##
## LEF for PtnCells ;
## created by Innovus v15.20-p005_1 on Mon Jun 14 16:49:06 2021
##

VERSION 5.7 ;

BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO DSP
  CLASS BLOCK ;
  SIZE 210.2200 BY 444.7200 ;
  FOREIGN DSP 0.0000 0.0000 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y R90 ;
  PIN top_N1BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.02765 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.209 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 16.6692 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 83.2685 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 14.9768 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 74.648 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 13.9450 444.3900 14.1150 444.7200 ;
    END
  END top_N1BEG[3]
  PIN top_N1BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.60565 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.889 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.1716 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.7805 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.5417 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.5375 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 43.633 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 233.176 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 41.2308 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 220.368 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 12.5650 444.3900 12.7350 444.7200 ;
    END
  END top_N1BEG[2]
  PIN top_N1BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 25.996 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 129.903 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 11.9628 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 59.696 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 11.1850 444.3900 11.3550 444.7200 ;
    END
  END top_N1BEG[1]
  PIN top_N1BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.54785 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.821 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.0832 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.1413 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.5565 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 52.351 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 279.672 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 48.2088 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 257.584 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 10.2650 444.3900 10.4350 444.7200 ;
    END
  END top_N1BEG[0]
  PIN top_N2BEG[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.91205 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.073 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.6868 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 3.3565 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.9784 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.774 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 24.9850 444.3900 25.1550 444.7200 ;
    END
  END top_N2BEG[7]
  PIN top_N2BEG[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.27625 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.325 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.0564 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 5.2045 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.1829 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.6685 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.1249 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.136 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 33.6078 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 179.712 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 23.6050 444.3900 23.7750 444.7200 ;
    END
  END top_N2BEG[6]
  PIN top_N2BEG[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.25885 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.481 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.3308 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 6.5765 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 10.4116 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 51.94 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 22.2250 444.3900 22.3950 444.7200 ;
    END
  END top_N2BEG[5]
  PIN top_N2BEG[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.16065 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.189 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 3.1984 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 15.9145 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.3308 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 11.536 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 20.8450 444.3900 21.0150 444.7200 ;
    END
  END top_N2BEG[4]
  PIN top_N2BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.62305 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.733 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 6.9686 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 34.7655 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 10.84 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 54.082 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 19.4650 444.3900 19.6350 444.7200 ;
    END
  END top_N2BEG[3]
  PIN top_N2BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.60565 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.889 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 13.13 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 65.5725 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.4072 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.918 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 18.0850 444.3900 18.2550 444.7200 ;
    END
  END top_N2BEG[2]
  PIN top_N2BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.50745 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.597 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 11.506 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 57.4525 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 8.0244 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 39.886 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 16.7050 444.3900 16.8750 444.7200 ;
    END
  END top_N2BEG[1]
  PIN top_N2BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.73865 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.869 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 6.1104 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 30.4745 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.3411 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.5345 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 25.6716 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 137.856 LAYER met3  ;
    PORT
      LAYER li1 ;
        RECT 15.3250 444.3900 15.4950 444.7200 ;
    END
  END top_N2BEG[0]
  PIN top_N2BEGb[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.91205 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.073 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.1716 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.7805 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.6687 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.1725 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.538 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 3.336 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 49.0518 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 262.08 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 35.5650 444.3900 35.7350 444.7200 ;
    END
  END top_N2BEGb[7]
  PIN top_N2BEGb[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.79645 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.937 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 2.7952 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 13.8985 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 16.0887 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 80.2725 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.262 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.864 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 4.7418 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 25.76 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 34.1850 444.3900 34.3550 444.7200 ;
    END
  END top_N2BEGb[6]
  PIN top_N2BEGb[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.33405 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.393 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 5.9032 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 29.4385 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 11.716 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 58.226 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 33.2650 444.3900 33.4350 444.7200 ;
    END
  END top_N2BEGb[5]
  PIN top_N2BEGb[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.25885 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.481 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.524 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 7.5425 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 3.0419 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.9205 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.642 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 9.224 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 55.6968 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 297.52 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 31.8850 444.3900 32.0550 444.7200 ;
    END
  END top_N2BEGb[4]
  PIN top_N2BEGb[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.136 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.16 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.0832 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.1335 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.5355 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 5.92 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 32.04 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 44.5248 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 237.936 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 30.5050 444.3900 30.6750 444.7200 ;
    END
  END top_N2BEGb[3]
  PIN top_N2BEGb[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.39185 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.461 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.8292 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 9.0685 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 18.9276 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 94.402 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 29.1250 444.3900 29.2950 444.7200 ;
    END
  END top_N2BEGb[2]
  PIN top_N2BEGb[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.39185 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.461 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.6224 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 3.0345 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.9435 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.5465 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.1249 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.136 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 50.3328 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 268.912 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 27.7450 444.3900 27.9150 444.7200 ;
    END
  END top_N2BEGb[1]
  PIN top_N2BEGb[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.66345 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.957 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.3004 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.4245 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.6897 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.2775 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.883 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 5.176 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 44.9856 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 240.864 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 26.3650 444.3900 26.5350 444.7200 ;
    END
  END top_N2BEGb[0]
  PIN top_N4BEG[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.66345 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.957 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.236 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.1025 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 5.3423 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 26.5405 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 15.6618 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 84 LAYER met3  ;
    PORT
      LAYER li1 ;
        RECT 57.1850 444.3900 57.3550 444.7200 ;
    END
  END top_N4BEG[15]
  PIN top_N4BEG[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.79645 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.937 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 10.778 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 53.8125 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 6.5908 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 32.718 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 56.2650 444.3900 56.4350 444.7200 ;
    END
  END top_N4BEG[14]
  PIN top_N4BEG[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.20105 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.413 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.6224 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 3.0345 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 4.9979 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 24.8185 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 6.6598 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 36.456 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 30.7758 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 164.608 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 54.8850 444.3900 55.0550 444.7200 ;
    END
  END top_N4BEG[13]
  PIN top_N4BEG[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.43225 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.685 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.3004 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.4245 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 2.3715 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 11.6865 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 11.554 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 62.088 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 16.4058 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 87.968 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 53.5050 444.3900 53.6750 444.7200 ;
    END
  END top_N4BEG[12]
  PIN top_N4BEG[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.43225 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.685 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.1716 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.7805 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.8801 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.2295 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.159 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 6.648 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 105.584 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 563.584 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 52.1250 444.3900 52.2950 444.7200 ;
    END
  END top_N4BEG[11]
  PIN top_N4BEG[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.10285 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.121 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.9104 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 9.4745 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.2057 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.8575 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 23.446 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 125.512 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 81.4278 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 434.752 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 50.7450 444.3900 50.9150 444.7200 ;
    END
  END top_N4BEG[10]
  PIN top_N4BEG[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.43225 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.685 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.3648 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.7465 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 3.6033 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 17.7275 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.469 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.968 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 102.487 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 548.48 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 49.3650 444.3900 49.5350 444.7200 ;
    END
  END top_N4BEG[9]
  PIN top_N4BEG[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.79645 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.937 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.0832 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.1803 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.6615 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.297 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 7.384 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 113.819 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 607.504 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 47.9850 444.3900 48.1550 444.7200 ;
    END
  END top_N4BEG[8]
  PIN top_N4BEG[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.25885 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.481 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.0832 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.2295 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.9765 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 6.586 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 35.592 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 128.474 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 686.608 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 46.6050 444.3900 46.7750 444.7200 ;
    END
  END top_N4BEG[7]
  PIN top_N4BEG[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.31665 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.549 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 2.7784 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 13.8145 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 2.7439 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 13.5485 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 3.16 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 17.32 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 122.284 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 653.12 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 45.2250 444.3900 45.3950 444.7200 ;
    END
  END top_N4BEG[6]
  PIN top_N4BEG[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.25885 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.481 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.0832 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.2295 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.9765 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 5.827 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 31.544 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 126.08 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 672.896 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 43.8450 444.3900 44.0150 444.7200 ;
    END
  END top_N4BEG[5]
  PIN top_N4BEG[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.44965 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.529 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.1716 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.7805 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.4689 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.1735 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.1249 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.136 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 129.079 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 689.36 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 42.4650 444.3900 42.6350 444.7200 ;
    END
  END top_N4BEG[4]
  PIN top_N4BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.91205 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.073 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 2.0056 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 9.9505 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.1036 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.455 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.1249 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.136 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 121.805 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 651.04 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 41.0850 444.3900 41.2550 444.7200 ;
    END
  END top_N4BEG[3]
  PIN top_N4BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.79645 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.937 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.0832 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.1803 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.6615 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 2.746 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 15.112 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 129.238 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 690.208 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 39.7050 444.3900 39.8750 444.7200 ;
    END
  END top_N4BEG[2]
  PIN top_N4BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.43225 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.685 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.236 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.1025 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.55 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.632 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 38.3250 444.3900 38.4950 444.7200 ;
    END
  END top_N4BEG[1]
  PIN top_N4BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.21845 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.257 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 20.5668 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 102.757 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.8828 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.296 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 36.9450 444.3900 37.1150 444.7200 ;
    END
  END top_N4BEG[0]
  PIN top_NN4BEG[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.16065 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.189 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.6868 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 3.3565 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 6.8457 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 33.9395 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 1.9128 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 10.672 LAYER met3  ;
    PORT
      LAYER li1 ;
        RECT 79.2650 444.3900 79.4350 444.7200 ;
    END
  END top_NN4BEG[15]
  PIN top_NN4BEG[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.68085 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.801 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.4936 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 2.3905 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 15.8716 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 79.24 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 77.8850 444.3900 78.0550 444.7200 ;
    END
  END top_NN4BEG[14]
  PIN top_NN4BEG[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.91205 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.073 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 6.5948 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 32.8965 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 6.8892 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 34.328 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 76.5050 444.3900 76.6750 444.7200 ;
    END
  END top_NN4BEG[13]
  PIN top_NN4BEG[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.39185 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.461 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.0732 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 5.2885 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 11.0582 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 55.055 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 75.1250 444.3900 75.2950 444.7200 ;
    END
  END top_NN4BEG[12]
  PIN top_NN4BEG[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.91205 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.073 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.0832 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.6253 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.9555 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.573 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 8.856 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 80.5128 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 429.872 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 73.7450 444.3900 73.9150 444.7200 ;
    END
  END top_NN4BEG[11]
  PIN top_NN4BEG[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.68085 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.801 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.0564 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 5.2045 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 4.1173 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 20.4155 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.469 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.968 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 107.303 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 572.752 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 72.3650 444.3900 72.5350 444.7200 ;
    END
  END top_NN4BEG[10]
  PIN top_NN4BEG[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.16065 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.189 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.0832 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.1945 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.8015 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 26.986 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 144.392 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 102.464 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 546.944 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 70.9850 444.3900 71.1550 444.7200 ;
    END
  END top_NN4BEG[9]
  PIN top_NN4BEG[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.68085 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.801 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.0832 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.2785 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.2215 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 18.5968 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 100.12 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 75.3168 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 402.16 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 69.6050 444.3900 69.7750 444.7200 ;
    END
  END top_NN4BEG[8]
  PIN top_NN4BEG[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.91205 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.073 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.7512 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 3.6785 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 2.0957 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.3075 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.607 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 3.704 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 121.576 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 649.344 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 68.2250 444.3900 68.3950 444.7200 ;
    END
  END top_NN4BEG[7]
  PIN top_NN4BEG[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.43225 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.685 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.3648 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.7465 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 2.9049 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.3535 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.814 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 4.808 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 118.784 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 633.984 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 66.8450 444.3900 67.0150 444.7200 ;
    END
  END top_NN4BEG[6]
  PIN top_NN4BEG[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.43225 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.685 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.0832 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.55 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.632 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 65.4650 444.3900 65.6350 444.7200 ;
    END
  END top_NN4BEG[5]
  PIN top_NN4BEG[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.31665 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.549 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.236 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.1025 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.0736 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.25 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 64.0850 444.3900 64.2550 444.7200 ;
    END
  END top_NN4BEG[4]
  PIN top_NN4BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.20105 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.413 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.88 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 4.3225 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.2771 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.2145 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.331 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.232 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 128.045 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 683.376 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 62.7050 444.3900 62.8750 444.7200 ;
    END
  END top_NN4BEG[3]
  PIN top_NN4BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.91205 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.073 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.0832 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.9784 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.774 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 61.3250 444.3900 61.4950 444.7200 ;
    END
  END top_NN4BEG[2]
  PIN top_NN4BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.73865 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.869 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.6868 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 3.3565 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.2309 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.9835 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.331 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.232 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 130.25 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 695.136 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 59.9450 444.3900 60.1150 444.7200 ;
    END
  END top_NN4BEG[1]
  PIN top_NN4BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.43225 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.685 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.1716 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.7805 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.5692 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.728 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 58.5650 444.3900 58.7350 444.7200 ;
    END
  END top_NN4BEG[0]
  PIN top_S1END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.43225 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.685 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.7512 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 3.6785 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 3.0547 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 15.1025 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.745 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 4.44 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.5156 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 6.8496 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 37.472 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 84.3250 444.3900 84.4950 444.7200 ;
    END
  END top_S1END[3]
  PIN top_S1END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.20105 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.413 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.8156 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 4.0005 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.2771 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.2145 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.331 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.232 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.5156 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 29.4024 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 157.744 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 82.9450 444.3900 83.1150 444.7200 ;
    END
  END top_S1END[2]
  PIN top_S1END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.33405 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.393 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.6224 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 3.0345 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.5012 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 25.4784 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 125.986 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 81.5650 444.3900 81.7350 444.7200 ;
    END
  END top_S1END[1]
  PIN top_S1END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.10285 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.121 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 2.3444 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 11.6445 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.1872 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 3.5879 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 17.6505 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.5012 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 13.3476 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 72.128 LAYER met3  ;
    PORT
      LAYER li1 ;
        RECT 80.1850 444.3900 80.3550 444.7200 ;
    END
  END top_S1END[0]
  PIN top_S2MID[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.66345 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.957 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.1716 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.7805 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.6057 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.8575 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 9.208 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 49.576 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.8792 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 48.9168 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 261.36 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 105.9450 444.3900 106.1150 444.7200 ;
    END
  END top_S2MID[7]
  PIN top_S2MID[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.43225 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.685 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.0832 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.1595 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.6055 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 6.679 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 36.088 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.512 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 57.4155 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 307.152 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 104.5650 444.3900 104.7350 444.7200 ;
    END
  END top_S2MID[6]
  PIN top_S2MID[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.43225 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.685 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.0832 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.1115 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.3865 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 4.354 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 23.688 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.692 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 59.9916 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 320.896 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 103.1850 444.3900 103.3550 444.7200 ;
    END
  END top_S2MID[5]
  PIN top_S2MID[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.58865 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.869 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.0832 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 2.3071 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 11.3645 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 2.677 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 14.744 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.512 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 116.421 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 623.728 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 102.2650 444.3900 102.4350 444.7200 ;
    END
  END top_S2MID[4]
  PIN top_S2MID[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.62305 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.733 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.2664 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 6.2545 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.5217 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.4375 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 7 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 37.8 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.8828 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 86.8311 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 464.976 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 100.8850 444.3900 101.0550 444.7200 ;
    END
  END top_S2MID[3]
  PIN top_S2MID[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.96985 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.141 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.4596 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 7.2205 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.5777 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.7175 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 2.677 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 14.744 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.7028 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 78.5292 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 420.704 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 99.5050 444.3900 99.6750 444.7200 ;
    END
  END top_S2MID[2]
  PIN top_S2MID[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.31665 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.549 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.2664 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 6.2545 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.8913 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.2855 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.711 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 9.592 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.8756 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 111.181 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 594.832 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 98.1250 444.3900 98.2950 444.7200 ;
    END
  END top_S2MID[1]
  PIN top_S2MID[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.43225 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.685 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.7512 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 3.6785 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 3.7603 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 18.6305 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.504 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 8.488 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.6992 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 95.8941 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 513.312 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 96.7450 444.3900 96.9150 444.7200 ;
    END
  END top_S2MID[0]
  PIN top_S2END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.68085 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.801 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 2.0392 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 10.1185 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.3744 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 20.0221 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 99.5855 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.5652 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 10.5208 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 57.048 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.1304 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 6.7167 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 36.288 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 95.3650 444.3900 95.5350 444.7200 ;
    END
  END top_S2END[7]
  PIN top_S2END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.31665 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.549 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 4.0356 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 20.1005 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.6089 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.8735 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 10.588 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 56.936 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.9432 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 32.616 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 175.824 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 93.9850 444.3900 94.1550 444.7200 ;
    END
  END top_S2END[6]
  PIN top_S2END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.20105 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.413 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.6868 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 3.3565 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.9432 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 7.3756 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 36.19 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 92.6050 444.3900 92.7750 444.7200 ;
    END
  END top_S2END[5]
  PIN top_S2END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.25925 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.305 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 8.3686 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 41.7655 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.756 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 19.1945 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 95.3295 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.9432 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 3.4308 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 18.768 LAYER met3  ;
    PORT
      LAYER li1 ;
        RECT 91.2250 444.3900 91.3950 444.7200 ;
    END
  END top_S2END[4]
  PIN top_S2END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.33405 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.393 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 5.0016 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 24.9305 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.5652 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 7.7209 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 37.9715 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.1304 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 9.4746 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 50.992 LAYER met3  ;
    PORT
      LAYER li1 ;
        RECT 89.8450 444.3900 90.0150 444.7200 ;
    END
  END top_S2END[3]
  PIN top_S2END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.39185 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.461 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 14.9808 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 74.8265 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.9432 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 28.8437 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 142.887 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.9432 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 1.228 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 7.016 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.1304 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 4.7418 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 25.76 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 88.4650 444.3900 88.6350 444.7200 ;
    END
  END top_S2END[2]
  PIN top_S2END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.66345 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.957 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.0832 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 6.5589 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 32.6235 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.1304 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 31.0416 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 166.016 LAYER met3  ;
    PORT
      LAYER li1 ;
        RECT 87.0850 444.3900 87.2550 444.7200 ;
    END
  END top_S2END[1]
  PIN top_S2END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.20105 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.413 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.3648 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.7465 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 4.2055 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 20.8565 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.5688 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 18.0598 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 96.776 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.134 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 22.0626 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 118.608 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 85.7050 444.3900 85.8750 444.7200 ;
    END
  END top_S2END[0]
  PIN top_S4END[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.37445 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.617 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 16.1708 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 80.7765 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 4.834 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 24.052 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 10.8527 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 41.9306 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 127.5650 444.3900 127.7350 444.7200 ;
    END
  END top_S4END[15]
  PIN top_S4END[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.50745 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.597 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 4.6936 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 23.3905 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 3.5752 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 17.64 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 8.08613 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 37.5859 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 126.1850 444.3900 126.3550 444.7200 ;
    END
  END top_S4END[14]
  PIN top_S4END[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.91205 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.073 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 12.232 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 61.0085 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 30.4729 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 151.721 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 6.8808 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 37.168 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met3  ;
    ANTENNAMAXAREACAR 13.5457 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 70.0458 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.123098 LAYER via3  ;
    PORT
      LAYER li1 ;
        RECT 125.2650 444.3900 125.4350 444.7200 ;
    END
  END top_S4END[13]
  PIN top_S4END[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.43225 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.685 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 2.6188 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 13.0165 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 9.8656 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 49.21 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 13.6954 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 67.1731 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 123.8850 444.3900 124.0550 444.7200 ;
    END
  END top_S4END[12]
  PIN top_S4END[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.14325 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.345 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 2.0868 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 10.3565 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 2.2469 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 11.0635 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 11.3904 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 64.512 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met3  ;
    ANTENNAMAXAREACAR 22.0626 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 118.174 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.123098 LAYER via3  ;
    PORT
      LAYER li1 ;
        RECT 122.5050 444.3900 122.6750 444.7200 ;
    END
  END top_S4END[11]
  PIN top_S4END[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.73865 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.869 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.236 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.1025 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 9.8919 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 49.0525 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 7.494 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 42.32 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met3  ;
    ANTENNAMAXAREACAR 17.6998 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 93.497 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.123098 LAYER via3  ;
    PORT
      LAYER li1 ;
        RECT 121.1250 444.3900 121.2950 444.7200 ;
    END
  END top_S4END[10]
  PIN top_S4END[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.73865 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.869 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 3.5512 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 17.6785 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 28.7517 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 142.762 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.3416 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 8.096 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met3  ;
    ANTENNAMAXAREACAR 8.51077 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 41.9636 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.123098 LAYER via3  ;
    PORT
      LAYER li1 ;
        RECT 119.7450 444.3900 119.9150 444.7200 ;
    END
  END top_S4END[9]
  PIN top_S4END[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.66345 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.957 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.0832 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 5.17 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 25.732 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 7.37131 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 35.5529 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 118.3650 444.3900 118.5350 444.7200 ;
    END
  END top_S4END[8]
  PIN top_S4END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.62305 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.733 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.4428 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 7.1365 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.3261 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.4595 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.331 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.232 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.9504 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 96.1257 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 513.136 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 116.9850 444.3900 117.1550 444.7200 ;
    END
  END top_S4END[7]
  PIN top_S4END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.54785 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.821 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.88 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 4.3225 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.4433 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.0455 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.4 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.6 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.9432 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 104.957 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 560.24 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 115.6050 444.3900 115.7750 444.7200 ;
    END
  END top_S4END[6]
  PIN top_S4END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.136 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.16 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 6.3204 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 31.5245 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.2897 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.2775 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 15.676 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 84.072 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.9468 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 110.222 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 589.728 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 114.2250 444.3900 114.3950 444.7200 ;
    END
  END top_S4END[5]
  PIN top_S4END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.22145 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.437 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 19.6138 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 97.9545 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.9504 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 10.586 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 51.898 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 112.8450 444.3900 113.0150 444.7200 ;
    END
  END top_S4END[4]
  PIN top_S4END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.66345 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.957 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.0832 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.5688 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 12.4227 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 61.3725 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.5688 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 4.057 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 22.104 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.9468 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 1.7658 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 9.888 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 111.4650 444.3900 111.6350 444.7200 ;
    END
  END top_S4END[3]
  PIN top_S4END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.16065 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.189 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 5.3828 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 26.7995 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.3583 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.6205 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 12.403 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 66.616 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.9468 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 47.6601 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 256.064 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 110.0850 444.3900 110.2550 444.7200 ;
    END
  END top_S4END[2]
  PIN top_S4END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.68085 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.801 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.3784 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 6.8145 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 7.0475 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 35.0665 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.5724 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 21.976 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 118.128 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.9504 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 7.4868 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 40.4 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 108.7050 444.3900 108.8750 444.7200 ;
    END
  END top_S4END[1]
  PIN top_S4END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.20105 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.413 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 2.7952 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 13.8985 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.2771 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.2145 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.1249 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.136 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.9468 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 16.7556 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 90.304 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 107.3250 444.3900 107.4950 444.7200 ;
    END
  END top_S4END[0]
  PIN top_SS4END[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.12625 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.325 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.0832 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 2.202 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.892 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 3.66653 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 16.938 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 149.1850 444.3900 149.3550 444.7200 ;
    END
  END top_SS4END[15]
  PIN top_SS4END[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.68085 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.801 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 3.5848 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 17.8465 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.4544 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.154 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 2.74606 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 11.3421 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 148.2650 444.3900 148.4350 444.7200 ;
    END
  END top_SS4END[14]
  PIN top_SS4END[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.33405 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.393 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 8.092 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 40.376 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 38.698 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 193.018 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 53.1663 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 263.96 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 146.8850 444.3900 147.0550 444.7200 ;
    END
  END top_SS4END[13]
  PIN top_SS4END[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.91205 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.073 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.1716 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.7805 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 2.678 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 13.272 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 4.82801 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 22.7455 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 145.5050 444.3900 145.6750 444.7200 ;
    END
  END top_SS4END[12]
  PIN top_SS4END[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.20105 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.413 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.524 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 7.5425 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 7.4716 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 37.24 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 10.4711 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 51.0519 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 144.1250 444.3900 144.2950 444.7200 ;
    END
  END top_SS4END[11]
  PIN top_SS4END[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.54785 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.821 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.1376 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 5.6105 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 7.096 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 35.126 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 10.171 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 49.1428 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 142.7450 444.3900 142.9150 444.7200 ;
    END
  END top_SS4END[10]
  PIN top_SS4END[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.33405 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.393 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 2.0224 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 10.0345 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 2.4568 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 12.166 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 3.71717 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 17.2822 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 141.3650 444.3900 141.5350 444.7200 ;
    END
  END top_SS4END[9]
  PIN top_SS4END[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.79645 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.937 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 8.5548 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 42.6965 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.7065 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.3615 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.3416 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 8.096 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met3  ;
    ANTENNAMAXAREACAR 28.6875 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 143.773 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.123098 LAYER via3  ;
    PORT
      LAYER li1 ;
        RECT 139.9850 444.3900 140.1550 444.7200 ;
    END
  END top_SS4END[8]
  PIN top_SS4END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.79645 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.937 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.4936 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 2.3905 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.1803 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.6615 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.538 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 3.336 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.378 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 78.4506 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 419.344 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 138.6050 444.3900 138.7750 444.7200 ;
    END
  END top_SS4END[7]
  PIN top_SS4END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.66345 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.957 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.0832 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.2379 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.0185 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 8.977 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 48.344 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.5688 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 110.413 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 589.808 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 137.2250 444.3900 137.3950 444.7200 ;
    END
  END top_SS4END[6]
  PIN top_SS4END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.56525 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.665 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 4.8084 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 23.9645 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.1423 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.5405 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.1905 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.464 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.5688 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 122.045 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 652.32 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 135.8450 444.3900 136.0150 444.7200 ;
    END
  END top_SS4END[5]
  PIN top_SS4END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.56525 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.665 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.3308 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 6.5765 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 2.4457 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 12.0575 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.814 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 4.808 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.5652 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 109.133 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 583.92 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 134.4650 444.3900 134.6350 444.7200 ;
    END
  END top_SS4END[4]
  PIN top_SS4END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.37445 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.617 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.8156 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 4.0005 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.9029 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.3435 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.4 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.6 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.378 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 28.8576 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 154.848 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 133.0850 444.3900 133.2550 444.7200 ;
    END
  END top_SS4END[3]
  PIN top_SS4END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.37445 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.617 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.0832 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.4759 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.2085 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.331 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.232 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.5688 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 36.0348 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 192.656 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 131.7050 444.3900 131.8750 444.7200 ;
    END
  END top_SS4END[2]
  PIN top_SS4END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.96985 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.141 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.4596 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 7.2205 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.5688 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 17.6814 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 87.955 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 130.3250 444.3900 130.4950 444.7200 ;
    END
  END top_SS4END[1]
  PIN top_SS4END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.66345 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.957 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.7512 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 3.6785 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.378 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 13.0328 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 64.659 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.5652 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 13.1478 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 70.592 LAYER met3  ;
    PORT
      LAYER li1 ;
        RECT 128.9450 444.3900 129.1150 444.7200 ;
    END
  END top_SS4END[0]
  PIN top_E1BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2063 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.7315 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 16.0788 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 86.224 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 209.7350 309.8400 210.2200 309.9800 ;
    END
  END top_E1BEG[3]
  PIN top_E1BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.9342 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.445 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 209.7350 308.4800 210.2200 308.6200 ;
    END
  END top_E1BEG[2]
  PIN top_E1BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 7.1327 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 35.4375 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 209.7350 306.7800 210.2200 306.9200 ;
    END
  END top_E1BEG[1]
  PIN top_E1BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 8.2212 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 40.88 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 209.7350 305.4200 210.2200 305.5600 ;
    END
  END top_E1BEG[0]
  PIN top_E2BEG[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.2433 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.9375 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 24.2208 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 129.648 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 209.7350 321.7400 210.2200 321.8800 ;
    END
  END top_E2BEG[7]
  PIN top_E2BEG[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1253 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.4655 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 35.4858 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 189.728 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 209.7350 320.0400 210.2200 320.1800 ;
    END
  END top_E2BEG[6]
  PIN top_E2BEG[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1449 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.5635 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 40.6848 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 217.456 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 209.7350 318.6800 210.2200 318.8200 ;
    END
  END top_E2BEG[5]
  PIN top_E2BEG[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1645 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.6615 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 16.108 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 86.376 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 0.8508 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 5.008 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 209.7350 317.3200 210.2200 317.4600 ;
    END
  END top_E2BEG[4]
  PIN top_E2BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.3481 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.6325 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 209.7350 315.6200 210.2200 315.7600 ;
    END
  END top_E2BEG[3]
  PIN top_E2BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.198 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.882 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 209.7350 314.2600 210.2200 314.4000 ;
    END
  END top_E2BEG[2]
  PIN top_E2BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 4.8204 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 23.758 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 209.7350 312.9000 210.2200 313.0400 ;
    END
  END top_E2BEG[1]
  PIN top_E2BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.1028 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 209.7350 311.2000 210.2200 311.3400 ;
    END
  END top_E2BEG[0]
  PIN top_E2BEGb[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.5409 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.4255 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 35.9928 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 192.432 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 209.7350 333.3000 210.2200 333.4400 ;
    END
  END top_E2BEGb[7]
  PIN top_E2BEGb[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.5264 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.471 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 16.2648 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 87.216 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 209.7350 331.9400 210.2200 332.0800 ;
    END
  END top_E2BEGb[6]
  PIN top_E2BEGb[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.2515 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.1495 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 209.7350 330.5800 210.2200 330.7200 ;
    END
  END top_E2BEGb[5]
  PIN top_E2BEGb[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.198 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.882 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 209.7350 328.8800 210.2200 329.0200 ;
    END
  END top_E2BEGb[4]
  PIN top_E2BEGb[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.266 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.169 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 35.149 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 187.928 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 2.3148 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 12.816 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 209.7350 327.5200 210.2200 327.6600 ;
    END
  END top_E2BEGb[3]
  PIN top_E2BEGb[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1841 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.7595 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 25.2738 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 135.264 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 209.7350 326.1600 210.2200 326.3000 ;
    END
  END top_E2BEGb[2]
  PIN top_E2BEGb[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.9631 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.7075 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 209.7350 324.4600 210.2200 324.6000 ;
    END
  END top_E2BEGb[1]
  PIN top_E2BEGb[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.5572 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.56 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 209.7350 323.1000 210.2200 323.2400 ;
    END
  END top_E2BEGb[0]
  PIN top_EE4BEG[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.42 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.939 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 32.7288 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 175.024 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 209.7350 357.1000 210.2200 357.2400 ;
    END
  END top_EE4BEG[15]
  PIN top_EE4BEG[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.3083 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.2355 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 38.2938 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 204.704 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 209.7350 355.4000 210.2200 355.5400 ;
    END
  END top_EE4BEG[14]
  PIN top_EE4BEG[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.8393 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 18.9175 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 22.384 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 119.848 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 0.4848 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 3.056 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 209.7350 354.0400 210.2200 354.1800 ;
    END
  END top_EE4BEG[13]
  PIN top_EE4BEG[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1673 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.6755 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 26.9328 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 144.112 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 209.7350 352.6800 210.2200 352.8200 ;
    END
  END top_EE4BEG[12]
  PIN top_EE4BEG[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1491 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.5845 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 29.8278 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 159.552 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 209.7350 350.9800 210.2200 351.1200 ;
    END
  END top_EE4BEG[11]
  PIN top_EE4BEG[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1687 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.6825 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 11.968 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 64.296 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 0.4848 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 3.056 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 209.7350 349.6200 210.2200 349.7600 ;
    END
  END top_EE4BEG[10]
  PIN top_EE4BEG[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1883 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.7805 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 25.327 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 135.544 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 2.4336 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 13.92 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 209.7350 348.2600 210.2200 348.4000 ;
    END
  END top_EE4BEG[9]
  PIN top_EE4BEG[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1365 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.5215 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 15.877 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 85.144 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 1.3356 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 8.064 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 209.7350 346.5600 210.2200 346.7000 ;
    END
  END top_EE4BEG[8]
  PIN top_EE4BEG[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.288 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.279 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 31.123 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 166.456 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 1.5186 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 9.04 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 209.7350 345.2000 210.2200 345.3400 ;
    END
  END top_EE4BEG[7]
  PIN top_EE4BEG[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1239 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.4585 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 38.5218 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 205.92 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 209.7350 343.8400 210.2200 343.9800 ;
    END
  END top_EE4BEG[6]
  PIN top_EE4BEG[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2009 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.8435 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 7.183 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 38.776 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 1.3356 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 8.064 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 209.7350 342.1400 210.2200 342.2800 ;
    END
  END top_EE4BEG[5]
  PIN top_EE4BEG[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.399 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.834 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 11.509 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 61.848 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 1.3356 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 8.064 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 209.7350 340.7800 210.2200 340.9200 ;
    END
  END top_EE4BEG[4]
  PIN top_EE4BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.1028 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 209.7350 339.4200 210.2200 339.5600 ;
    END
  END top_EE4BEG[3]
  PIN top_EE4BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1799 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.7385 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 17.0548 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 91.896 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 1.5186 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 9.04 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 209.7350 337.7200 210.2200 337.8600 ;
    END
  END top_EE4BEG[2]
  PIN top_EE4BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.2278 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.978 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 56.9148 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 304.016 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 209.7350 336.3600 210.2200 336.5000 ;
    END
  END top_EE4BEG[1]
  PIN top_EE4BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.0468 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.126 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 209.7350 335.0000 210.2200 335.1400 ;
    END
  END top_EE4BEG[0]
  PIN top_E6BEG[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1477 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.5775 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 28.6788 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 153.424 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 209.7350 374.7800 210.2200 374.9200 ;
    END
  END top_E6BEG[11]
  PIN top_E6BEG[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.4098 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.888 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 52.216 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 278.952 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 1.3356 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 8.064 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 209.7350 373.0800 210.2200 373.2200 ;
    END
  END top_E6BEG[10]
  PIN top_E6BEG[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1575 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.6265 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 26.0568 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 139.44 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 209.7350 371.7200 210.2200 371.8600 ;
    END
  END top_E6BEG[9]
  PIN top_E6BEG[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.6132 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.905 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 10.0998 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 54.336 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 209.7350 370.3600 210.2200 370.5000 ;
    END
  END top_E6BEG[8]
  PIN top_E6BEG[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1561 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.6195 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 36.019 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 192.568 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 2.5524 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 15.024 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 209.7350 368.6600 210.2200 368.8000 ;
    END
  END top_E6BEG[7]
  PIN top_E6BEG[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7404 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.423 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 10.543 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 56.696 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 0.6678 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 4.032 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 209.7350 367.3000 210.2200 367.4400 ;
    END
  END top_E6BEG[6]
  PIN top_E6BEG[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1897 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.7875 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 16.2618 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 87.2 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 209.7350 365.9400 210.2200 366.0800 ;
    END
  END top_E6BEG[5]
  PIN top_E6BEG[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1351 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.5145 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 9.4068 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 50.64 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 209.7350 364.2400 210.2200 364.3800 ;
    END
  END top_E6BEG[4]
  PIN top_E6BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.3267 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.3545 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 12.8568 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 69.04 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 209.7350 362.8800 210.2200 363.0200 ;
    END
  END top_E6BEG[3]
  PIN top_E6BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1813 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.7455 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 28.6368 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 153.2 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 209.7350 361.5200 210.2200 361.6600 ;
    END
  END top_E6BEG[2]
  PIN top_E6BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1995 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.8365 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 40.063 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 214.136 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 0.6678 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 4.032 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 209.7350 359.8200 210.2200 359.9600 ;
    END
  END top_E6BEG[1]
  PIN top_E6BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.1028 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 209.7350 358.4600 210.2200 358.6000 ;
    END
  END top_E6BEG[0]
  PIN top_E1END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.1872 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.7701 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.4105 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via2  ;
    ANTENNADIFFAREA 0.3744 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 6.2753 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 34.4 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via3  ;
    ANTENNADIFFAREA 2.0736 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 24.1881 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 130.88 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 309.8400 0.4850 309.9800 ;
    END
  END top_E1END[3]
  PIN top_E1END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.3113 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.2775 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 4.0646 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 22.136 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via3  ;
    ANTENNADIFFAREA 2.0736 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 12.6654 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 68.96 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 308.4800 0.4850 308.6200 ;
    END
  END top_E1END[2]
  PIN top_E1END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1883 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.7805 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 3.781 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 20.632 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.6992 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 7.9782 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 44.432 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 306.7800 0.4850 306.9200 ;
    END
  END top_E1END[1]
  PIN top_E1END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.8232 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.955 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 4.954 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 26.888 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.6992 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 26.6925 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 145.648 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 305.4200 0.4850 305.5600 ;
    END
  END top_E1END[0]
  PIN top_E2MID[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1435 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.5565 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 20.7386 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 111.064 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via3  ;
    ANTENNADIFFAREA 0.7632 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 13.4616 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 72.736 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 20.621 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 110.189 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 321.7400 0.4850 321.8800 ;
    END
  END top_E2MID[7]
  PIN top_E2MID[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1813 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.7455 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.5688 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 30.5016 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 163.616 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met3  ;
    ANTENNAMAXAREACAR 46.0671 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 243.134 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.123098 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 320.0400 0.4850 320.1800 ;
    END
  END top_E2MID[6]
  PIN top_E2MID[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1617 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.6475 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.262 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.864 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.7632 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 48.9792 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 263.104 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 74.0106 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 394.63 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 318.6800 0.4850 318.8200 ;
    END
  END top_E2MID[5]
  PIN top_E2MID[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.9773 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.6075 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 2.47 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 13.64 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.5688 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 44.0064 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 236.112 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 75.821 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 403.005 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 317.3200 0.4850 317.4600 ;
    END
  END top_E2MID[4]
  PIN top_E2MID[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1603 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.6405 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.7632 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 11.8458 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 63.648 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met3  ;
    ANTENNAMAXAREACAR 29.7908 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 152.527 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.153401 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 315.6200 0.4850 315.7600 ;
    END
  END top_E2MID[3]
  PIN top_E2MID[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1407 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.5425 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.5688 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 19.8018 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 106.08 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met3  ;
    ANTENNAMAXAREACAR 37.1356 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 192.954 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.123098 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 314.2600 0.4850 314.4000 ;
    END
  END top_E2MID[2]
  PIN top_E2MID[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2791 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.1165 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.7632 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 50.2713 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 269.52 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met3  ;
    ANTENNAMAXAREACAR 80.3962 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 424.978 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.123098 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 312.9000 0.4850 313.0400 ;
    END
  END top_E2MID[1]
  PIN top_E2MID[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 7.5689 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 37.5655 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 6.5917 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 36.096 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.5688 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 19.2198 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 105.328 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 51.4245 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 276.451 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 311.2000 0.4850 311.3400 ;
    END
  END top_E2MID[0]
  PIN top_E2END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.5724 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 6.1059 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 29.6905 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.954 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 5.0868 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 27.6 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 333.3000 0.4850 333.4400 ;
    END
  END top_E2END[7]
  PIN top_E2END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1673 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.6755 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.7632 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 9.1588 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 49.304 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.1448 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 2.0034 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 12.096 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 331.9400 0.4850 332.0800 ;
    END
  END top_E2END[6]
  PIN top_E2END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.1448 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 12.7972 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 62.482 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 330.5800 0.4850 330.7200 ;
    END
  END top_E2END[5]
  PIN top_E2END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.6069 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.8735 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 11.968 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 64.296 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.9468 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 7.3248 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 41.888 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 328.8800 0.4850 329.0200 ;
    END
  END top_E2END[4]
  PIN top_E2END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.8359 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.9005 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 10.057 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 54.104 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.5156 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 5.9346 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 32.592 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 327.5200 0.4850 327.6600 ;
    END
  END top_E2END[3]
  PIN top_E2END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.5985 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 17.7135 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.332 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 39.9186 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 213.36 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 326.1600 0.4850 326.3000 ;
    END
  END top_E2END[2]
  PIN top_E2END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.8701 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 19.0715 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.1905 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.464 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.756 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 4.5108 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 24.528 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 324.4600 0.4850 324.6000 ;
    END
  END top_E2END[1]
  PIN top_E2END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1239 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.4585 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 11.1926 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 60.152 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via3  ;
    ANTENNADIFFAREA 0.7632 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 27.2415 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 148.576 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 323.1000 0.4850 323.2400 ;
    END
  END top_E2END[0]
  PIN top_EE4END[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.5054 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.366 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 30.2418 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 161.76 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met3  ;
    ANTENNAMAXAREACAR 44.6877 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 235.487 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.123098 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 357.1000 0.4850 357.2400 ;
    END
  END top_EE4END[15]
  PIN top_EE4END[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1785 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.7315 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 36.7758 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 196.608 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met3  ;
    ANTENNAMAXAREACAR 51.0821 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 268.589 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.123098 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 355.4000 0.4850 355.5400 ;
    END
  END top_EE4END[14]
  PIN top_EE4END[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.0468 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.126 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 3.27919 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 15.0148 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 354.0400 0.4850 354.1800 ;
    END
  END top_EE4END[13]
  PIN top_EE4END[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7217 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.4475 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 22.6098 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 121.056 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met3  ;
    ANTENNAMAXAREACAR 33.7989 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 178.312 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.123098 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 352.6800 0.4850 352.8200 ;
    END
  END top_EE4END[12]
  PIN top_EE4END[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.224 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.894 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 7.2565 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 34.0465 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 350.9800 0.4850 351.1200 ;
    END
  END top_EE4END[11]
  PIN top_EE4END[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1379 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.5285 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 15.922 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 85.384 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 3.1014 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 17.952 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 6.8936 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 37.0411 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 349.6200 0.4850 349.7600 ;
    END
  END top_EE4END[10]
  PIN top_EE4END[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.1764 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.656 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 5.73387 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 27.1293 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 348.2600 0.4850 348.4000 ;
    END
  END top_EE4END[9]
  PIN top_EE4END[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1365 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.5215 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 34.1988 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 182.864 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met3  ;
    ANTENNAMAXAREACAR 52.7727 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 278.384 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.123098 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 346.5600 0.4850 346.7000 ;
    END
  END top_EE4END[8]
  PIN top_EE4END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.1219 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.3305 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 31.876 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 170.472 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 2.0676 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 11.968 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 14.9472 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 79.2162 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 345.2000 0.4850 345.3400 ;
    END
  END top_EE4END[7]
  PIN top_EE4END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.164 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.712 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 4.4369 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 20.8034 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 343.8400 0.4850 343.9800 ;
    END
  END top_EE4END[6]
  PIN top_EE4END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.2156 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.852 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 3.29212 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 14.9205 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 342.1400 0.4850 342.2800 ;
    END
  END top_EE4END[5]
  PIN top_EE4END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1813 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.7455 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 58.324 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 311.528 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.4848 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 3.056 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 3.29024 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 16.5253 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 340.7800 0.4850 340.9200 ;
    END
  END top_EE4END[4]
  PIN top_EE4END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.504 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.359 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.378 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 38.8878 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 207.872 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 339.4200 0.4850 339.5600 ;
    END
  END top_EE4END[3]
  PIN top_EE4END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.7918 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 23.695 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.1908 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 22.9459 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 122.84 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.5652 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 3.8334 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 21.856 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 337.7200 0.4850 337.8600 ;
    END
  END top_EE4END[2]
  PIN top_EE4END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.3361 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.4015 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 23.281 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 124.632 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.5724 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 3.3084 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 19.056 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 336.3600 0.4850 336.5000 ;
    END
  END top_EE4END[1]
  PIN top_EE4END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1407 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.5425 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.5724 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 34.5585 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 185.248 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 335.0000 0.4850 335.1400 ;
    END
  END top_EE4END[0]
  PIN top_E6END[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2331 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.0045 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 26.8428 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 143.632 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met3  ;
    ANTENNAMAXAREACAR 40.1614 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 211.032 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.123098 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 374.7800 0.4850 374.9200 ;
    END
  END top_E6END[11]
  PIN top_E6END[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.0673 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.0575 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 38.599 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 206.328 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.6678 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 4.032 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 7.19232 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 37.4451 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 373.0800 0.4850 373.2200 ;
    END
  END top_E6END[10]
  PIN top_E6END[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.9818 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.683 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 4.53845 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 21.1522 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 371.7200 0.4850 371.8600 ;
    END
  END top_E6END[9]
  PIN top_E6END[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1725 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.6405 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 36.0378 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 192.672 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met3  ;
    ANTENNAMAXAREACAR 50.2372 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 266.464 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.123098 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 370.3600 0.4850 370.5000 ;
    END
  END top_E6END[8]
  PIN top_E6END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2359 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.0185 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 20.197 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 108.184 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 1.8204 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 11.12 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 11.2176 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 58.9912 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 368.6600 0.4850 368.8000 ;
    END
  END top_E6END[7]
  PIN top_E6END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.1457 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.4495 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 36.5898 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 195.616 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met3  ;
    ANTENNAMAXAREACAR 51.697 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 272.927 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.123098 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 367.3000 0.4850 367.4400 ;
    END
  END top_E6END[6]
  PIN top_E6END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1897 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.7875 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 26.383 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 141.176 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 1.7016 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 10.016 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 27.549 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 146.943 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 365.9400 0.4850 366.0800 ;
    END
  END top_E6END[5]
  PIN top_E6END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.4732 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.205 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 28.0848 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 150.256 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met3  ;
    ANTENNAMAXAREACAR 42.5623 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 224.587 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.123098 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 364.2400 0.4850 364.3800 ;
    END
  END top_E6END[4]
  PIN top_E6END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1911 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.7945 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 11.83 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 63.56 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 1.2168 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 6.96 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 4.35993 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 20.9643 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 362.8800 0.4850 363.0200 ;
    END
  END top_E6END[3]
  PIN top_E6END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1253 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.4655 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 49.1898 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 262.816 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met3  ;
    ANTENNAMAXAREACAR 69.8845 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 369.977 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.123098 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 361.5200 0.4850 361.6600 ;
    END
  END top_E6END[2]
  PIN top_E6END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.4789 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.1155 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 15.577 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 83.544 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 2.2716 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 7.9878 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 43.072 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 359.8200 0.4850 359.9600 ;
    END
  END top_E6END[1]
  PIN top_E6END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.6305 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.8735 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 8.701 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 46.872 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 2.2752 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 2.0676 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 11.968 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 358.4600 0.4850 358.6000 ;
    END
  END top_E6END[0]
  PIN top_W1BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1253 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.4655 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 41.9268 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 224.08 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 239.1200 0.4850 239.2600 ;
    END
  END top_W1BEG[3]
  PIN top_W1BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.0304 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.991 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 27.19 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 145.48 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 1.1526 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 7.088 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 237.7600 0.4850 237.9000 ;
    END
  END top_W1BEG[2]
  PIN top_W1BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1351 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.5145 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 39.0768 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 208.88 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 236.4000 0.4850 236.5400 ;
    END
  END top_W1BEG[1]
  PIN top_W1BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2373 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.0255 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 53.1498 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 283.936 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 235.0400 0.4850 235.1800 ;
    END
  END top_W1BEG[0]
  PIN top_W2BEG[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1379 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.5285 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 26.0298 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 139.296 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 251.0200 0.4850 251.1600 ;
    END
  END top_W2BEG[7]
  PIN top_W2BEG[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.6775 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.2795 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 249.6600 0.4850 249.8000 ;
    END
  END top_W2BEG[6]
  PIN top_W2BEG[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 3.128 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 15.414 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 247.9600 0.4850 248.1000 ;
    END
  END top_W2BEG[5]
  PIN top_W2BEG[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.5409 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.4255 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 8.611 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 46.392 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 1.2168 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 6.96 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 246.6000 0.4850 246.7400 ;
    END
  END top_W2BEG[4]
  PIN top_W2BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1281 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.4795 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 31.0758 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 166.208 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 245.2400 0.4850 245.3800 ;
    END
  END top_W2BEG[3]
  PIN top_W2BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 10.9093 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 54.2675 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 38.6568 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 206.64 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 243.5400 0.4850 243.6800 ;
    END
  END top_W2BEG[2]
  PIN top_W2BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.9847 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.6445 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 50.0208 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 267.248 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 242.1800 0.4850 242.3200 ;
    END
  END top_W2BEG[1]
  PIN top_W2BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1995 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.8365 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 19.393 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 103.896 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 0.6678 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 4.032 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 240.8200 0.4850 240.9600 ;
    END
  END top_W2BEG[0]
  PIN top_W2BEGb[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1799 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.7385 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 5.7768 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 31.28 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 262.9200 0.4850 263.0600 ;
    END
  END top_W2BEGb[7]
  PIN top_W2BEGb[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.5823 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.8035 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 261.2200 0.4850 261.3600 ;
    END
  END top_W2BEGb[6]
  PIN top_W2BEGb[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1253 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.4655 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 29.0478 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 155.392 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 259.8600 0.4850 260.0000 ;
    END
  END top_W2BEGb[5]
  PIN top_W2BEGb[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.4648 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.163 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 14.4228 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 77.392 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 258.5000 0.4850 258.6400 ;
    END
  END top_W2BEGb[4]
  PIN top_W2BEGb[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.2456 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.12 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 256.8000 0.4850 256.9400 ;
    END
  END top_W2BEGb[3]
  PIN top_W2BEGb[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.1028 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 255.4400 0.4850 255.5800 ;
    END
  END top_W2BEGb[2]
  PIN top_W2BEGb[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.8288 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.983 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 28.7268 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 153.68 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 254.0800 0.4850 254.2200 ;
    END
  END top_W2BEGb[1]
  PIN top_W2BEGb[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2037 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.8575 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 21.5088 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 115.184 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 252.3800 0.4850 252.5200 ;
    END
  END top_W2BEGb[0]
  PIN top_WW4BEG[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.9041 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.2415 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 4.333 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 23.576 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 0.8508 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 5.008 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 286.3800 0.4850 286.5200 ;
    END
  END top_WW4BEG[15]
  PIN top_WW4BEG[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 7.3743 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 36.5925 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 7.0188 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 37.904 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 285.0200 0.4850 285.1600 ;
    END
  END top_WW4BEG[14]
  PIN top_WW4BEG[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 15.7323 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 78.3825 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 21.6468 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 115.92 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 283.3200 0.4850 283.4600 ;
    END
  END top_WW4BEG[13]
  PIN top_WW4BEG[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.6555 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.8805 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 5.8218 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 31.52 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 281.9600 0.4850 282.1000 ;
    END
  END top_WW4BEG[12]
  PIN top_WW4BEG[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.2716 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.132 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 280.6000 0.4850 280.7400 ;
    END
  END top_WW4BEG[11]
  PIN top_WW4BEG[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2485 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.0815 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 9.37 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 50.44 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 2.1318 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 11.84 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 278.9000 0.4850 279.0400 ;
    END
  END top_WW4BEG[10]
  PIN top_WW4BEG[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.9155 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.4695 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 277.5400 0.4850 277.6800 ;
    END
  END top_WW4BEG[9]
  PIN top_WW4BEG[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.198 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.882 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 276.1800 0.4850 276.3200 ;
    END
  END top_WW4BEG[8]
  PIN top_WW4BEG[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.0688 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.236 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 274.4800 0.4850 274.6200 ;
    END
  END top_WW4BEG[7]
  PIN top_WW4BEG[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1883 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.7805 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 12.841 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 68.952 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 3.0468 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 16.72 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 273.1200 0.4850 273.2600 ;
    END
  END top_WW4BEG[6]
  PIN top_WW4BEG[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7005 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.2235 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 58.9518 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 314.88 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 271.7600 0.4850 271.9000 ;
    END
  END top_WW4BEG[5]
  PIN top_WW4BEG[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1869 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.7735 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 15.3438 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 82.304 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 270.0600 0.4850 270.2000 ;
    END
  END top_WW4BEG[4]
  PIN top_WW4BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.5409 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.4255 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 15.649 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 83.928 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 3.5958 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 19.648 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 268.7000 0.4850 268.8400 ;
    END
  END top_WW4BEG[3]
  PIN top_WW4BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1589 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.6335 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 59.3568 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 317.04 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 267.3400 0.4850 267.4800 ;
    END
  END top_WW4BEG[2]
  PIN top_WW4BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.2456 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.12 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 265.6400 0.4850 265.7800 ;
    END
  END top_WW4BEG[1]
  PIN top_WW4BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.2256 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.02 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 264.2800 0.4850 264.4200 ;
    END
  END top_WW4BEG[0]
  PIN top_W6BEG[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.3731 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.5295 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 8.5368 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 46 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 304.0600 0.4850 304.2000 ;
    END
  END top_W6BEG[11]
  PIN top_W6BEG[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1617 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.6475 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.469 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.968 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 21.3948 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 114.576 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 302.7000 0.4850 302.8400 ;
    END
  END top_W6BEG[10]
  PIN top_W6BEG[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.702 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.402 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 301.0000 0.4850 301.1400 ;
    END
  END top_W6BEG[9]
  PIN top_W6BEG[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.0468 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.126 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 299.6400 0.4850 299.7800 ;
    END
  END top_W6BEG[8]
  PIN top_W6BEG[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.2929 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.3035 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 24.916 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 133.352 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 2.5056 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 14.304 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 298.2800 0.4850 298.4200 ;
    END
  END top_W6BEG[7]
  PIN top_W6BEG[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1647 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.6195 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 16.474 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 88.328 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 1.4544 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 9.168 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 296.5800 0.4850 296.7200 ;
    END
  END top_W6BEG[6]
  PIN top_W6BEG[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.8666 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.172 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 10.336 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 55.592 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 0.6678 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 4.032 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 295.2200 0.4850 295.3600 ;
    END
  END top_W6BEG[5]
  PIN top_W6BEG[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.0468 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.126 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 293.8600 0.4850 294.0000 ;
    END
  END top_W6BEG[4]
  PIN top_W6BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.2675 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.0585 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 24.3658 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 130.888 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 1.3356 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 8.064 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 292.1600 0.4850 292.3000 ;
    END
  END top_W6BEG[3]
  PIN top_W6BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.0468 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.126 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 290.8000 0.4850 290.9400 ;
    END
  END top_W6BEG[2]
  PIN top_W6BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.6972 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.325 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 22.939 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 122.808 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 1.2168 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 6.96 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 289.4400 0.4850 289.5800 ;
    END
  END top_W6BEG[1]
  PIN top_W6BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2065 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.8715 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 57.8868 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 309.2 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 287.7400 0.4850 287.8800 ;
    END
  END top_W6BEG[0]
  PIN top_W1END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1813 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.7455 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 2.677 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 14.744 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 2.088 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 57.1116 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 305.536 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 209.7350 239.1200 210.2200 239.2600 ;
    END
  END top_W1END[3]
  PIN top_W1END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.5246 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.462 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 3.781 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 20.632 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 2.088 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 58.7427 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 316.112 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 209.7350 237.7600 210.2200 237.9000 ;
    END
  END top_W1END[2]
  PIN top_W1END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1351 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.5145 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 31.975 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 171 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.692 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 41.8104 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 224.4 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 209.7350 236.4000 210.2200 236.5400 ;
    END
  END top_W1END[1]
  PIN top_W1END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.0059 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.8685 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 11.092 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 59.624 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.5012 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 66.9438 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 359.856 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 209.7350 235.0400 210.2200 235.1800 ;
    END
  END top_W1END[0]
  PIN top_W2MID[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.4261 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.8515 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.5724 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 33.9859 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 181.72 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.7632 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 3.7146 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 20.752 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 11.5665 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 61.3791 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 209.7350 251.0200 210.2200 251.1600 ;
    END
  END top_W2MID[7]
  PIN top_W2MID[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1575 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.6265 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.5616 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 52.3095 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 279.92 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met3  ;
    ANTENNAMAXAREACAR 73.0443 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 388.5 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.123098 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 209.7350 249.6600 210.2200 249.8000 ;
    END
  END top_W2MID[6]
  PIN top_W2MID[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1673 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.6755 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 15.925 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 85.4 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.7632 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 1.0338 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 5.984 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 18.3888 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 93.4949 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 209.7350 247.9600 210.2200 248.1000 ;
    END
  END top_W2MID[5]
  PIN top_W2MID[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.8461 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.9515 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 13.303 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 71.416 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.5616 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 1.7496 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 10.272 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 27.3414 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 144.459 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 209.7350 246.6000 210.2200 246.7400 ;
    END
  END top_W2MID[4]
  PIN top_W2MID[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.4061 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.7515 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 21.898 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 117.256 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.7632 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 12.6351 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 69.264 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 37.9254 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 203.632 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 209.7350 245.2400 210.2200 245.3800 ;
    END
  END top_W2MID[3]
  PIN top_W2MID[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.5054 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.366 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 31.579 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 168.888 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.5616 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 11.9268 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 64.08 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 61.9248 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 328.23 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 209.7350 243.5400 210.2200 243.6800 ;
    END
  END top_W2MID[2]
  PIN top_W2MID[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1799 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.7385 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.7632 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 31.6125 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 169.536 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met3  ;
    ANTENNAMAXAREACAR 43.4669 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 231.321 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.123098 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 209.7350 242.1800 210.2200 242.3200 ;
    END
  END top_W2MID[1]
  PIN top_W2MID[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.5495 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 17.4685 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 16.705 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 89.56 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.5616 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 1.7016 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 10.016 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 13.5911 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 69.835 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.207273 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 209.7350 240.8200 210.2200 240.9600 ;
    END
  END top_W2MID[0]
  PIN top_W2END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1799 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.7385 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.5652 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 38.0277 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 203.28 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met3  ;
    ANTENNAMAXAREACAR 62.6822 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 329.18 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.123098 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 209.7350 262.9200 210.2200 263.0600 ;
    END
  END top_W2END[7]
  PIN top_W2END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 8.9094 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 44.268 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 28.87 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 154.44 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.3816 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 5.8464 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 32.592 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 209.7350 261.2200 210.2200 261.3600 ;
    END
  END top_W2END[6]
  PIN top_W2END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.3897 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.6695 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.3816 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 22.2858 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 119.328 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 209.7350 259.8600 210.2200 260.0000 ;
    END
  END top_W2END[5]
  PIN top_W2END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1911 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.7945 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.3176 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 14.5416 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 78.496 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met3  ;
    ANTENNAMAXAREACAR 44.3886 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 226.638 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 209.7350 258.5000 210.2200 258.6400 ;
    END
  END top_W2END[4]
  PIN top_W2END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1239 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.4585 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.378 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 31.6108 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 169.528 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met3  ;
    ANTENNAMAXAREACAR 69.9775 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 362.981 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.230842 LAYER via3  ;
    ANTENNADIFFAREA 1.1268 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 7.9878 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 43.072 LAYER met4  ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 80.7355 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 420.991 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.230842 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 209.7350 256.8000 210.2200 256.9400 ;
    END
  END top_W2END[3]
  PIN top_W2END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.5499 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 12.4705 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.1872 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 5.6248 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 30.936 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.1268 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 5.0436 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 27.84 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 209.7350 255.4400 210.2200 255.5800 ;
    END
  END top_W2END[2]
  PIN top_W2END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 17.0973 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 85.2075 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.1304 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 18.6885 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 100.608 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 209.7350 254.0800 210.2200 254.2200 ;
    END
  END top_W2END[1]
  PIN top_W2END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.5801 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.6215 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 11.758 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 63.176 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.378 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 7.7952 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 43.456 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 19.0126 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 100.448 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 209.7350 252.3800 210.2200 252.5200 ;
    END
  END top_W2END[0]
  PIN top_WW4END[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1407 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.5425 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 37.594 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 200.968 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 1.3356 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 8.064 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 33.0385 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 176.28 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 209.7350 286.3800 210.2200 286.5200 ;
    END
  END top_WW4END[15]
  PIN top_WW4END[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.6776 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.162 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 4.84579 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 22.6889 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 209.7350 285.0200 210.2200 285.1600 ;
    END
  END top_WW4END[14]
  PIN top_WW4END[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2493 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.9765 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 7.528 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 40.616 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 3.5862 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 21.008 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 27.8568 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 150.139 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 209.7350 283.3200 210.2200 283.4600 ;
    END
  END top_WW4END[13]
  PIN top_WW4END[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1617 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.6475 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 17.995 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 96.44 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 2.9184 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 16.976 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 15.6219 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 82.3219 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 209.7350 281.9600 210.2200 282.1000 ;
    END
  END top_WW4END[12]
  PIN top_WW4END[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1813 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.7455 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 60.715 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 324.28 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.4848 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 3.056 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 3.21145 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 16.7441 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 209.7350 280.6000 210.2200 280.7400 ;
    END
  END top_WW4END[11]
  PIN top_WW4END[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.3793 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.5365 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 46.483 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 248.376 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.6678 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 4.032 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 2.58303 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 13.2525 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 209.7350 278.9000 210.2200 279.0400 ;
    END
  END top_WW4END[10]
  PIN top_WW4END[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.8432 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.99 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 1.74976 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 7.20875 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 209.7350 277.5400 210.2200 277.6800 ;
    END
  END top_WW4END[9]
  PIN top_WW4END[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1897 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.7875 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 47.4858 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 253.728 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met3  ;
    ANTENNAMAXAREACAR 66.4931 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 352.951 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.123098 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 209.7350 276.1800 210.2200 276.3200 ;
    END
  END top_WW4END[8]
  PIN top_WW4END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.4107 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.7745 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 42.6648 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 228.016 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met3  ;
    ANTENNAMAXAREACAR 61.4369 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 325.506 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.123098 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 209.7350 274.4800 210.2200 274.6200 ;
    END
  END top_WW4END[7]
  PIN top_WW4END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.0336 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.942 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 2.09293 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 8.92458 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 209.7350 273.1200 210.2200 273.2600 ;
    END
  END top_WW4END[6]
  PIN top_WW4END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1687 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.6825 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 57.364 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 306.408 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 2.0676 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 11.968 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 3.81508 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 20.7333 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 209.7350 271.7600 210.2200 271.9000 ;
    END
  END top_WW4END[5]
  PIN top_WW4END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.5083 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.2625 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 50.2548 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 268.496 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met3  ;
    ANTENNAMAXAREACAR 75.0757 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 397.107 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.123098 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 209.7350 270.0600 210.2200 270.2000 ;
    END
  END top_WW4END[4]
  PIN top_WW4END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1393 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.5355 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.1908 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 6.6124 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 35.728 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.5688 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 17.5998 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 94.336 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 209.7350 268.7000 210.2200 268.8400 ;
    END
  END top_WW4END[3]
  PIN top_WW4END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.6282 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.98 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.1249 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.136 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.5688 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 11.6316 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 62.976 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 209.7350 267.3400 210.2200 267.4800 ;
    END
  END top_WW4END[2]
  PIN top_WW4END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2261 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.9695 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.1905 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.464 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.5688 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 19.8828 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 106.512 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 209.7350 265.6400 210.2200 265.7800 ;
    END
  END top_WW4END[1]
  PIN top_WW4END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.5054 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.366 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 14.2 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 76.2 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.5688 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 20.8155 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 111.952 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 209.7350 264.2800 210.2200 264.4200 ;
    END
  END top_WW4END[0]
  PIN top_W6END[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.245 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.064 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 31.126 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 166.472 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 3.0372 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 18.08 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 32.3845 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 174.02 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 209.7350 304.0600 210.2200 304.2000 ;
    END
  END top_W6END[11]
  PIN top_W6END[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.2054 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.866 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 55.6408 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 297.688 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 3.0036 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 16.96 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 4.8497 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 26.3232 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 209.7350 302.7000 210.2200 302.8400 ;
    END
  END top_W6END[10]
  PIN top_W6END[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.198 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.882 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 3.93535 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 18.2956 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 209.7350 301.0000 210.2200 301.1400 ;
    END
  END top_W6END[9]
  PIN top_W6END[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.6061 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.9225 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 4.11919 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 19.2148 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 209.7350 299.6400 210.2200 299.7800 ;
    END
  END top_W6END[8]
  PIN top_W6END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1239 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.4585 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 43.6758 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 233.408 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met3  ;
    ANTENNAMAXAREACAR 60.6156 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 321.803 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.123098 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 209.7350 298.2800 210.2200 298.4200 ;
    END
  END top_W6END[7]
  PIN top_W6END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.9693 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.5675 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 47.203 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 252.216 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 1.0338 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 5.984 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 7.16835 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 36.4633 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 209.7350 296.5800 210.2200 296.7200 ;
    END
  END top_W6END[6]
  PIN top_W6END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7251 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.5175 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 4.40768 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 20.6572 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 209.7350 295.2200 210.2200 295.3600 ;
    END
  END top_W6END[5]
  PIN top_W6END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.4149 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.7955 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 53.299 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 284.728 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 1.6614 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 10.272 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 5.40997 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 29.3791 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 209.7350 293.8600 210.2200 294.0000 ;
    END
  END top_W6END[4]
  PIN top_W6END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.4135 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.7885 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 33.0948 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 176.976 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met3  ;
    ANTENNAMAXAREACAR 46.4193 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 246.093 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.123098 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 209.7350 292.1600 210.2200 292.3000 ;
    END
  END top_W6END[3]
  PIN top_W6END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.198 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.882 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 4.45542 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 19.9024 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 209.7350 290.8000 210.2200 290.9400 ;
    END
  END top_W6END[2]
  PIN top_W6END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.246 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.069 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.9044 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 27.3345 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 146.72 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 209.7350 289.4400 210.2200 289.5800 ;
    END
  END top_W6END[1]
  PIN top_W6END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.1908 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.2891 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.0585 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.5228 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 7.3258 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 40.008 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.7136 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 0.8508 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 5.008 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 209.7350 287.7400 210.2200 287.8800 ;
    END
  END top_W6END[0]
  PIN bot_E1BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 9.0907 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 45.1745 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 33.8778 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 181.152 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 209.7350 84.7600 210.2200 84.9000 ;
    END
  END bot_E1BEG[3]
  PIN bot_E1BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.2456 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.12 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 209.7350 83.4000 210.2200 83.5400 ;
    END
  END bot_E1BEG[2]
  PIN bot_E1BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.6165 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.8035 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 41.7666 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 223.696 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 209.7350 81.7000 210.2200 81.8400 ;
    END
  END bot_E1BEG[1]
  PIN bot_E1BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.3967 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.7045 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 7.093 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 38.296 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 2.1318 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 11.84 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 209.7350 80.3400 210.2200 80.4800 ;
    END
  END bot_E1BEG[0]
  PIN bot_E2BEG[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2674 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.176 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 2.194 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 12.168 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 24.3708 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 130.448 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 209.7350 96.6600 210.2200 96.8000 ;
    END
  END bot_E2BEG[7]
  PIN bot_E2BEG[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.2456 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.12 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 209.7350 94.9600 210.2200 95.1000 ;
    END
  END bot_E2BEG[6]
  PIN bot_E2BEG[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.0468 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.126 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 209.7350 93.6000 210.2200 93.7400 ;
    END
  END bot_E2BEG[5]
  PIN bot_E2BEG[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.1028 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 209.7350 92.2400 210.2200 92.3800 ;
    END
  END bot_E2BEG[4]
  PIN bot_E2BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1617 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.6475 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 30.2898 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 162.016 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 209.7350 90.5400 210.2200 90.6800 ;
    END
  END bot_E2BEG[3]
  PIN bot_E2BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.4158 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.918 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 13.6848 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 73.456 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 209.7350 89.1800 210.2200 89.3200 ;
    END
  END bot_E2BEG[2]
  PIN bot_E2BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 3.2652 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 16.1 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 209.7350 87.8200 210.2200 87.9600 ;
    END
  END bot_E2BEG[1]
  PIN bot_E2BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.756 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.619 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 51.1308 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 273.168 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 209.7350 86.1200 210.2200 86.2600 ;
    END
  END bot_E2BEG[0]
  PIN bot_E2BEGb[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.5908 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.793 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 10.84 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 58.28 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 1.5186 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 9.04 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 209.7350 108.2200 210.2200 108.3600 ;
    END
  END bot_E2BEGb[7]
  PIN bot_E2BEGb[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1407 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.5425 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 27.325 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 146.2 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 0.6678 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 4.032 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 209.7350 106.8600 210.2200 107.0000 ;
    END
  END bot_E2BEGb[6]
  PIN bot_E2BEGb[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2065 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.8715 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 43.3458 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 231.648 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 209.7350 105.5000 210.2200 105.6400 ;
    END
  END bot_E2BEGb[5]
  PIN bot_E2BEGb[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.0468 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.126 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 209.7350 103.8000 210.2200 103.9400 ;
    END
  END bot_E2BEGb[4]
  PIN bot_E2BEGb[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.198 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.882 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 209.7350 102.4400 210.2200 102.5800 ;
    END
  END bot_E2BEGb[3]
  PIN bot_E2BEGb[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.0037 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.9105 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 209.7350 101.0800 210.2200 101.2200 ;
    END
  END bot_E2BEGb[2]
  PIN bot_E2BEGb[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.3141 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.2915 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 16.129 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 86.488 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 1.7496 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 10.272 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 209.7350 99.3800 210.2200 99.5200 ;
    END
  END bot_E2BEGb[1]
  PIN bot_E2BEGb[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1841 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.7595 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 8.815 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 47.48 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 3.1656 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 17.824 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 209.7350 98.0200 210.2200 98.1600 ;
    END
  END bot_E2BEGb[0]
  PIN bot_EE4BEG[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.9429 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 19.4355 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 9.5028 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 51.152 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 209.7350 132.0200 210.2200 132.1600 ;
    END
  END bot_EE4BEG[15]
  PIN bot_EE4BEG[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2121 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.8995 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 12.8406 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 69.424 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 209.7350 130.3200 210.2200 130.4600 ;
    END
  END bot_EE4BEG[14]
  PIN bot_EE4BEG[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 9.0795 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 45.1185 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 15.8028 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 84.752 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 209.7350 128.9600 210.2200 129.1000 ;
    END
  END bot_EE4BEG[13]
  PIN bot_EE4BEG[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2688 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.183 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 16.4448 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 88.176 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 209.7350 127.6000 210.2200 127.7400 ;
    END
  END bot_EE4BEG[12]
  PIN bot_EE4BEG[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2219 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.7735 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 8.035 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 43.32 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 2.9184 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 16.976 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 209.7350 125.9000 210.2200 126.0400 ;
    END
  END bot_EE4BEG[11]
  PIN bot_EE4BEG[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1673 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.6755 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 16.108 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 86.376 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 1.3356 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 8.064 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 209.7350 124.5400 210.2200 124.6800 ;
    END
  END bot_EE4BEG[10]
  PIN bot_EE4BEG[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.4395 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.0895 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 209.7350 123.1800 210.2200 123.3200 ;
    END
  END bot_EE4BEG[9]
  PIN bot_EE4BEG[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1687 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.6825 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 47.4948 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 253.776 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 209.7350 121.4800 210.2200 121.6200 ;
    END
  END bot_EE4BEG[8]
  PIN bot_EE4BEG[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1883 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.7805 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 6.6498 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 35.936 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 209.7350 120.1200 210.2200 120.2600 ;
    END
  END bot_EE4BEG[7]
  PIN bot_EE4BEG[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.198 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.882 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 209.7350 118.7600 210.2200 118.9000 ;
    END
  END bot_EE4BEG[6]
  PIN bot_EE4BEG[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.5726 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.702 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 50.2488 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 268.464 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 209.7350 117.0600 210.2200 117.2000 ;
    END
  END bot_EE4BEG[5]
  PIN bot_EE4BEG[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1239 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.4585 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 21.0888 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 112.944 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 209.7350 115.7000 210.2200 115.8400 ;
    END
  END bot_EE4BEG[4]
  PIN bot_EE4BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.4871 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.3275 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 209.7350 114.3400 210.2200 114.4800 ;
    END
  END bot_EE4BEG[3]
  PIN bot_EE4BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2107 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.8925 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 38.3868 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 205.2 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 209.7350 112.6400 210.2200 112.7800 ;
    END
  END bot_EE4BEG[2]
  PIN bot_EE4BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.0468 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.126 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 209.7350 111.2800 210.2200 111.4200 ;
    END
  END bot_EE4BEG[1]
  PIN bot_EE4BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2275 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.9765 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 17.788 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 95.336 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 3.7146 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 20.752 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 209.7350 109.9200 210.2200 110.0600 ;
    END
  END bot_EE4BEG[0]
  PIN bot_E6BEG[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.0468 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.126 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 209.7350 149.7000 210.2200 149.8400 ;
    END
  END bot_E6BEG[11]
  PIN bot_E6BEG[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.0468 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.126 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 209.7350 148.0000 210.2200 148.1400 ;
    END
  END bot_E6BEG[10]
  PIN bot_E6BEG[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.616 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.919 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 46.3428 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 247.632 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 209.7350 146.6400 210.2200 146.7800 ;
    END
  END bot_E6BEG[9]
  PIN bot_E6BEG[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.198 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.882 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 209.7350 145.2800 210.2200 145.4200 ;
    END
  END bot_E6BEG[8]
  PIN bot_E6BEG[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.658 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.129 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 26.9808 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 144.368 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 209.7350 143.5800 210.2200 143.7200 ;
    END
  END bot_E6BEG[7]
  PIN bot_E6BEG[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.497 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.324 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 31.309 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 167.448 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 3.2844 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 18.928 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 209.7350 142.2200 210.2200 142.3600 ;
    END
  END bot_E6BEG[6]
  PIN bot_E6BEG[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.1462 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.623 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 209.7350 140.8600 210.2200 141.0000 ;
    END
  END bot_E6BEG[5]
  PIN bot_E6BEG[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1365 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.5215 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 14.866 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 79.752 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 1.1526 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 7.088 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 209.7350 139.1600 210.2200 139.3000 ;
    END
  END bot_E6BEG[4]
  PIN bot_E6BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7868 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.773 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 17.992 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 96.424 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 0.9696 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 6.112 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 209.7350 137.8000 210.2200 137.9400 ;
    END
  END bot_E6BEG[3]
  PIN bot_E6BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.4281 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 11.8615 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 39.8598 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 213.056 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 209.7350 136.4400 210.2200 136.5800 ;
    END
  END bot_E6BEG[2]
  PIN bot_E6BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1911 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.7945 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 19.3266 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 104.016 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 209.7350 134.7400 210.2200 134.8800 ;
    END
  END bot_E6BEG[1]
  PIN bot_E6BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1253 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.4655 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 43.726 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 233.672 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 1.1526 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 7.088 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 209.7350 133.3800 210.2200 133.5200 ;
    END
  END bot_E6BEG[0]
  PIN bot_E1END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.1872 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.6169 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 12.6875 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.378 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 28.5988 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 153.464 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 2.0736 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 3.6408 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 22.24 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 84.7600 0.4850 84.9000 ;
    END
  END bot_E1END[3]
  PIN bot_E1END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.1872 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.1547 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.2675 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.134 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 7.5568 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 41.24 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 2.0736 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 30.3456 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 162.784 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 83.4000 0.4850 83.5400 ;
    END
  END bot_E1END[2]
  PIN bot_E1END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.6104 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.891 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 27.514 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 147.208 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.6992 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 2.9826 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 16.848 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 81.7000 0.4850 81.8400 ;
    END
  END bot_E1END[1]
  PIN bot_E1END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 5.3441 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 26.3235 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.7596 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 25.7913 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 138.472 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.6992 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 14.8953 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 80.848 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 80.3400 0.4850 80.4800 ;
    END
  END bot_E1END[0]
  PIN bot_E2MID[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.3729 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.5855 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.952 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 5.544 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.7632 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 9.1404 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 50.16 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 40.1903 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 214.94 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.230842 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 96.6600 0.4850 96.8000 ;
    END
  END bot_E2MID[7]
  PIN bot_E2MID[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.9173 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.4255 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.756 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 26.0856 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 140.064 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met3  ;
    ANTENNAMAXAREACAR 53.2702 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 276.892 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 94.9600 0.4850 95.1000 ;
    END
  END bot_E2MID[6]
  PIN bot_E2MID[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1435 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.5565 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.7632 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 6.8778 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 37.152 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met3  ;
    ANTENNAMAXAREACAR 17.5617 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 88.1434 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.153401 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 93.6000 0.4850 93.7400 ;
    END
  END bot_E2MID[5]
  PIN bot_E2MID[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1631 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.6545 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 24.5758 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 132.008 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.5688 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 5.4738 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 29.664 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 60.471 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 320.331 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 92.2400 0.4850 92.3800 ;
    END
  END bot_E2MID[4]
  PIN bot_E2MID[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.1285 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.3635 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.7632 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 56.7606 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 303.184 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met3  ;
    ANTENNAMAXAREACAR 77.4059 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 411.757 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.123098 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 90.5400 0.4850 90.6800 ;
    END
  END bot_E2MID[3]
  PIN bot_E2MID[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1645 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.6615 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 6.838 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 36.936 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.5688 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 25.4352 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 137.536 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 36.8906 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 197.572 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 89.1800 0.4850 89.3200 ;
    END
  END bot_E2MID[2]
  PIN bot_E2MID[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.953 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.604 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.7632 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 20.3826 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 109.648 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met3  ;
    ANTENNAMAXAREACAR 28.9534 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 153.719 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.123098 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 87.8200 0.4850 87.9600 ;
    END
  END bot_E2MID[1]
  PIN bot_E2MID[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1659 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.6685 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.7596 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 27.3438 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 146.304 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met3  ;
    ANTENNAMAXAREACAR 51.4991 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 268.185 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.123098 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 86.1200 0.4850 86.2600 ;
    END
  END bot_E2MID[0]
  PIN bot_E2END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 6.8283 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 33.8625 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 31.3768 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 168.28 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.954 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 2.0034 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 12.096 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 108.2200 0.4850 108.3600 ;
    END
  END bot_E2END[7]
  PIN bot_E2END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1659 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.6685 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.262 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.864 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.1448 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 25.0068 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 133.84 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 106.8600 0.4850 107.0000 ;
    END
  END bot_E2END[6]
  PIN bot_E2END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.7113 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.2775 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 22.981 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 123.032 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.1448 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 1.5186 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 9.04 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 105.5000 0.4850 105.6400 ;
    END
  END bot_E2END[5]
  PIN bot_E2END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 7.3379 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 36.4105 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.9468 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 8.2515 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 44.944 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 103.8000 0.4850 103.9400 ;
    END
  END bot_E2END[4]
  PIN bot_E2END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.8489 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.9655 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 20.5316 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 109.96 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via3  ;
    ANTENNADIFFAREA 1.5156 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 3.3486 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 18.8 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 102.4400 0.4850 102.5800 ;
    END
  END bot_E2END[3]
  PIN bot_E2END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.4779 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.1105 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.332 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 22.8858 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 122.528 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 101.0800 0.4850 101.2200 ;
    END
  END bot_E2END[2]
  PIN bot_E2END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.1872 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.0881 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.0435 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.1872 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.331 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.232 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.756 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 5.0598 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 27.456 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 99.3800 0.4850 99.5200 ;
    END
  END bot_E2END[1]
  PIN bot_E2END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1841 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.7595 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 11.296 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 60.712 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.7632 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 5.9586 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 32.72 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 98.0200 0.4850 98.1600 ;
    END
  END bot_E2END[0]
  PIN bot_EE4END[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1617 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.6475 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 10.8798 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 58.496 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met3  ;
    ANTENNAMAXAREACAR 21.0687 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 109.395 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.123098 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 132.0200 0.4850 132.1600 ;
    END
  END bot_EE4END[15]
  PIN bot_EE4END[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.4956 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.252 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 4.53657 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 21.1428 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 130.3200 0.4850 130.4600 ;
    END
  END bot_EE4END[14]
  PIN bot_EE4END[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.5661 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.5515 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 54.1668 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 289.36 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met3  ;
    ANTENNAMAXAREACAR 75.278 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 399.875 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.123098 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 128.9600 0.4850 129.1000 ;
    END
  END bot_EE4END[13]
  PIN bot_EE4END[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.178 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.782 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 12.1411 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 59.3246 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 127.6000 0.4850 127.7400 ;
    END
  END bot_EE4END[12]
  PIN bot_EE4END[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1589 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.6335 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 30.8278 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 165.352 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 1.5186 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 9.04 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 24.5666 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 131.098 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 125.9000 0.4850 126.0400 ;
    END
  END bot_EE4END[11]
  PIN bot_EE4END[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1393 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.5355 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 10.516 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 56.552 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 1.3356 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 8.064 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 49.2917 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 262.411 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 124.5400 0.4850 124.6800 ;
    END
  END bot_EE4END[10]
  PIN bot_EE4END[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.3112 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.33 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 1.2064 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 3.49832 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 123.1800 0.4850 123.3200 ;
    END
  END bot_EE4END[9]
  PIN bot_EE4END[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1379 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.5285 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 24.607 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 131.704 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 1.8846 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 10.992 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 26.0648 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 139.752 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 121.4800 0.4850 121.6200 ;
    END
  END bot_EE4END[8]
  PIN bot_EE4END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.2647 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.0445 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 52.9248 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 282.736 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met3  ;
    ANTENNAMAXAREACAR 74.2294 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 394.074 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.123098 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 120.1200 0.4850 120.2600 ;
    END
  END bot_EE4END[7]
  PIN bot_EE4END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.3752 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.715 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 11.8938 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 63.904 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met3  ;
    ANTENNAMAXAREACAR 19.6853 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 102.933 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.123098 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 118.7600 0.4850 118.9000 ;
    END
  END bot_EE4END[6]
  PIN bot_EE4END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.1172 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.425 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 37.495 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 200.44 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 2.0676 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 11.968 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 17.1258 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 91.0276 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 117.0600 0.4850 117.2000 ;
    END
  END bot_EE4END[5]
  PIN bot_EE4END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1827 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.7525 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 20.341 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 108.952 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 1.9488 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 10.864 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 3.87111 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 20.1751 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 115.7000 0.4850 115.8400 ;
    END
  END bot_EE4END[4]
  PIN bot_EE4END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.8638 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.158 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 7.9468 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 43.32 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.378 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 1.9488 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 10.864 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 114.3400 0.4850 114.4800 ;
    END
  END bot_EE4END[3]
  PIN bot_EE4END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.6781 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.1115 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 13.21 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 70.92 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.5652 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 30.7923 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 165.632 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 112.6400 0.4850 112.7800 ;
    END
  END bot_EE4END[2]
  PIN bot_EE4END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 6.2795 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 31.1185 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.5724 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 4.9587 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 26.912 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 111.2800 0.4850 111.4200 ;
    END
  END bot_EE4END[1]
  PIN bot_EE4END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.3001 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.2215 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 5.251 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 28.472 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.5724 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 26.0181 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 140.64 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 109.9200 0.4850 110.0600 ;
    END
  END bot_EE4END[0]
  PIN bot_E6END[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1603 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.6405 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 13.1808 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 70.768 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met3  ;
    ANTENNAMAXAREACAR 22.1568 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 115.173 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.123098 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 149.7000 0.4850 149.8400 ;
    END
  END bot_E6END[11]
  PIN bot_E6END[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.3202 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.44 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 52.3476 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 280.128 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met3  ;
    ANTENNAMAXAREACAR 73.584 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 391.222 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.123098 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 148.0000 0.4850 148.1400 ;
    END
  END bot_E6END[10]
  PIN bot_E6END[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1589 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.6335 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 35.1678 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 188.032 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met3  ;
    ANTENNAMAXAREACAR 48.8489 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 259.291 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.123098 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 146.6400 0.4850 146.7800 ;
    END
  END bot_E6END[9]
  PIN bot_E6END[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2247 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.9625 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 12.4428 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 66.832 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met3  ;
    ANTENNAMAXAREACAR 18.5014 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 97.2606 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.123098 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 145.2800 0.4850 145.4200 ;
    END
  END bot_E6END[8]
  PIN bot_E6END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.252 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.099 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 53.4708 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 285.648 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met3  ;
    ANTENNAMAXAREACAR 75.883 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 402.587 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.123098 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 143.5800 0.4850 143.7200 ;
    END
  END bot_E6END[7]
  PIN bot_E6END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7322 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.5 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 38.9388 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 208.144 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met3  ;
    ANTENNAMAXAREACAR 53.762 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 285.459 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.123098 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 142.2200 0.4850 142.3600 ;
    END
  END bot_E6END[6]
  PIN bot_E6END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.6052 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.8 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 5.14471 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 23.4875 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 140.8600 0.4850 141.0000 ;
    END
  END bot_E6END[5]
  PIN bot_E6END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.9464 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.506 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 7.00626 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 32.4976 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 139.1600 0.4850 139.3000 ;
    END
  END bot_E6END[4]
  PIN bot_E6END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.9709 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.6935 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 28.045 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 150.04 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 2.3694 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 14.048 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 5.29791 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 29.0707 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 137.8000 0.4850 137.9400 ;
    END
  END bot_E6END[3]
  PIN bot_E6END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1827 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.7525 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 16.1688 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 86.704 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met3  ;
    ANTENNAMAXAREACAR 22.6824 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 119.838 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.123098 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 136.4400 0.4850 136.5800 ;
    END
  END bot_E6END[2]
  PIN bot_E6END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.5036 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 22.239 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.378 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 2.2288 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 12.824 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 2.2644 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 5.0598 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 27.456 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 134.7400 0.4850 134.8800 ;
    END
  END bot_E6END[1]
  PIN bot_E6END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 15.5979 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 77.7105 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 2.268 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 24.3456 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 131.24 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 133.3800 0.4850 133.5200 ;
    END
  END bot_E6END[0]
  PIN bot_W1BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.3755 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.7165 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.1905 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.464 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 11.6076 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 62.848 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 14.0400 0.4850 14.1800 ;
    END
  END bot_W1BEG[3]
  PIN bot_W1BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 7.0422 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 34.867 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 12.6800 0.4850 12.8200 ;
    END
  END bot_W1BEG[2]
  PIN bot_W1BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1337 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.5075 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 6.8328 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 36.912 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 11.3200 0.4850 11.4600 ;
    END
  END bot_W1BEG[1]
  PIN bot_W1BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1533 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.6055 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.262 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.864 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 27.3858 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 146.528 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 9.9600 0.4850 10.1000 ;
    END
  END bot_W1BEG[0]
  PIN bot_W2BEG[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1365 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.5215 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 28.9998 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 155.136 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 25.9400 0.4850 26.0800 ;
    END
  END bot_W2BEG[7]
  PIN bot_W2BEG[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 16.4848 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 82.145 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 10.7448 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 57.776 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 24.5800 0.4850 24.7200 ;
    END
  END bot_W2BEG[6]
  PIN bot_W2BEG[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 10.9666 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 54.607 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 22.8800 0.4850 23.0200 ;
    END
  END bot_W2BEG[5]
  PIN bot_W2BEG[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.7188 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.486 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 21.5200 0.4850 21.6600 ;
    END
  END bot_W2BEG[4]
  PIN bot_W2BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1295 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.4865 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 11.83 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 63.56 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 1.5828 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 8.912 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 20.1600 0.4850 20.3000 ;
    END
  END bot_W2BEG[3]
  PIN bot_W2BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.0925 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.1835 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 9.691 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 52.152 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 7.4388 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 40.144 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 18.4600 0.4850 18.6000 ;
    END
  END bot_W2BEG[2]
  PIN bot_W2BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1281 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.4795 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 19.1598 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 102.656 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 17.1000 0.4850 17.2400 ;
    END
  END bot_W2BEG[1]
  PIN bot_W2BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.4224 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 11.886 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 15.7400 0.4850 15.8800 ;
    END
  END bot_W2BEG[0]
  PIN bot_W2BEGb[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7999 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.7205 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 9.4548 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 50.896 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 37.8400 0.4850 37.9800 ;
    END
  END bot_W2BEGb[7]
  PIN bot_W2BEGb[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1603 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.6405 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 10.6968 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 57.52 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 36.1400 0.4850 36.2800 ;
    END
  END bot_W2BEGb[6]
  PIN bot_W2BEGb[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.4395 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.0895 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 34.7800 0.4850 34.9200 ;
    END
  END bot_W2BEGb[5]
  PIN bot_W2BEGb[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1995 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.8365 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 8.287 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 44.664 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 1.2168 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 6.96 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 33.4200 0.4850 33.5600 ;
    END
  END bot_W2BEGb[4]
  PIN bot_W2BEGb[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2443 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.0605 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 28.2678 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 151.232 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 31.7200 0.4850 31.8600 ;
    END
  END bot_W2BEGb[3]
  PIN bot_W2BEGb[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.6501 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.9715 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 18.6078 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 99.712 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 30.3600 0.4850 30.5000 ;
    END
  END bot_W2BEGb[2]
  PIN bot_W2BEGb[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.1462 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.623 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 29.0000 0.4850 29.1400 ;
    END
  END bot_W2BEGb[1]
  PIN bot_W2BEGb[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.0135 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.9595 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 27.3000 0.4850 27.4400 ;
    END
  END bot_W2BEGb[0]
  PIN bot_WW4BEG[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1393 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.5355 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.676 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 4.072 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 8.7198 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 46.976 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 61.3000 0.4850 61.4400 ;
    END
  END bot_WW4BEG[15]
  PIN bot_WW4BEG[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1589 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.6335 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.469 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.968 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 23.2248 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 124.336 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 59.9400 0.4850 60.0800 ;
    END
  END bot_WW4BEG[14]
  PIN bot_WW4BEG[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2261 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.9695 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 24.544 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 131.368 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 2.79 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 17.232 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 58.2400 0.4850 58.3800 ;
    END
  END bot_WW4BEG[13]
  PIN bot_WW4BEG[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1603 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.6405 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 5.182 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 28.104 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 18.6018 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 99.68 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 56.8800 0.4850 57.0200 ;
    END
  END bot_WW4BEG[12]
  PIN bot_WW4BEG[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1799 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.7385 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 40.921 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 218.712 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 0.6678 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 4.032 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 55.5200 0.4850 55.6600 ;
    END
  END bot_WW4BEG[11]
  PIN bot_WW4BEG[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.4155 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.7535 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 39.3978 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 210.592 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 53.8200 0.4850 53.9600 ;
    END
  END bot_WW4BEG[10]
  PIN bot_WW4BEG[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1253 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.4655 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 47.059 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 251.448 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 0.6678 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 4.032 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 52.4600 0.4850 52.6000 ;
    END
  END bot_WW4BEG[9]
  PIN bot_WW4BEG[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.2456 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.12 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 51.1000 0.4850 51.2400 ;
    END
  END bot_WW4BEG[8]
  PIN bot_WW4BEG[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.5116 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.45 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 49.4000 0.4850 49.5400 ;
    END
  END bot_WW4BEG[7]
  PIN bot_WW4BEG[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.0384 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.084 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 48.0400 0.4850 48.1800 ;
    END
  END bot_WW4BEG[6]
  PIN bot_WW4BEG[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1365 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.5215 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 3.7068 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 20.24 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 46.6800 0.4850 46.8200 ;
    END
  END bot_WW4BEG[5]
  PIN bot_WW4BEG[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1883 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.7805 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 11.527 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 61.944 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 1.9392 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 12.224 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 44.9800 0.4850 45.1200 ;
    END
  END bot_WW4BEG[4]
  PIN bot_WW4BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.5991 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.8875 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 43.6200 0.4850 43.7600 ;
    END
  END bot_WW4BEG[3]
  PIN bot_WW4BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.1938 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.861 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 42.2600 0.4850 42.4000 ;
    END
  END bot_WW4BEG[2]
  PIN bot_WW4BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1673 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.6755 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 30.2898 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 162.016 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 40.5600 0.4850 40.7000 ;
    END
  END bot_WW4BEG[1]
  PIN bot_WW4BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.6167 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.9225 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 11.785 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 63.32 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 1.7658 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 9.888 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 39.2000 0.4850 39.3400 ;
    END
  END bot_WW4BEG[0]
  PIN bot_W6BEG[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2436 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.057 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 10.885 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 58.52 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 12.2514 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 66.752 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 78.9800 0.4850 79.1200 ;
    END
  END bot_W6BEG[11]
  PIN bot_W6BEG[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1463 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.5705 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 33.7 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 180.2 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 1.7016 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 10.016 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 77.6200 0.4850 77.7600 ;
    END
  END bot_W6BEG[10]
  PIN bot_W6BEG[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.3673 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.5575 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 20.476 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 109.672 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 0.9696 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 6.112 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 75.9200 0.4850 76.0600 ;
    END
  END bot_W6BEG[9]
  PIN bot_W6BEG[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1617 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.6475 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 12.6708 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 68.048 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 74.5600 0.4850 74.7000 ;
    END
  END bot_W6BEG[8]
  PIN bot_W6BEG[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.6068 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.926 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 73.2000 0.4850 73.3400 ;
    END
  END bot_W6BEG[7]
  PIN bot_W6BEG[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.8428 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.053 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 14.656 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 78.632 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 1.6308 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 9.168 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 71.5000 0.4850 71.6400 ;
    END
  END bot_W6BEG[6]
  PIN bot_W6BEG[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.3015 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.2285 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 57.3348 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 306.256 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 70.1400 0.4850 70.2800 ;
    END
  END bot_W6BEG[5]
  PIN bot_W6BEG[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2023 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.8505 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 10.2378 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 55.072 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 68.7800 0.4850 68.9200 ;
    END
  END bot_W6BEG[4]
  PIN bot_W6BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1841 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.7595 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 10.0548 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 54.096 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 67.0800 0.4850 67.2200 ;
    END
  END bot_W6BEG[3]
  PIN bot_W6BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.5719 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.6985 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 28.3128 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 151.472 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 65.7200 0.4850 65.8600 ;
    END
  END bot_W6BEG[2]
  PIN bot_W6BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.3645 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.5435 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 8.8098 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 47.456 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 64.3600 0.4850 64.5000 ;
    END
  END bot_W6BEG[1]
  PIN bot_W6BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.0468 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.126 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 62.6600 0.4850 62.8000 ;
    END
  END bot_W6BEG[0]
  PIN bot_W1END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.5192 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 21.493 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 105.777 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via2  ;
    ANTENNADIFFAREA 2.088 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 6.7275 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 36.816 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 209.7350 14.0400 210.2200 14.1800 ;
    END
  END bot_W1END[3]
  PIN bot_W1END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.378 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 6.9022 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 33.481 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via2  ;
    ANTENNADIFFAREA 0.5688 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 3.2788 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 18.424 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 2.088 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 36.0186 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 193.04 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 209.7350 12.6800 210.2200 12.8200 ;
    END
  END bot_W1END[2]
  PIN bot_W1END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.1872 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.3681 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.4435 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.9432 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 25.3072 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 135.424 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.692 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 7.3038 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 39.424 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 209.7350 11.3200 210.2200 11.4600 ;
    END
  END bot_W1END[1]
  PIN bot_W1END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3744 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 6.7001 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 32.7495 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.3744 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.1905 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.464 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.5012 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 51.3285 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 274.688 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 209.7350 9.9600 210.2200 10.1000 ;
    END
  END bot_W1END[0]
  PIN bot_W2MID[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.0932 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.187 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 43.2907 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 231.824 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met3  ;
    ANTENNAMAXAREACAR 63.1139 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 334.429 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.261145 LAYER via3  ;
    ANTENNADIFFAREA 0.7632 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 40.1088 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 214.384 LAYER met4  ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 117.133 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 623.162 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.261145 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 209.7350 25.9400 210.2200 26.0800 ;
    END
  END bot_W2MID[7]
  PIN bot_W2MID[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 11.2035 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 55.3945 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 17.3284 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 84.567 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.123098 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.331 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.232 LAYER met3  ;
    ANTENNAGATEAREA 0.7425 LAYER met3  ;
    ANTENNAMAXAREACAR 17.7741 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 87.5731 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via3  ;
    ANTENNADIFFAREA 0.5616 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 32.3826 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 173.648 LAYER met4  ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 61.3871 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 321.442 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 209.7350 24.5800 210.2200 24.7200 ;
    END
  END bot_W2MID[6]
  PIN bot_W2MID[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.5988 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.833 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 50.62 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 270.44 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.7632 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 16.2807 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 87.296 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 37.3883 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 198.308 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 209.7350 22.8800 210.2200 23.0200 ;
    END
  END bot_W2MID[5]
  PIN bot_W2MID[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.369 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.566 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 34.0927 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 182.768 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met3  ;
    ANTENNAMAXAREACAR 52.6154 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 277.807 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.261145 LAYER via3  ;
    ANTENNADIFFAREA 0.5616 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 28.2618 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 151.2 LAYER met4  ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 90.6784 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 481.443 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.261145 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 209.7350 21.5200 210.2200 21.6600 ;
    END
  END bot_W2MID[4]
  PIN bot_W2MID[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1771 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.7245 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 28.8971 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 155.04 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met3  ;
    ANTENNAMAXAREACAR 40.7714 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 216.606 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via3  ;
    ANTENNADIFFAREA 0.7632 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 34.4904 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 185.36 LAYER met4  ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 87.2232 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 466.249 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 209.7350 20.1600 210.2200 20.3000 ;
    END
  END bot_W2MID[3]
  PIN bot_W2MID[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2443 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.0605 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 35.1988 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 188.664 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met3  ;
    ANTENNAMAXAREACAR 50.7205 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 269.075 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.230842 LAYER via3  ;
    ANTENNADIFFAREA 0.5616 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 29.0808 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 155.568 LAYER met4  ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 89.8866 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 478.594 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.230842 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 209.7350 18.4600 210.2200 18.6000 ;
    END
  END bot_W2MID[2]
  PIN bot_W2MID[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1785 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.7315 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 42.85 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 229 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.7632 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 18.5715 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 99.984 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 36.2804 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 193.002 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 209.7350 17.1000 210.2200 17.2400 ;
    END
  END bot_W2MID[1]
  PIN bot_W2MID[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1981 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.8295 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 60.8663 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 325.552 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via3  ;
    ANTENNADIFFAREA 0.7488 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 37.2756 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 199.744 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 51.2947 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 274.041 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 209.7350 15.7400 210.2200 15.8800 ;
    END
  END bot_W2MID[0]
  PIN bot_W2END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.3636 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.657 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.5652 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 26.0598 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 139.456 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met3  ;
    ANTENNAMAXAREACAR 66.0521 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 339.737 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.153401 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 209.7350 37.8400 210.2200 37.9800 ;
    END
  END bot_W2END[7]
  PIN bot_W2END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2457 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.0675 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 4.492 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 24.424 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.3816 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 34.7058 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 185.568 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 209.7350 36.1400 210.2200 36.2800 ;
    END
  END bot_W2END[6]
  PIN bot_W2END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1799 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.7385 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 3.919 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 21.368 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.3816 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 8.6394 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 47.488 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 209.7350 34.7800 210.2200 34.9200 ;
    END
  END bot_W2END[5]
  PIN bot_W2END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2297 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.7945 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.5688 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 39.0988 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 208.984 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.3176 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 1.8846 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 10.992 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 21.3026 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 112.292 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.207273 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 209.7350 33.4200 210.2200 33.5600 ;
    END
  END bot_W2END[4]
  PIN bot_W2END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.4621 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.0315 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 39.2644 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 209.872 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met3  ;
    ANTENNAMAXAREACAR 55.0057 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 291.811 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via3  ;
    ANTENNADIFFAREA 1.1268 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 21.6966 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 116.656 LAYER met4  ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 84.2267 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 448.924 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 209.7350 31.7200 210.2200 31.8600 ;
    END
  END bot_W2END[3]
  PIN bot_W2END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2953 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.2005 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 13.324 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 71.528 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.1268 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 0.6678 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 4.032 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 209.7350 30.3600 210.2200 30.5000 ;
    END
  END bot_W2END[2]
  PIN bot_W2END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.8404 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 13.923 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.1304 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 34.6578 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 185.312 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 209.7350 29.0000 210.2200 29.1400 ;
    END
  END bot_W2END[1]
  PIN bot_W2END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2926 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.302 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.378 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 33.5988 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 179.664 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met3  ;
    ANTENNAMAXAREACAR 59.1605 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 309.56 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.153401 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 209.7350 27.3000 210.2200 27.4400 ;
    END
  END bot_W2END[0]
  PIN bot_WW4END[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.413 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.904 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 19.0218 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 101.92 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met3  ;
    ANTENNAMAXAREACAR 30.03 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 157.857 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.123098 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 209.7350 61.3000 210.2200 61.4400 ;
    END
  END bot_WW4END[15]
  PIN bot_WW4END[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.5381 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.4115 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 17.7348 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 95.056 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met3  ;
    ANTENNAMAXAREACAR 27.1692 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 142.975 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.123098 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 209.7350 59.9400 210.2200 60.0800 ;
    END
  END bot_WW4END[14]
  PIN bot_WW4END[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.8041 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.7415 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 5.2248 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 28.336 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met3  ;
    ANTENNAMAXAREACAR 10.7705 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 55.4828 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.123098 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 209.7350 58.2400 210.2200 58.3800 ;
    END
  END bot_WW4END[13]
  PIN bot_WW4END[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2571 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.9975 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 7.99 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 43.08 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 4.3518 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 23.68 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 73.0808 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 389.044 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 209.7350 56.8800 210.2200 57.0200 ;
    END
  END bot_WW4END[12]
  PIN bot_WW4END[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1267 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.4725 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 25.924 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 138.728 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 2.4978 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 13.792 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 51.3304 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 272.5 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 209.7350 55.5200 210.2200 55.6600 ;
    END
  END bot_WW4END[11]
  PIN bot_WW4END[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.6916 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.297 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 25.672 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 137.384 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 2.3934 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 14.176 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 23.6481 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 122.292 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 209.7350 53.8200 210.2200 53.9600 ;
    END
  END bot_WW4END[10]
  PIN bot_WW4END[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.399 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.834 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 37.0548 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 198.096 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met3  ;
    ANTENNAMAXAREACAR 54.8352 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 289.82 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.123098 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 209.7350 52.4600 210.2200 52.6000 ;
    END
  END bot_WW4END[9]
  PIN bot_WW4END[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2009 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.8435 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 30.343 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 162.296 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 2.1318 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 11.84 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 5.92741 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 30.6316 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 209.7350 51.1000 210.2200 51.2400 ;
    END
  END bot_WW4END[8]
  PIN bot_WW4END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1239 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.4585 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 45.3288 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 242.224 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met3  ;
    ANTENNAMAXAREACAR 64.7212 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 343.123 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.123098 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 209.7350 49.4000 210.2200 49.5400 ;
    END
  END bot_WW4END[7]
  PIN bot_WW4END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7425 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.4335 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 53.1948 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 284.176 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met3  ;
    ANTENNAMAXAREACAR 74.1782 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 393.939 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.123098 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 209.7350 48.0400 210.2200 48.1800 ;
    END
  END bot_WW4END[6]
  PIN bot_WW4END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1701 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.6895 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 23.0718 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 123.52 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met3  ;
    ANTENNAMAXAREACAR 33.4234 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 176.484 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.123098 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 209.7350 46.6800 210.2200 46.8200 ;
    END
  END bot_WW4END[5]
  PIN bot_WW4END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.6557 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.9995 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 33.9666 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 182.096 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met3  ;
    ANTENNAMAXAREACAR 49.658 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 263.34 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.123098 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 209.7350 44.9800 210.2200 45.1200 ;
    END
  END bot_WW4END[4]
  PIN bot_WW4END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.5278 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.478 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 18.061 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 96.792 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.5688 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 10.0185 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 54.368 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 209.7350 43.6200 210.2200 43.7600 ;
    END
  END bot_WW4END[3]
  PIN bot_WW4END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.1247 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.3445 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.1908 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 28.7344 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 153.712 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.5688 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 20.2185 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 108.768 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 209.7350 42.2600 210.2200 42.4000 ;
    END
  END bot_WW4END[2]
  PIN bot_WW4END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.3701 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.5715 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 13.807 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 74.104 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.5688 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 9.2046 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 50.032 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 209.7350 40.5600 210.2200 40.7000 ;
    END
  END bot_WW4END[1]
  PIN bot_WW4END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1589 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.6335 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.1905 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.464 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.5688 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 38.9148 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 208.016 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 209.7350 39.2000 210.2200 39.3400 ;
    END
  END bot_WW4END[0]
  PIN bot_W6END[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1407 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.5425 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 21.0438 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 112.704 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met3  ;
    ANTENNAMAXAREACAR 31.7539 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 167.385 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.123098 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 209.7350 78.9800 210.2200 79.1200 ;
    END
  END bot_W6END[11]
  PIN bot_W6END[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1463 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.5705 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 6.586 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 35.592 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 1.2168 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 6.96 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 65.5883 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 348.853 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 209.7350 77.6200 210.2200 77.7600 ;
    END
  END bot_W6END[10]
  PIN bot_W6END[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.2073 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.7575 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 28.363 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 151.736 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 2.6166 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 14.896 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 38.4481 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 204.431 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 209.7350 75.9200 210.2200 76.0600 ;
    END
  END bot_W6END[9]
  PIN bot_W6END[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.6061 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.9225 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 3.83636 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 17.8007 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 209.7350 74.5600 210.2200 74.7000 ;
    END
  END bot_W6END[8]
  PIN bot_W6END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.0384 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.084 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 3.72283 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 17.1832 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 209.7350 73.2000 210.2200 73.3400 ;
    END
  END bot_W6END[7]
  PIN bot_W6END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1631 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.6545 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 53.0088 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 283.184 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met3  ;
    ANTENNAMAXAREACAR 72.6415 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 386.263 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.123098 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 209.7350 71.5000 210.2200 71.6400 ;
    END
  END bot_W6END[6]
  PIN bot_W6END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1239 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.4585 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 11.896 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 63.912 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 2.0034 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 12.096 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 8.19798 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 43.0128 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 209.7350 70.1400 210.2200 70.2800 ;
    END
  END bot_W6END[5]
  PIN bot_W6END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1897 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.7875 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 18.361 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 98.392 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.9696 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 6.112 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 19.8447 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 106.168 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 209.7350 68.7800 210.2200 68.9200 ;
    END
  END bot_W6END[4]
  PIN bot_W6END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.9315 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.3785 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 5.827 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 31.544 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 1.3356 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 8.064 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 60.9033 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 324.393 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 209.7350 67.0800 210.2200 67.2200 ;
    END
  END bot_W6END[3]
  PIN bot_W6END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1883 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.7805 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 51.775 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 276.6 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 2.0676 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 11.968 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 6.67354 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 35.029 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 209.7350 65.7200 210.2200 65.8600 ;
    END
  END bot_W6END[2]
  PIN bot_W6END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 9.2125 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 45.7835 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.1872 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 7.9069 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 42.632 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.8972 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 1.8846 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 10.992 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 209.7350 64.3600 210.2200 64.5000 ;
    END
  END bot_W6END[1]
  PIN bot_W6END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1869 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.7735 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 2.836 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 15.592 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.7064 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 7.3038 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 39.424 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 209.7350 62.6600 210.2200 62.8000 ;
    END
  END bot_W6END[0]
  PIN bot_S1BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.27625 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.325 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.1894 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 5.8695 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 5.0777 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 25.2175 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.883 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 5.176 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 17.7828 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 95.312 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 84.3250 0.0000 84.4950 0.3300 ;
    END
  END bot_S1BEG[3]
  PIN bot_S1BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.62305 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.733 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 4.002 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 19.9325 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 3.5824 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 17.794 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 82.9450 0.0000 83.1150 0.3300 ;
    END
  END bot_S1BEG[2]
  PIN bot_S1BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.81685 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.961 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 8.0256 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 40.0505 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 8.3312 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 41.538 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 81.5650 0.0000 81.7350 0.3300 ;
    END
  END bot_S1BEG[1]
  PIN bot_S1BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.62305 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.733 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.3004 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.4245 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 11.344 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 56.602 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 80.1850 0.0000 80.3550 0.3300 ;
    END
  END bot_S1BEG[0]
  PIN bot_S2BEG[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.10285 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.121 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.0832 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.1049 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.4585 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.1905 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.464 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 52.7358 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 281.728 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 105.9450 0.0000 106.1150 0.3300 ;
    END
  END bot_S2BEG[7]
  PIN bot_S2BEG[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.16065 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.189 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.6224 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 3.0345 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.1751 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.6475 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.331 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.232 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 33.6408 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 179.888 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 104.5650 0.0000 104.7350 0.3300 ;
    END
  END bot_S2BEG[6]
  PIN bot_S2BEG[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.68085 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.801 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.524 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 7.5425 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 2.9973 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.8155 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.1905 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.464 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 39.9018 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 213.28 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 103.1850 0.0000 103.3550 0.3300 ;
    END
  END bot_S2BEG[5]
  PIN bot_S2BEG[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.73865 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.869 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.3648 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.7465 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 7.5696 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 37.73 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 102.2650 0.0000 102.4350 0.3300 ;
    END
  END bot_S2BEG[4]
  PIN bot_S2BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.73865 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.869 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.1716 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.7805 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.3592 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.678 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 100.8850 0.0000 101.0550 0.3300 ;
    END
  END bot_S2BEG[3]
  PIN bot_S2BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.73865 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.869 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.0832 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 6.6148 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 32.956 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 99.5050 0.0000 99.6750 0.3300 ;
    END
  END bot_S2BEG[2]
  PIN bot_S2BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.73865 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.869 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.0832 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.1212 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.488 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 98.1250 0.0000 98.2950 0.3300 ;
    END
  END bot_S2BEG[1]
  PIN bot_S2BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.73865 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.869 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.8632 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 4.2385 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.1212 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.488 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 96.7450 0.0000 96.9150 0.3300 ;
    END
  END bot_S2BEG[0]
  PIN bot_S2BEGb[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.79645 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.937 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.9104 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 9.4745 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 3.4579 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 17.1185 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.711 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 9.592 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 41.6208 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 222.448 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 95.3650 0.0000 95.5350 0.3300 ;
    END
  END bot_S2BEGb[7]
  PIN bot_S2BEGb[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.10285 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.121 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.0832 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 21.9308 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 109.536 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 93.9850 0.0000 94.1550 0.3300 ;
    END
  END bot_S2BEGb[6]
  PIN bot_S2BEGb[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.54785 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.821 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.4292 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 2.0685 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 11.8816 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 59.29 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 92.6050 0.0000 92.7750 0.3300 ;
    END
  END bot_S2BEGb[5]
  PIN bot_S2BEGb[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.73865 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.869 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.6224 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 3.0345 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.6439 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.0485 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.1249 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.136 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 38.8998 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 207.936 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 91.2250 0.0000 91.3950 0.3300 ;
    END
  END bot_S2BEGb[4]
  PIN bot_S2BEGb[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.16065 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.189 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 4.4192 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 22.0185 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.1075 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.4655 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.1249 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.136 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 29.2638 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 156.544 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 89.8450 0.0000 90.0150 0.3300 ;
    END
  END bot_S2BEGb[3]
  PIN bot_S2BEGb[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.27625 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.325 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.9104 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 9.4745 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 17.9476 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 89.502 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 88.4650 0.0000 88.6350 0.3300 ;
    END
  END bot_S2BEGb[2]
  PIN bot_S2BEGb[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.10285 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.121 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.88 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 4.3225 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 15.285 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 76.307 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 87.0850 0.0000 87.2550 0.3300 ;
    END
  END bot_S2BEGb[1]
  PIN bot_S2BEGb[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.73865 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.869 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.1716 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.7805 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 18.1368 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 90.566 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 85.7050 0.0000 85.8750 0.3300 ;
    END
  END bot_S2BEGb[0]
  PIN bot_S4BEG[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.39185 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.461 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 13.053 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 65.1875 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 4.568 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 22.722 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 127.5650 0.0000 127.7350 0.3300 ;
    END
  END bot_S4BEG[15]
  PIN bot_S4BEG[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.33405 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.393 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.992 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 4.8825 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 18.1256 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 90.51 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 126.1850 0.0000 126.3550 0.3300 ;
    END
  END bot_S4BEG[14]
  PIN bot_S4BEG[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.49005 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.753 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.6224 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 3.0345 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 12.282 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 61.292 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 125.2650 0.0000 125.4350 0.3300 ;
    END
  END bot_S4BEG[13]
  PIN bot_S4BEG[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.10285 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.121 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.4596 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 7.2205 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 6.5796 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 32.662 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 123.8850 0.0000 124.0550 0.3300 ;
    END
  END bot_S4BEG[12]
  PIN bot_S4BEG[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.16065 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.189 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.558 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 2.7125 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.1751 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.6475 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.09 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 6.28 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 102.218 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 545.632 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 122.5050 0.0000 122.6750 0.3300 ;
    END
  END bot_S4BEG[11]
  PIN bot_S4BEG[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.79645 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.937 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 2.6832 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 13.3385 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.2795 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.2265 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.09 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 6.28 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 97.0938 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 518.304 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 121.1250 0.0000 121.2950 0.3300 ;
    END
  END bot_S4BEG[10]
  PIN bot_S4BEG[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.75905 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.893 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 8.5576 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 42.7105 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.7769 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.7135 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.262 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.864 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 91.4688 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 488.304 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 119.7450 0.0000 119.9150 0.3300 ;
    END
  END bot_S4BEG[9]
  PIN bot_S4BEG[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.27625 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.325 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNADIFFAREA 1.782 LAYER met1  ;
    ANTENNAPARTIALMETALAREA 13.291 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 66.381 LAYER met1  ;
    PORT
      LAYER li1 ;
        RECT 118.3650 0.0000 118.5350 0.3300 ;
    END
  END bot_S4BEG[8]
  PIN bot_S4BEG[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.35745 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.597 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 17.5348 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 87.5595 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.3596 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.68 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 116.9850 0.0000 117.1550 0.3300 ;
    END
  END bot_S4BEG[7]
  PIN bot_S4BEG[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.50745 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.597 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 11.9876 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 59.8605 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.9197 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.4275 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 7.618 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 41.096 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 120.056 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 640.768 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 115.6050 0.0000 115.7750 0.3300 ;
    END
  END bot_S4BEG[6]
  PIN bot_S4BEG[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.02765 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.209 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.9444 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 4.6445 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.8832 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.298 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 114.2250 0.0000 114.3950 0.3300 ;
    END
  END bot_S4BEG[5]
  PIN bot_S4BEG[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.02765 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.209 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.8156 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 4.0005 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.4059 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.8585 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.1905 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.464 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 104.876 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 559.808 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 112.8450 0.0000 113.0150 0.3300 ;
    END
  END bot_S4BEG[4]
  PIN bot_S4BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.73865 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.869 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.88 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 4.3225 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.4544 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.154 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 111.4650 0.0000 111.6350 0.3300 ;
    END
  END bot_S4BEG[3]
  PIN bot_S4BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.10285 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.121 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.236 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.1025 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.5972 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.868 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 110.0850 0.0000 110.2550 0.3300 ;
    END
  END bot_S4BEG[2]
  PIN bot_S4BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.73865 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.869 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.0832 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.4544 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.154 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 108.7050 0.0000 108.8750 0.3300 ;
    END
  END bot_S4BEG[1]
  PIN bot_S4BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.10285 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.121 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.4292 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 2.0685 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.1049 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.4585 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.573 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 8.856 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 121.664 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 649.344 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 107.3250 0.0000 107.4950 0.3300 ;
    END
  END bot_S4BEG[0]
  PIN bot_SS4BEG[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 3.8396 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 19.1205 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.2281 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.9695 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.745 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 4.44 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 38.0478 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 203.392 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 149.1850 0.0000 149.3550 0.3300 ;
    END
  END bot_SS4BEG[15]
  PIN bot_SS4BEG[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.25885 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.481 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.236 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.1025 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 6.0464 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 30.114 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 148.2650 0.0000 148.4350 0.3300 ;
    END
  END bot_SS4BEG[14]
  PIN bot_SS4BEG[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.10285 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.121 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 5.416 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 27.0025 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.1751 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.6475 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.331 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.232 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 22.3578 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 119.712 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 146.8850 0.0000 147.0550 0.3300 ;
    END
  END bot_SS4BEG[13]
  PIN bot_SS4BEG[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.39185 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.461 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 2.2156 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 11.0005 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.6948 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 13.356 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 145.5050 0.0000 145.6750 0.3300 ;
    END
  END bot_SS4BEG[12]
  PIN bot_SS4BEG[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.54785 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.821 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.1716 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.7805 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.6855 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.2565 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.021 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 5.912 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 108.352 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 578.816 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 144.1250 0.0000 144.2950 0.3300 ;
    END
  END bot_SS4BEG[11]
  PIN bot_SS4BEG[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.50745 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.597 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 3.246 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 16.1525 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 4.3161 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 21.4095 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.366 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 7.752 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 90.1878 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 481.472 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 142.7450 0.0000 142.9150 0.3300 ;
    END
  END bot_SS4BEG[10]
  PIN bot_SS4BEG[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.10285 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.121 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.0832 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.1049 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.4585 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.952 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 5.544 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 110.5 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 590.272 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 141.3650 0.0000 141.5350 0.3300 ;
    END
  END bot_SS4BEG[9]
  PIN bot_SS4BEG[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.10285 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.121 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.4292 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 2.0685 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.1049 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.4585 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.504 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 8.488 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 89.1366 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 476.336 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 139.9850 0.0000 140.1550 0.3300 ;
    END
  END bot_SS4BEG[8]
  PIN bot_SS4BEG[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.56525 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.665 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 6.1916 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 30.8805 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.9155 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.4065 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.952 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 5.544 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 127.552 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 681.216 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 138.6050 0.0000 138.7750 0.3300 ;
    END
  END bot_SS4BEG[7]
  PIN bot_SS4BEG[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.49005 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.753 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.236 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.1025 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.5375 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.5165 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.4 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.6 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 125.554 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 670.56 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 137.2250 0.0000 137.3950 0.3300 ;
    END
  END bot_SS4BEG[6]
  PIN bot_SS4BEG[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.54785 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.821 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.1376 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 5.6105 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.3596 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.68 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 135.8450 0.0000 136.0150 0.3300 ;
    END
  END bot_SS4BEG[5]
  PIN bot_SS4BEG[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.16065 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.189 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 3.8564 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 19.2045 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.1751 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.6475 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.262 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.864 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 125.228 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 668.352 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 134.4650 0.0000 134.6350 0.3300 ;
    END
  END bot_SS4BEG[4]
  PIN bot_SS4BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.39185 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.461 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 2.9884 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 14.8645 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 2.3771 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 11.7145 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.676 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 4.072 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 112.841 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 602.288 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 133.0850 0.0000 133.2550 0.3300 ;
    END
  END bot_SS4BEG[3]
  PIN bot_SS4BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.136 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.16 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.3648 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.7465 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.1903 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.7805 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.09 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 6.28 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 114.805 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 613.232 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 131.7050 0.0000 131.8750 0.3300 ;
    END
  END bot_SS4BEG[2]
  PIN bot_SS4BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.10285 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.121 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.0832 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.1049 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.4585 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.331 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.232 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 124.568 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 664.832 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 130.3250 0.0000 130.4950 0.3300 ;
    END
  END bot_SS4BEG[1]
  PIN bot_SS4BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.16065 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.189 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.6868 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 3.3565 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.5496 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.63 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 128.9450 0.0000 129.1150 0.3300 ;
    END
  END bot_SS4BEG[0]
  PIN bot_N1END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.54785 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.821 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.8156 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 4.0005 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.3744 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 14.3331 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 71.0325 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.3744 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 4.402 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 23.944 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.872 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 26.1366 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 140.336 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 13.9450 0.0000 14.1150 0.3300 ;
    END
  END bot_N1END[3]
  PIN bot_N1END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 5.6736 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 28.2905 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.3744 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 6.0627 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 29.7675 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.3744 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.952 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 5.544 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.872 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 49.5927 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 265.896 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 12.5650 0.0000 12.7350 0.3300 ;
    END
  END bot_N1END[2]
  PIN bot_N1END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.27625 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.325 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 4.498 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 22.3755 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.5011 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.3345 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 12.745 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 68.44 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.872 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 27.1932 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 146.912 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 11.1850 0.0000 11.3550 0.3300 ;
    END
  END bot_N1END[1]
  PIN bot_N1END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.56825 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.845 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 14.1436 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 70.6405 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.1872 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 3.0475 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.9485 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.7488 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 6.8668 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 37.56 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.872 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 39.0576 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 209.248 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 10.2650 0.0000 10.4350 0.3300 ;
    END
  END bot_N1END[0]
  PIN bot_N2MID[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.16065 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.189 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.3648 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.7465 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.1751 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.6475 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.331 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.232 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.8864 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 50.4918 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 269.76 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 24.9850 0.0000 25.1550 0.3300 ;
    END
  END bot_N2MID[7]
  PIN bot_N2MID[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.10285 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.121 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.0832 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.1049 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.4585 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.1905 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.464 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.6992 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 101.192 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 541.568 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 23.6050 0.0000 23.7750 0.3300 ;
    END
  END bot_N2MID[6]
  PIN bot_N2MID[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.50745 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.597 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.2664 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 6.2545 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.5175 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.4165 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.469 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.968 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.6992 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 120.478 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 643.488 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 22.2250 0.0000 22.3950 0.3300 ;
    END
  END bot_N2MID[5]
  PIN bot_N2MID[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.10285 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.121 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.0832 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.1049 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.4585 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.1905 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.464 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.692 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 77.2482 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 413.872 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 20.8450 0.0000 21.0150 0.3300 ;
    END
  END bot_N2MID[4]
  PIN bot_N2MID[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.10285 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.121 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.0832 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.1049 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.4585 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.1905 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.464 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.8792 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 60.8361 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 326.336 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 19.4650 0.0000 19.6350 0.3300 ;
    END
  END bot_N2MID[3]
  PIN bot_N2MID[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.16065 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.189 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.9148 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 9.527 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.1036 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.455 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.5616 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 51.8008 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 277.208 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.5048 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 41.4762 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 223.088 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 18.0850 0.0000 18.2550 0.3300 ;
    END
  END bot_N2MID[2]
  PIN bot_N2MID[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.62305 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.733 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 2.5852 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 12.8485 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.4867 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.2625 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.331 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.232 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.692 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 98.142 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 525.776 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 16.7050 0.0000 16.8750 0.3300 ;
    END
  END bot_N2MID[1]
  PIN bot_N2MID[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.73865 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.869 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.6224 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 3.0345 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 9.2721 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 46.1895 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.883 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 5.176 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.8864 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 112.807 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 606.8 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 15.3250 0.0000 15.4950 0.3300 ;
    END
  END bot_N2MID[0]
  PIN bot_N2END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.54785 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.821 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.0832 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.6607 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.1325 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 31.585 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 168.92 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.1376 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 50.6838 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 270.784 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 35.5650 0.0000 35.7350 0.3300 ;
    END
  END bot_N2END[7]
  PIN bot_N2END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.25885 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.481 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 13.9812 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 69.8285 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.7279 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.4685 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.09 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 6.28 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.9504 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 50.6118 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 270.4 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 34.1850 0.0000 34.3550 0.3300 ;
    END
  END bot_N2END[6]
  PIN bot_N2END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.0782 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.092 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 14.8422 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 74.1335 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.9504 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 18.2764 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 90.566 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 33.2650 0.0000 33.4350 0.3300 ;
    END
  END bot_N2END[5]
  PIN bot_N2END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.70425 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 2.005 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.0832 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.1304 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 8.485 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 41.727 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 31.8850 0.0000 32.0550 0.3300 ;
    END
  END bot_N2END[4]
  PIN bot_N2END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.12625 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.325 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 14.8044 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 73.9445 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.1304 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 16.124 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 79.912 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 30.5050 0.0000 30.6750 0.3300 ;
    END
  END bot_N2END[3]
  PIN bot_N2END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.16065 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.189 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.8292 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 9.0685 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.1872 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 7.5649 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 37.2995 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.9432 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.5328 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 3.312 LAYER met3  ;
    PORT
      LAYER li1 ;
        RECT 29.1250 0.0000 29.2950 0.3300 ;
    END
  END bot_N2END[2]
  PIN bot_N2END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.21845 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.257 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.5072 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 7.4585 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.9432 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 15.4104 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 76.482 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 27.7450 0.0000 27.9150 0.3300 ;
    END
  END bot_N2END[1]
  PIN bot_N2END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.3648 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.7465 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.2379 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.0185 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 19.789 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 106.008 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.3248 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 61.6041 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 329.952 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 26.3650 0.0000 26.5350 0.3300 ;
    END
  END bot_N2END[0]
  PIN bot_N4END[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.62305 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.733 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.236 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.1025 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.9304 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.534 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 3.00822 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 13.7374 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 57.1850 0.0000 57.3550 0.3300 ;
    END
  END bot_N4END[15]
  PIN bot_N4END[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.27625 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.325 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.4292 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 2.0685 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 2.216 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.962 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 3.94559 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 18.3333 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 56.2650 0.0000 56.4350 0.3300 ;
    END
  END bot_N4END[14]
  PIN bot_N4END[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.62305 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.733 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.1208 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 5.5265 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 2.0592 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.178 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 3.73441 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 17.2774 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 54.8850 0.0000 55.0550 0.3300 ;
    END
  END bot_N4END[13]
  PIN bot_N4END[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.16065 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.189 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.7004 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 8.4245 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.7876 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.82 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 3.19481 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 13.5859 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 53.5050 0.0000 53.6750 0.3300 ;
    END
  END bot_N4END[12]
  PIN bot_N4END[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.54785 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.821 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.0832 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 4.12 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 20.482 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 8.54626 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 41.3367 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 52.1250 0.0000 52.2950 0.3300 ;
    END
  END bot_N4END[11]
  PIN bot_N4END[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.68085 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.801 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.2328 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 6.0865 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.5356 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.56 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 4.74983 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 21.6586 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 50.7450 0.0000 50.9150 0.3300 ;
    END
  END bot_N4END[10]
  PIN bot_N4END[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.27625 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.325 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 2.1512 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 10.6785 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.5764 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.646 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 1.3037 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 4.96498 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 49.3650 0.0000 49.5350 0.3300 ;
    END
  END bot_N4END[9]
  PIN bot_N4END[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.10285 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.121 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 8.5408 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 42.6265 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 10.3986 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 51.639 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 14.8792 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 72.6835 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 47.9850 0.0000 48.1550 0.3300 ;
    END
  END bot_N4END[8]
  PIN bot_N4END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.45265 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.709 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 8.5384 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 42.5775 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.2981 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.3195 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 11.44 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 61.48 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.9432 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 29.079 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 157.44 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 46.6050 0.0000 46.7750 0.3300 ;
    END
  END bot_N4END[7]
  PIN bot_N4END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.43225 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.685 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.4596 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 7.2205 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.1335 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.5355 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.883 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 5.176 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.9432 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 73.4388 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 392.144 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 45.2250 0.0000 45.3950 0.3300 ;
    END
  END bot_N4END[6]
  PIN bot_N4END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.14325 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.345 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.9444 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 4.6445 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.3107 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.3825 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.331 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.232 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.9432 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 107.22 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 574.192 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 43.8450 0.0000 44.0150 0.3300 ;
    END
  END bot_N4END[5]
  PIN bot_N4END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.62305 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.733 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.5072 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 7.4585 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.0331 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.9945 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.273 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 7.256 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.9432 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 99.0363 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 529.6 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 42.4650 0.0000 42.6350 0.3300 ;
    END
  END bot_N4END[4]
  PIN bot_N4END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.31665 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.549 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.202 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 5.9325 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 3.1643 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 15.4875 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.4 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.6 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.9432 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 45.8715 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 245.584 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 41.0850 0.0000 41.2550 0.3300 ;
    END
  END bot_N4END[3]
  PIN bot_N4END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.16065 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.189 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.1716 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.7805 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.9432 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 11.7056 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 57.722 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 39.7050 0.0000 39.8750 0.3300 ;
    END
  END bot_N4END[2]
  PIN bot_N4END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.54785 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.821 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.0832 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.9603 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.6305 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.814 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 4.808 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.9432 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 14.0988 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 75.664 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 38.3250 0.0000 38.4950 0.3300 ;
    END
  END bot_N4END[1]
  PIN bot_N4END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.14325 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.345 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.4292 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 2.0685 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.1908 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.9507 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.4745 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.1908 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 2.746 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 15.112 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.9432 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 14.0748 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 75.536 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 36.9450 0.0000 37.1150 0.3300 ;
    END
  END bot_N4END[0]
  PIN bot_NN4END[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.62305 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.733 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.3004 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.4245 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.9304 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.534 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 3.90788 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 18.1448 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 79.2650 0.0000 79.4350 0.3300 ;
    END
  END bot_NN4END[15]
  PIN bot_NN4END[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.21845 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.257 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.1852 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 5.8485 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 2.2636 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 11.2 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 4.0097 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 18.6539 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 77.8850 0.0000 78.0550 0.3300 ;
    END
  END bot_NN4END[14]
  PIN bot_NN4END[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.16065 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.189 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.558 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 2.7125 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 15.4729 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 76.4855 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 12.1608 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 70.032 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met3  ;
    ANTENNAMAXAREACAR 32.6924 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 174.106 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.123098 LAYER via3  ;
    PORT
      LAYER li1 ;
        RECT 76.5050 0.0000 76.6750 0.3300 ;
    END
  END bot_NN4END[13]
  PIN bot_NN4END[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.37445 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.617 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.846 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 9.1525 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.2095 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.8765 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 13.3512 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 75.44 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met3  ;
    ANTENNAMAXAREACAR 33.3924 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 175.673 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.123098 LAYER via3  ;
    PORT
      LAYER li1 ;
        RECT 75.1250 0.0000 75.2950 0.3300 ;
    END
  END bot_NN4END[12]
  PIN bot_NN4END[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.10285 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.121 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.524 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 7.5425 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.8352 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.058 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 3.25892 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 13.9064 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 73.7450 0.0000 73.9150 0.3300 ;
    END
  END bot_NN4END[11]
  PIN bot_NN4END[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.62305 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.733 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 16.5996 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 82.887 LAYER met1  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met1  ;
    ANTENNAMAXAREACAR 22.9904 LAYER met1  ;
    ANTENNAMAXSIDEAREACAR 112.38 LAYER met1  ;
    ANTENNAMAXCUTCAR 0.0389226 LAYER via  ;
    PORT
      LAYER li1 ;
        RECT 72.3650 0.0000 72.5350 0.3300 ;
    END
  END bot_NN4END[10]
  PIN bot_NN4END[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.27625 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.325 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.992 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 4.8825 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 2.216 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.962 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 3.94559 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 18.3333 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 70.9850 0.0000 71.1550 0.3300 ;
    END
  END bot_NN4END[9]
  PIN bot_NN4END[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.44965 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.529 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.2664 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 6.2545 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 14.0201 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 69.4575 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 11.2812 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 64.4 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met3  ;
    ANTENNAMAXAREACAR 18.6436 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 101.345 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.123098 LAYER via3  ;
    PORT
      LAYER li1 ;
        RECT 69.6050 0.0000 69.7750 0.3300 ;
    END
  END bot_NN4END[8]
  PIN bot_NN4END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.68085 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.801 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 2.6188 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 13.0165 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.0331 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.9945 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.1249 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.136 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.5616 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 109.117 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 582.896 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 68.2250 0.0000 68.3950 0.3300 ;
    END
  END bot_NN4END[7]
  PIN bot_NN4END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.16065 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.189 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.88 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 4.3225 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 5.2753 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 26.1205 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.469 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.968 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.5616 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 70.7418 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 377.76 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 66.8450 0.0000 67.0150 0.3300 ;
    END
  END bot_NN4END[6]
  PIN bot_NN4END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.21845 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.257 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.558 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 2.7125 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.0723 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.1905 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.1905 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.464 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.5616 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 85.9146 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 459.152 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 65.4650 0.0000 65.6350 0.3300 ;
    END
  END bot_NN4END[5]
  PIN bot_NN4END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.33405 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.393 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.6528 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 8.1865 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 3.8597 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 19.1275 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.159 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 6.648 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.3744 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 59.0136 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 315.68 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 64.0850 0.0000 64.2550 0.3300 ;
    END
  END bot_NN4END[4]
  PIN bot_NN4END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.56525 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.665 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 2.6664 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 13.2545 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.0009 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.8335 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.952 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 5.544 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.5616 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 34.4742 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 185.744 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 62.7050 0.0000 62.8750 0.3300 ;
    END
  END bot_NN4END[3]
  PIN bot_NN4END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.54785 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.821 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.0832 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.1872 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 6.6759 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 32.8545 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.1872 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 5.851 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 31.672 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.5616 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 3.0948 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 16.976 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 61.3250 0.0000 61.4950 0.3300 ;
    END
  END bot_NN4END[2]
  PIN bot_NN4END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.68085 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.801 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.0832 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.1872 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 11.4588 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 56.854 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via2  ;
    ANTENNADIFFAREA 0.5616 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 14.8656 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 80.224 LAYER met3  ;
    PORT
      LAYER li1 ;
        RECT 59.9450 0.0000 60.1150 0.3300 ;
    END
  END bot_NN4END[1]
  PIN bot_NN4END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.16065 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.189 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.1376 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 5.6105 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.2487 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.0725 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.435 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 8.12 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.3744 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 18.4908 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 99.088 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 58.5650 0.0000 58.7350 0.3300 ;
    END
  END bot_NN4END[0]
  PIN UserCLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.0114 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 16.056 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 4.608 LAYER met4  ;
    ANTENNAMAXAREACAR 7.70864 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 40.2318 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.0473307 LAYER via4  ;
    PORT
      LAYER met4 ;
        RECT 89.5500 0.0000 89.8500 0.8000 ;
    END
  END UserCLK
  PIN top_FrameData[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 9.5215 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 46.6305 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.113 LAYER met2  ;
    ANTENNAMAXAREACAR 42.6454 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 208.223 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.500719 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.538 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 3.336 LAYER met3  ;
    ANTENNAGATEAREA 1.113 LAYER met3  ;
    ANTENNAMAXAREACAR 43.1287 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 211.221 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.536658 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 19.0497 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 102.064 LAYER met4  ;
    ANTENNAGATEAREA 2.8095 LAYER met4  ;
    ANTENNAMAXAREACAR 59.3483 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 294.966 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.548637 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 434.2800 0.4850 434.4200 ;
    END
  END top_FrameData[31]
  PIN top_FrameData[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 30.464 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 150.311 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.067 LAYER met2  ;
    ANTENNAMAXAREACAR 67.2049 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 330.927 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.625641 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 5.3628 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 29.072 LAYER met3  ;
    ANTENNAGATEAREA 2.8095 LAYER met3  ;
    ANTENNAMAXAREACAR 69.1137 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 341.275 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.625641 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 432.5800 0.4850 432.7200 ;
    END
  END top_FrameData[30]
  PIN top_FrameData[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1561 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.6195 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 23.0724 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 123.984 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.8095 LAYER met3  ;
    ANTENNAMAXAREACAR 47.2458 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 234.215 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.632495 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 430.8800 0.4850 431.0200 ;
    END
  END top_FrameData[29]
  PIN top_FrameData[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 11.1845 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 54.7225 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.6965 LAYER met2  ;
    ANTENNAMAXAREACAR 16.1722 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 78.6272 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.346848 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 12.5266 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 68.216 LAYER met3  ;
    ANTENNAGATEAREA 2.1735 LAYER met3  ;
    ANTENNAMAXAREACAR 40.0463 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 196.524 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.986328 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 27.0537 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 144.752 LAYER met4  ;
    ANTENNAGATEAREA 2.8095 LAYER met4  ;
    ANTENNAMAXAREACAR 49.6757 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 248.046 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.986328 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 429.1800 0.4850 429.3200 ;
    END
  END top_FrameData[28]
  PIN top_FrameData[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2555 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.1165 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 22.6378 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 121.672 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.3325 LAYER met3  ;
    ANTENNAMAXAREACAR 46.8364 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 232.896 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.516227 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 1.3998 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 7.936 LAYER met4  ;
    ANTENNAGATEAREA 2.8095 LAYER met4  ;
    ANTENNAMAXAREACAR 47.3346 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 235.721 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.516227 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 427.4800 0.4850 427.6200 ;
    END
  END top_FrameData[27]
  PIN top_FrameData[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.6056 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.749 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 7.77966 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 37.1414 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.153401 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.331 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.232 LAYER met3  ;
    ANTENNAGATEAREA 0.7425 LAYER met3  ;
    ANTENNAMAXAREACAR 8.22545 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 40.1475 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.207273 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 11.3298 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 60.896 LAYER met4  ;
    ANTENNAGATEAREA 2.8095 LAYER met4  ;
    ANTENNAMAXAREACAR 41.479 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 208.16 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.609918 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 425.7800 0.4850 425.9200 ;
    END
  END top_FrameData[26]
  PIN top_FrameData[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 15.9911 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 78.9355 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.0605 LAYER met2  ;
    ANTENNAMAXAREACAR 18.3011 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 88.169 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.398707 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 5.144 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 28.368 LAYER met3  ;
    ANTENNAGATEAREA 1.0605 LAYER met3  ;
    ANTENNAMAXAREACAR 23.1517 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 114.919 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.474143 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 19.6131 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 106.48 LAYER met4  ;
    ANTENNAGATEAREA 2.8095 LAYER met4  ;
    ANTENNAMAXAREACAR 39.2867 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 198.854 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.07799 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 424.0800 0.4850 424.2200 ;
    END
  END top_FrameData[25]
  PIN top_FrameData[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 17.512 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 86.422 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.0605 LAYER met2  ;
    ANTENNAMAXAREACAR 23.313 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 112.045 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.398707 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.4848 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 8.856 LAYER met3  ;
    ANTENNAGATEAREA 1.2195 LAYER met3  ;
    ANTENNAMAXAREACAR 24.5305 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 119.307 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.607643 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 8.6796 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 47.232 LAYER met4  ;
    ANTENNAGATEAREA 2.8095 LAYER met4  ;
    ANTENNAMAXAREACAR 39.5632 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 199.226 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.779245 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 422.0400 0.4850 422.1800 ;
    END
  END top_FrameData[24]
  PIN top_FrameData[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 18.8565 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 93.5515 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.3785 LAYER met2  ;
    ANTENNAMAXAREACAR 26.3998 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 127.343 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.493797 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 13.1808 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 70.768 LAYER met3  ;
    ANTENNAGATEAREA 2.8095 LAYER met3  ;
    ANTENNAMAXAREACAR 49.3615 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 243.947 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.634242 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 420.3400 0.4850 420.4800 ;
    END
  END top_FrameData[23]
  PIN top_FrameData[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 19.6636 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 97.426 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.3785 LAYER met2  ;
    ANTENNAMAXAREACAR 27.1488 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 131.65 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.522814 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 31.4296 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 169.032 LAYER met3  ;
    ANTENNAGATEAREA 2.1735 LAYER met3  ;
    ANTENNAMAXAREACAR 88.595 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 442.166 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.986328 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 1.5828 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 8.912 LAYER met4  ;
    ANTENNAGATEAREA 2.8095 LAYER met4  ;
    ANTENNAMAXAREACAR 89.1583 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 445.338 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.986328 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 418.6400 0.4850 418.7800 ;
    END
  END top_FrameData[22]
  PIN top_FrameData[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 18.9117 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 93.6845 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.636 LAYER met2  ;
    ANTENNAMAXAREACAR 42.1002 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 205.68 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.527673 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 20.8036 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 112.36 LAYER met3  ;
    ANTENNAGATEAREA 1.8555 LAYER met3  ;
    ANTENNAMAXAREACAR 53.312 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 266.235 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.73791 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 20.8296 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 112.032 LAYER met4  ;
    ANTENNAGATEAREA 2.8095 LAYER met4  ;
    ANTENNAMAXAREACAR 60.726 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 306.111 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.857862 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 416.9400 0.4850 417.0800 ;
    END
  END top_FrameData[21]
  PIN top_FrameData[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 17.7632 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 88.095 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.3785 LAYER met2  ;
    ANTENNAMAXAREACAR 21.7677 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 104.189 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.493797 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 7.4638 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 40.744 LAYER met3  ;
    ANTENNAGATEAREA 1.8555 LAYER met3  ;
    ANTENNAMAXAREACAR 42.9638 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 210.357 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.795562 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 2.0676 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 11.968 LAYER met4  ;
    ANTENNAGATEAREA 2.8095 LAYER met4  ;
    ANTENNAMAXAREACAR 51.2107 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 252.536 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.795562 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 415.2400 0.4850 415.3800 ;
    END
  END top_FrameData[20]
  PIN top_FrameData[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2051 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.8645 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 9.067 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 48.824 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 3.4032 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 20.032 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.8095 LAYER met4  ;
    ANTENNAMAXAREACAR 38.4332 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 191.348 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.677394 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 413.5400 0.4850 413.6800 ;
    END
  END top_FrameData[19]
  PIN top_FrameData[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1757 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.7175 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 49.605 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 265.472 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.8095 LAYER met3  ;
    ANTENNAMAXAREACAR 53.0447 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 265.907 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.706918 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 411.5000 0.4850 411.6400 ;
    END
  END top_FrameData[18]
  PIN top_FrameData[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.2187 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.9325 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 25.2483 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 136.064 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.8095 LAYER met3  ;
    ANTENNAMAXAREACAR 54.0778 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 268.341 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.590566 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 409.8000 0.4850 409.9400 ;
    END
  END top_FrameData[17]
  PIN top_FrameData[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1267 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.4725 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 29.9512 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 160.672 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.4915 LAYER met3  ;
    ANTENNAMAXAREACAR 41.8206 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 208.406 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.526575 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 10.9158 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 58.688 LAYER met4  ;
    ANTENNAGATEAREA 2.8095 LAYER met4  ;
    ANTENNAMAXAREACAR 45.7059 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 229.295 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.716352 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 408.1000 0.4850 408.2400 ;
    END
  END top_FrameData[16]
  PIN top_FrameData[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1449 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.5635 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 13.645 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 73.24 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 42.0516 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 227.088 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.8095 LAYER met4  ;
    ANTENNAMAXAREACAR 74.5375 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 375.021 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.07799 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 406.4000 0.4850 406.5400 ;
    END
  END top_FrameData[15]
  PIN top_FrameData[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2297 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.7945 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 29.8854 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 160.8 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.8095 LAYER met3  ;
    ANTENNAMAXAREACAR 46.8217 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 233.246 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.632495 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 404.7000 0.4850 404.8400 ;
    END
  END top_FrameData[14]
  PIN top_FrameData[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.0215 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.7105 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 28.6626 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 153.808 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.8095 LAYER met3  ;
    ANTENNAMAXAREACAR 71.6446 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 356.79 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.635306 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 403.0000 0.4850 403.1400 ;
    END
  END top_FrameData[13]
  PIN top_FrameData[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.3631 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.5365 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 9.988 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 53.736 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 36.8085 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 197.248 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.8095 LAYER met4  ;
    ANTENNAMAXAREACAR 83.3345 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 435.421 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.2195 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 400.9600 0.4850 401.1000 ;
    END
  END top_FrameData[12]
  PIN top_FrameData[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 5.0405 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 24.9235 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 60.187 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 323.336 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.4915 LAYER met3  ;
    ANTENNAMAXAREACAR 97.5532 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 491.222 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.983979 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.6678 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 4.032 LAYER met4  ;
    ANTENNAGATEAREA 2.8095 LAYER met4  ;
    ANTENNAMAXAREACAR 97.7909 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 492.657 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.983979 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 399.2600 0.4850 399.4000 ;
    END
  END top_FrameData[11]
  PIN top_FrameData[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2037 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.8575 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 24.13 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 129.16 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 15.1566 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 81.776 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.8095 LAYER met4  ;
    ANTENNAMAXAREACAR 48.6699 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 247.083 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.752291 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 397.5600 0.4850 397.7000 ;
    END
  END top_FrameData[10]
  PIN top_FrameData[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.858 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.011 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 25.12 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 134.44 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 47.3409 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 254.832 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.6505 LAYER met4  ;
    ANTENNAMAXAREACAR 71.2749 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 365.687 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.07799 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 395.8600 0.4850 396.0000 ;
    END
  END top_FrameData[9]
  PIN top_FrameData[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1699 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.6335 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 44.7272 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 239.944 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.3785 LAYER met3  ;
    ANTENNAMAXAREACAR 51.497 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 264.225 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.690529 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 47.9586 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 259.072 LAYER met4  ;
    ANTENNAGATEAREA 2.6505 LAYER met4  ;
    ANTENNAMAXAREACAR 69.5912 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 361.97 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.07799 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 394.1600 0.4850 394.3000 ;
    END
  END top_FrameData[8]
  PIN top_FrameData[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2429 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.0535 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.469 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.968 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 41.4315 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 221.904 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.6505 LAYER met4  ;
    ANTENNAMAXAREACAR 46.7344 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 234.707 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.826415 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 392.4600 0.4850 392.6000 ;
    END
  END top_FrameData[7]
  PIN top_FrameData[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2135 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.9065 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 34.186 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 182.792 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 77.5098 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 414.792 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.6505 LAYER met4  ;
    ANTENNAMAXAREACAR 58.1264 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 301.053 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.07574 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 390.4200 0.4850 390.5600 ;
    END
  END top_FrameData[6]
  PIN top_FrameData[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2317 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.9975 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.262 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.864 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 22.1976 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 119.328 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.6505 LAYER met4  ;
    ANTENNAMAXAREACAR 41.3361 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 207.577 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.530186 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 388.7200 0.4850 388.8600 ;
    END
  END top_FrameData[5]
  PIN top_FrameData[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.1514 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 15.596 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 2.125 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 11.8 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 36.3207 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 196.528 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.6505 LAYER met4  ;
    ANTENNAMAXAREACAR 41.7442 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 216.402 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.842138 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 387.0200 0.4850 387.1600 ;
    END
  END top_FrameData[4]
  PIN top_FrameData[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 10.6469 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 52.6015 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.477 LAYER met2  ;
    ANTENNAMAXAREACAR 46.1627 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 225.732 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.548637 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 10.9804 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 59.024 LAYER met3  ;
    ANTENNAGATEAREA 0.954 LAYER met3  ;
    ANTENNAMAXAREACAR 57.6725 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 287.602 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.590566 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 20.5746 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 110.672 LAYER met4  ;
    ANTENNAGATEAREA 2.6505 LAYER met4  ;
    ANTENNAMAXAREACAR 65.4351 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 329.357 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.826415 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 385.3200 0.4850 385.4600 ;
    END
  END top_FrameData[3]
  PIN top_FrameData[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.5502 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.59 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 10.129 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 54.488 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 40.4892 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 217.824 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.6505 LAYER met4  ;
    ANTENNAMAXAREACAR 72.7333 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 383.481 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.07799 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 383.6200 0.4850 383.7600 ;
    END
  END top_FrameData[2]
  PIN top_FrameData[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1337 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.5075 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 18.7178 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 101.232 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 19.881 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 108.384 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.6505 LAYER met4  ;
    ANTENNAMAXAREACAR 55.5544 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 277.129 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.826415 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 381.9200 0.4850 382.0600 ;
    END
  END top_FrameData[1]
  PIN top_FrameData[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7033 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.2375 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 8.563 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 46.136 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 37.6419 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 203.104 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.6505 LAYER met4  ;
    ANTENNAMAXAREACAR 50.8841 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 257.831 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.27153 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 380.2200 0.4850 380.3600 ;
    END
  END top_FrameData[0]
  PIN top_FrameData_O[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.9342 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.445 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 209.7350 434.2800 210.2200 434.4200 ;
    END
  END top_FrameData_O[31]
  PIN top_FrameData_O[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.6635 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.2095 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 209.7350 432.5800 210.2200 432.7200 ;
    END
  END top_FrameData_O[30]
  PIN top_FrameData_O[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.7151 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.3495 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 209.7350 430.8800 210.2200 431.0200 ;
    END
  END top_FrameData_O[29]
  PIN top_FrameData_O[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2352 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.015 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 51.0798 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 272.896 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 209.7350 429.1800 210.2200 429.3200 ;
    END
  END top_FrameData_O[28]
  PIN top_FrameData_O[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.4282 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.862 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 22.8888 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 122.544 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 209.7350 427.4800 210.2200 427.6200 ;
    END
  END top_FrameData_O[27]
  PIN top_FrameData_O[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2107 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.8925 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 53.0178 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 283.232 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 209.7350 425.7800 210.2200 425.9200 ;
    END
  END top_FrameData_O[26]
  PIN top_FrameData_O[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.672 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.199 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 54.355 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 290.36 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 0.6678 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 4.032 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 209.7350 424.0800 210.2200 424.2200 ;
    END
  END top_FrameData_O[25]
  PIN top_FrameData_O[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.8411 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 13.9265 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 42.391 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 226.552 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 11.9106 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 64.464 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 209.7350 422.0400 210.2200 422.1800 ;
    END
  END top_FrameData_O[24]
  PIN top_FrameData_O[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.3626 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.652 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 57.0588 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 304.784 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 209.7350 420.3400 210.2200 420.4800 ;
    END
  END top_FrameData_O[23]
  PIN top_FrameData_O[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1561 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.6195 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 57.1023 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 305.016 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 209.7350 418.6400 210.2200 418.7800 ;
    END
  END top_FrameData_O[22]
  PIN top_FrameData_O[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2408 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.043 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 38.506 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 205.832 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 0.6678 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 4.032 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 209.7350 416.9400 210.2200 417.0800 ;
    END
  END top_FrameData_O[21]
  PIN top_FrameData_O[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1869 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.7735 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 57.2418 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 305.76 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 209.7350 415.2400 210.2200 415.3800 ;
    END
  END top_FrameData_O[20]
  PIN top_FrameData_O[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.4338 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.89 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 10.7448 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 57.776 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 209.7350 413.5400 210.2200 413.6800 ;
    END
  END top_FrameData_O[19]
  PIN top_FrameData_O[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1757 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.7175 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 11.8008 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 63.408 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 209.7350 411.5000 210.2200 411.6400 ;
    END
  END top_FrameData_O[18]
  PIN top_FrameData_O[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1939 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.8085 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 13.6848 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 73.456 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 209.7350 409.8000 210.2200 409.9400 ;
    END
  END top_FrameData_O[17]
  PIN top_FrameData_O[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1267 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.4725 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 6.9708 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 37.648 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 209.7350 408.1000 210.2200 408.2400 ;
    END
  END top_FrameData_O[16]
  PIN top_FrameData_O[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.1609 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.6965 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 209.7350 406.4000 210.2200 406.5400 ;
    END
  END top_FrameData_O[15]
  PIN top_FrameData_O[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.1028 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 209.7350 404.7000 210.2200 404.8400 ;
    END
  END top_FrameData_O[14]
  PIN top_FrameData_O[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.0468 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.126 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 209.7350 403.0000 210.2200 403.1400 ;
    END
  END top_FrameData_O[13]
  PIN top_FrameData_O[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.1462 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.623 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 209.7350 400.9600 210.2200 401.1000 ;
    END
  END top_FrameData_O[12]
  PIN top_FrameData_O[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.5203 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.4935 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 209.7350 399.2600 210.2200 399.4000 ;
    END
  END top_FrameData_O[11]
  PIN top_FrameData_O[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.0468 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.126 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 209.7350 397.5600 210.2200 397.7000 ;
    END
  END top_FrameData_O[10]
  PIN top_FrameData_O[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.1938 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.861 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 209.7350 395.8600 210.2200 396.0000 ;
    END
  END top_FrameData_O[9]
  PIN top_FrameData_O[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.2456 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.12 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 209.7350 394.1600 210.2200 394.3000 ;
    END
  END top_FrameData_O[8]
  PIN top_FrameData_O[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.1938 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.861 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 209.7350 392.4600 210.2200 392.6000 ;
    END
  END top_FrameData_O[7]
  PIN top_FrameData_O[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.4107 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 11.9455 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 209.7350 390.4200 210.2200 390.5600 ;
    END
  END top_FrameData_O[6]
  PIN top_FrameData_O[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.1028 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 209.7350 388.7200 210.2200 388.8600 ;
    END
  END top_FrameData_O[5]
  PIN top_FrameData_O[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.2456 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.12 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 209.7350 387.0200 210.2200 387.1600 ;
    END
  END top_FrameData_O[4]
  PIN top_FrameData_O[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.1938 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.861 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 209.7350 385.3200 210.2200 385.4600 ;
    END
  END top_FrameData_O[3]
  PIN top_FrameData_O[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.4395 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.0895 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 209.7350 383.6200 210.2200 383.7600 ;
    END
  END top_FrameData_O[2]
  PIN top_FrameData_O[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.2456 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.12 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 209.7350 381.9200 210.2200 382.0600 ;
    END
  END top_FrameData_O[1]
  PIN top_FrameData_O[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.3668 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.608 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 209.7350 380.2200 210.2200 380.3600 ;
    END
  END top_FrameData_O[0]
  PIN bot_FrameData[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1379 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.5285 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 50.8783 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 273.224 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.0145 LAYER met3  ;
    ANTENNAMAXAREACAR 54.8538 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 279.071 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.987781 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 8.7198 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 46.976 LAYER met4  ;
    ANTENNAGATEAREA 2.8095 LAYER met4  ;
    ANTENNAMAXAREACAR 57.9575 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 295.792 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.987781 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 209.5400 0.4850 209.6800 ;
    END
  END bot_FrameData[31]
  PIN bot_FrameData[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.6559 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.1185 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 57.9904 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 310.68 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.3325 LAYER met3  ;
    ANTENNAMAXAREACAR 58.9102 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 298.243 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.649644 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 1.0338 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 5.984 LAYER met4  ;
    ANTENNAGATEAREA 2.8095 LAYER met4  ;
    ANTENNAMAXAREACAR 59.2782 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 300.373 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.6587 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 207.8400 0.4850 207.9800 ;
    END
  END bot_FrameData[30]
  PIN bot_FrameData[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.3981 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.7115 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 7.231 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 39.032 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 33.3402 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 179.216 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.8095 LAYER met4  ;
    ANTENNAMAXAREACAR 88.4758 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 456.349 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.32956 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 206.1400 0.4850 206.2800 ;
    END
  END bot_FrameData[29]
  PIN bot_FrameData[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.6303 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.9905 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 33.7097 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 181.192 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.113 LAYER met3  ;
    ANTENNAMAXAREACAR 91.3138 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 462.054 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.785984 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 44.5797 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 240.576 LAYER met4  ;
    ANTENNAGATEAREA 2.8095 LAYER met4  ;
    ANTENNAMAXAREACAR 107.181 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 547.683 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.07799 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 204.4400 0.4850 204.5800 ;
    END
  END bot_FrameData[28]
  PIN bot_FrameData[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.6373 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 22.9075 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 49.9252 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 268.136 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.8555 LAYER met3  ;
    ANTENNAMAXAREACAR 50.4425 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 257.125 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.863696 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 15.5388 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 83.344 LAYER met4  ;
    ANTENNAGATEAREA 2.8095 LAYER met4  ;
    ANTENNAMAXAREACAR 55.9733 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 286.79 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.863696 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 202.7400 0.4850 202.8800 ;
    END
  END bot_FrameData[27]
  PIN bot_FrameData[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1323 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.5005 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 22.9618 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 123.4 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.318 LAYER met3  ;
    ANTENNAMAXAREACAR 116.17 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 601.924 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.842138 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 27.0777 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 144.88 LAYER met4  ;
    ANTENNAGATEAREA 2.8095 LAYER met4  ;
    ANTENNAMAXAREACAR 125.808 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 653.492 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.842138 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 201.0400 0.4850 201.1800 ;
    END
  END bot_FrameData[26]
  PIN bot_FrameData[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7161 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.4195 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 47.3242 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 254.264 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.4915 LAYER met3  ;
    ANTENNAMAXAREACAR 42.5792 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 214.405 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.983979 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 26.9187 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 144.032 LAYER met4  ;
    ANTENNAGATEAREA 2.8095 LAYER met4  ;
    ANTENNAMAXAREACAR 52.1605 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 269.684 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.983979 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 199.0000 0.4850 199.1400 ;
    END
  END bot_FrameData[25]
  PIN bot_FrameData[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2289 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.9835 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 19.0558 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 102.568 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.318 LAYER met3  ;
    ANTENNAMAXAREACAR 87.5987 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 455.343 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.842138 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 16.5597 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 88.784 LAYER met4  ;
    ANTENNAGATEAREA 2.8095 LAYER met4  ;
    ANTENNAMAXAREACAR 93.4929 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 486.944 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.09371 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 197.3000 0.4850 197.4400 ;
    END
  END bot_FrameData[24]
  PIN bot_FrameData[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1253 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.4655 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 20.038 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 107.336 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 91.9029 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 491.056 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.8095 LAYER met4  ;
    ANTENNAMAXAREACAR 100.294 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 521.441 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.826415 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 195.6000 0.4850 195.7400 ;
    END
  END bot_FrameData[23]
  PIN bot_FrameData[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.4732 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.205 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 39.0172 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 209.024 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.8555 LAYER met3  ;
    ANTENNAMAXAREACAR 55.5795 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 281.418 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.515354 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 12.5868 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 67.6 LAYER met4  ;
    ANTENNAGATEAREA 2.8095 LAYER met4  ;
    ANTENNAMAXAREACAR 60.0596 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 305.479 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.548637 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 193.9000 0.4850 194.0400 ;
    END
  END bot_FrameData[22]
  PIN bot_FrameData[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1743 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.7105 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 31.813 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 170.136 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 25.6746 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 137.872 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.8095 LAYER met4  ;
    ANTENNAMAXAREACAR 71.1435 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 368.34 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.700601 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 192.2000 0.4850 192.3400 ;
    END
  END bot_FrameData[21]
  PIN bot_FrameData[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1883 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.7805 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 11.989 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 64.408 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 67.1223 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 359.392 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.8095 LAYER met4  ;
    ANTENNAMAXAREACAR 93.0252 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 492.188 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.07799 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 190.1600 0.4850 190.3000 ;
    END
  END bot_FrameData[20]
  PIN bot_FrameData[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2065 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.8715 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 45.1015 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 241.944 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.5375 LAYER met3  ;
    ANTENNAMAXAREACAR 56.3233 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 287.433 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.993941 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 4.9956 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 27.584 LAYER met4  ;
    ANTENNAGATEAREA 2.8095 LAYER met4  ;
    ANTENNAMAXAREACAR 58.1014 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 297.251 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.993941 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 188.4600 0.4850 188.6000 ;
    END
  END bot_FrameData[19]
  PIN bot_FrameData[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2247 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.9625 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 26.335 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 140.92 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 1.3998 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 7.936 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.8095 LAYER met4  ;
    ANTENNAMAXAREACAR 36.592 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 178.756 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.493255 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 186.7600 0.4850 186.9000 ;
    END
  END bot_FrameData[18]
  PIN bot_FrameData[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.987 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.774 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 48.109 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 257.504 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.5375 LAYER met3  ;
    ANTENNAMAXAREACAR 51.5485 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 263.846 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.600859 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 17.0172 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 92.64 LAYER met4  ;
    ANTENNAGATEAREA 2.8095 LAYER met4  ;
    ANTENNAMAXAREACAR 58.6706 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 299.694 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.826415 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 185.0600 0.4850 185.2000 ;
    END
  END bot_FrameData[17]
  PIN bot_FrameData[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.6275 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.9765 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 59.2485 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 318.8 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.8095 LAYER met3  ;
    ANTENNAMAXAREACAR 54.6097 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 274.945 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.842138 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 183.3600 0.4850 183.5000 ;
    END
  END bot_FrameData[16]
  PIN bot_FrameData[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1603 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.6405 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.676 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 4.072 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 70.6506 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 380.096 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.8095 LAYER met4  ;
    ANTENNAMAXAREACAR 86.4131 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 449.802 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.47107 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 181.3200 0.4850 181.4600 ;
    END
  END bot_FrameData[15]
  PIN bot_FrameData[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2499 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.0885 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 2.722 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 14.984 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 54.0138 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 290.896 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.8095 LAYER met4  ;
    ANTENNAMAXAREACAR 78.7458 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 402.884 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.32956 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 179.6200 0.4850 179.7600 ;
    END
  END bot_FrameData[14]
  PIN bot_FrameData[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1827 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.7525 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 18.454 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 98.888 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 20.4417 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 109.488 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.8095 LAYER met4  ;
    ANTENNAMAXAREACAR 68.9132 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 353.869 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.985074 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 177.9200 0.4850 178.0600 ;
    END
  END bot_FrameData[13]
  PIN bot_FrameData[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.4541 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.9915 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 4.44094 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 20.398 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.153401 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 22.5264 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 121.552 LAYER met3  ;
    ANTENNAGATEAREA 2.8095 LAYER met3  ;
    ANTENNAMAXAREACAR 73.9998 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 368.134 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.690147 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 176.2200 0.4850 176.3600 ;
    END
  END bot_FrameData[12]
  PIN bot_FrameData[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.1585 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.6315 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 12.796 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 68.712 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 8.7438 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 47.104 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.8095 LAYER met4  ;
    ANTENNAMAXAREACAR 49.5109 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 244.629 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.776274 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 174.5200 0.4850 174.6600 ;
    END
  END bot_FrameData[11]
  PIN bot_FrameData[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.5717 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.5795 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 38.7381 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 207.992 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.1735 LAYER met3  ;
    ANTENNAMAXAREACAR 47.9762 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 241.562 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.567041 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 6.9138 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 37.344 LAYER met4  ;
    ANTENNAGATEAREA 2.8095 LAYER met4  ;
    ANTENNAMAXAREACAR 50.4371 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 254.854 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.590566 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 172.4800 0.4850 172.6200 ;
    END
  END bot_FrameData[10]
  PIN bot_FrameData[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.1953 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 15.6975 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 33.3903 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 179.488 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.8095 LAYER met3  ;
    ANTENNAMAXAREACAR 49.4294 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 247.229 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.574843 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 170.7800 0.4850 170.9200 ;
    END
  END bot_FrameData[9]
  PIN bot_FrameData[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.6951 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.3145 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 48.1351 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 257.648 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.6505 LAYER met3  ;
    ANTENNAMAXAREACAR 40.8133 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 206.116 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.51581 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 14.5758 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 78.208 LAYER met4  ;
    ANTENNAGATEAREA 2.8095 LAYER met4  ;
    ANTENNAMAXAREACAR 46.0014 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 233.953 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.826415 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 169.0800 0.4850 169.2200 ;
    END
  END bot_FrameData[8]
  PIN bot_FrameData[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1589 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.6335 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 10.564 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 56.808 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 22.968 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 124.848 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.8095 LAYER met4  ;
    ANTENNAMAXAREACAR 77.8971 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 407.266 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.826415 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 167.3800 0.4850 167.5200 ;
    END
  END bot_FrameData[7]
  PIN bot_FrameData[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.3029 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.2355 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 11.899 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 63.928 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 49.644 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 266.64 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.8095 LAYER met4  ;
    ANTENNAMAXAREACAR 58.88 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 302.424 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.910273 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 165.6800 0.4850 165.8200 ;
    END
  END bot_FrameData[6]
  PIN bot_FrameData[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.5712 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.695 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 29.0802 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 156.496 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.8095 LAYER met3  ;
    ANTENNAMAXAREACAR 53.4409 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 266.088 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.967925 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 163.6400 0.4850 163.7800 ;
    END
  END bot_FrameData[5]
  PIN bot_FrameData[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2261 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.9695 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 18.0119 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 96.992 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 24.2655 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 132.704 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.8095 LAYER met4  ;
    ANTENNAMAXAREACAR 63.0634 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 320.757 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.826415 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 161.9400 0.4850 162.0800 ;
    END
  END bot_FrameData[4]
  PIN bot_FrameData[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2011 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.7175 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 31.0542 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 167.024 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.8095 LAYER met3  ;
    ANTENNAMAXAREACAR 46.9984 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 234.582 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.967925 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 160.2400 0.4850 160.3800 ;
    END
  END bot_FrameData[3]
  PIN bot_FrameData[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 6.9618 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 34.251 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 47.5069 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 229.899 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.967925 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 35.3374 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 189.864 LAYER met3  ;
    ANTENNAGATEAREA 1.6965 LAYER met3  ;
    ANTENNAMAXAREACAR 68.3365 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 341.814 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.991502 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.4848 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 3.056 LAYER met4  ;
    ANTENNAGATEAREA 2.8095 LAYER met4  ;
    ANTENNAMAXAREACAR 68.5091 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 342.902 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.991502 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 158.5400 0.4850 158.6800 ;
    END
  END bot_FrameData[2]
  PIN bot_FrameData[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 15.369 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 76.006 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.795 LAYER met2  ;
    ANTENNAMAXAREACAR 35.2931 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 171.284 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.515094 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 31.5132 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 169.472 LAYER met3  ;
    ANTENNAGATEAREA 2.8095 LAYER met3  ;
    ANTENNAMAXAREACAR 50.4418 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 251.045 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.967925 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 156.8400 0.4850 156.9800 ;
    END
  END bot_FrameData[1]
  PIN bot_FrameData[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 21.0062 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 103.754 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.113 LAYER met2  ;
    ANTENNAMAXAREACAR 40.9232 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 198.198 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.678167 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 38.4414 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 206.432 LAYER met3  ;
    ANTENNAGATEAREA 2.8095 LAYER met3  ;
    ANTENNAMAXAREACAR 54.6058 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 271.675 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.678167 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 155.1400 0.4850 155.2800 ;
    END
  END bot_FrameData[0]
  PIN bot_FrameData_O[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.0468 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.126 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 209.7350 209.5400 210.2200 209.6800 ;
    END
  END bot_FrameData_O[31]
  PIN bot_FrameData_O[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.1157 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.4705 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 209.7350 207.8400 210.2200 207.9800 ;
    END
  END bot_FrameData_O[30]
  PIN bot_FrameData_O[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.0468 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.126 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 209.7350 206.1400 210.2200 206.2800 ;
    END
  END bot_FrameData_O[29]
  PIN bot_FrameData_O[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.0468 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.126 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 209.7350 204.4400 210.2200 204.5800 ;
    END
  END bot_FrameData_O[28]
  PIN bot_FrameData_O[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.1938 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.861 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 209.7350 202.7400 210.2200 202.8800 ;
    END
  END bot_FrameData_O[27]
  PIN bot_FrameData_O[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.9869 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.8265 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 209.7350 201.0400 210.2200 201.1800 ;
    END
  END bot_FrameData_O[26]
  PIN bot_FrameData_O[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.0468 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.126 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 209.7350 199.0000 210.2200 199.1400 ;
    END
  END bot_FrameData_O[25]
  PIN bot_FrameData_O[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.1938 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.861 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 209.7350 197.3000 210.2200 197.4400 ;
    END
  END bot_FrameData_O[24]
  PIN bot_FrameData_O[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.1028 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 209.7350 195.6000 210.2200 195.7400 ;
    END
  END bot_FrameData_O[23]
  PIN bot_FrameData_O[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.5347 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.5655 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 209.7350 193.9000 210.2200 194.0400 ;
    END
  END bot_FrameData_O[22]
  PIN bot_FrameData_O[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.7489 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.6365 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 209.7350 192.2000 210.2200 192.3400 ;
    END
  END bot_FrameData_O[21]
  PIN bot_FrameData_O[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.9422 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.485 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 209.7350 190.1600 210.2200 190.3000 ;
    END
  END bot_FrameData_O[20]
  PIN bot_FrameData_O[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.2456 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.12 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 209.7350 188.4600 210.2200 188.6000 ;
    END
  END bot_FrameData_O[19]
  PIN bot_FrameData_O[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.7489 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.6365 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 209.7350 186.7600 210.2200 186.9000 ;
    END
  END bot_FrameData_O[18]
  PIN bot_FrameData_O[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.8432 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.99 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 209.7350 185.0600 210.2200 185.2000 ;
    END
  END bot_FrameData_O[17]
  PIN bot_FrameData_O[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 4.7249 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 23.5165 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 209.7350 183.3600 210.2200 183.5000 ;
    END
  END bot_FrameData_O[16]
  PIN bot_FrameData_O[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.8441 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.1125 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 209.7350 181.3200 210.2200 181.4600 ;
    END
  END bot_FrameData_O[15]
  PIN bot_FrameData_O[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.0468 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.126 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 209.7350 179.6200 210.2200 179.7600 ;
    END
  END bot_FrameData_O[14]
  PIN bot_FrameData_O[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1239 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.4585 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 59.887 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 319.864 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 15.5148 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 83.216 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 209.7350 177.9200 210.2200 178.0600 ;
    END
  END bot_FrameData_O[13]
  PIN bot_FrameData_O[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.6692 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.185 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 60.2298 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 321.696 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 209.7350 176.2200 210.2200 176.3600 ;
    END
  END bot_FrameData_O[12]
  PIN bot_FrameData_O[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.0468 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.126 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 209.7350 174.5200 210.2200 174.6600 ;
    END
  END bot_FrameData_O[11]
  PIN bot_FrameData_O[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.6061 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.9225 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 209.7350 172.4800 210.2200 172.6200 ;
    END
  END bot_FrameData_O[10]
  PIN bot_FrameData_O[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.1028 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 209.7350 170.7800 210.2200 170.9200 ;
    END
  END bot_FrameData_O[9]
  PIN bot_FrameData_O[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.2456 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.12 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 209.7350 169.0800 210.2200 169.2200 ;
    END
  END bot_FrameData_O[8]
  PIN bot_FrameData_O[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.6299 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.0415 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 209.7350 167.3800 210.2200 167.5200 ;
    END
  END bot_FrameData_O[7]
  PIN bot_FrameData_O[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.0468 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.126 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 209.7350 165.6800 210.2200 165.8200 ;
    END
  END bot_FrameData_O[6]
  PIN bot_FrameData_O[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2443 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.0605 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 25.8288 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 138.224 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 209.7350 163.6400 210.2200 163.7800 ;
    END
  END bot_FrameData_O[5]
  PIN bot_FrameData_O[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2261 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.9695 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 22.8888 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 122.544 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 209.7350 161.9400 210.2200 162.0800 ;
    END
  END bot_FrameData_O[4]
  PIN bot_FrameData_O[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2539 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.9905 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 11.737 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 63.064 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 0.9696 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 6.112 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 209.7350 160.2400 210.2200 160.3800 ;
    END
  END bot_FrameData_O[3]
  PIN bot_FrameData_O[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.4634 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.156 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 42.4338 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 226.784 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 209.7350 158.5400 210.2200 158.6800 ;
    END
  END bot_FrameData_O[2]
  PIN bot_FrameData_O[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2205 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.9415 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 8.0298 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 43.296 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 209.7350 156.8400 210.2200 156.9800 ;
    END
  END bot_FrameData_O[1]
  PIN bot_FrameData_O[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.1028 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 209.7350 155.1400 210.2200 155.2800 ;
    END
  END bot_FrameData_O[0]
  PIN FrameStrobe[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 12.6238 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 62.958 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 14.394 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 79.12 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met3  ;
    ANTENNAMAXAREACAR 24.4931 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 130.629 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.123098 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 199.8000 0.0000 199.9400 0.4850 ;
    END
  END FrameStrobe[19]
  PIN FrameStrobe[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.8731 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.2575 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 6.4101 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 30.6694 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 197.0400 0.0000 197.1800 0.4850 ;
    END
  END FrameStrobe[18]
  PIN FrameStrobe[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7307 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.5455 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 41.5993 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 205.869 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 194.7400 0.0000 194.8800 0.4850 ;
    END
  END FrameStrobe[17]
  PIN FrameStrobe[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.3343 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 21.5635 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 6.71178 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 32.1778 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 192.4400 0.0000 192.5800 0.4850 ;
    END
  END FrameStrobe[16]
  PIN FrameStrobe[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.1107 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 15.4455 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 4.7169 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 22.2034 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 190.1400 0.0000 190.2800 0.4850 ;
    END
  END FrameStrobe[15]
  PIN FrameStrobe[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 31.3754 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 155.89 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 6.1524 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 34.224 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met3  ;
    ANTENNAMAXAREACAR 9.20525 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 49.3138 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.123098 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 187.8400 0.0000 187.9800 0.4850 ;
    END
  END FrameStrobe[14]
  PIN FrameStrobe[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 25.6346 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 127.54 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 12.8604 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 72.352 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met3  ;
    ANTENNAMAXAREACAR 18.5623 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 102.187 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.123098 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 185.5400 0.0000 185.6800 0.4850 ;
    END
  END FrameStrobe[13]
  PIN FrameStrobe[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 25.1288 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 123.753 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.385 LAYER met2  ;
    ANTENNAMAXAREACAR 32.672 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 157.583 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.623061 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 17.9132 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 97.392 LAYER met3  ;
    ANTENNAGATEAREA 4.452 LAYER met3  ;
    ANTENNAMAXAREACAR 36.6957 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 179.459 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.985894 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 21.3306 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 114.704 LAYER met4  ;
    ANTENNAGATEAREA 5.2845 LAYER met4  ;
    ANTENNAMAXAREACAR 40.7321 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 201.165 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.985894 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 183.2400 0.0000 183.3800 0.4850 ;
    END
  END FrameStrobe[12]
  PIN FrameStrobe[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 14.3645 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 70.4235 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.59 LAYER met2  ;
    ANTENNAMAXAREACAR 27.6758 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 128.1 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.671698 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 15.8717 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 86.048 LAYER met3  ;
    ANTENNAGATEAREA 3.18 LAYER met3  ;
    ANTENNAMAXAREACAR 32.6669 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 155.159 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.728931 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 21.3951 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 115.984 LAYER met4  ;
    ANTENNAGATEAREA 5.2845 LAYER met4  ;
    ANTENNAMAXAREACAR 42.3201 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 209.062 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.826415 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 180.9400 0.0000 181.0800 0.4850 ;
    END
  END FrameStrobe[11]
  PIN FrameStrobe[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 36.8566 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 180.943 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.18 LAYER met2  ;
    ANTENNAMAXAREACAR 32.2065 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 154.319 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.12 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.644025 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 34.2984 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 184.336 LAYER met3  ;
    ANTENNAGATEAREA 5.2845 LAYER met3  ;
    ANTENNAMAXAREACAR 38.6969 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 189.201 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.644025 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 178.6400 0.0000 178.7800 0.4850 ;
    END
  END FrameStrobe[10]
  PIN FrameStrobe[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 42.8592 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 210.672 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 4.134 LAYER met2  ;
    ANTENNAMAXAREACAR 47.5782 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 226.936 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.625641 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 13.7136 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 74.08 LAYER met3  ;
    ANTENNAGATEAREA 5.2845 LAYER met3  ;
    ANTENNAMAXAREACAR 50.1732 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 240.954 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.625641 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 175.8800 0.0000 176.0200 0.4850 ;
    END
  END FrameStrobe[9]
  PIN FrameStrobe[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.133 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.504 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.1905 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.464 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 22.6836 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 121.92 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 5.2845 LAYER met4  ;
    ANTENNAMAXAREACAR 28.0537 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 128.973 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.723922 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 173.5800 0.0000 173.7200 0.4850 ;
    END
  END FrameStrobe[8]
  PIN FrameStrobe[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.4574 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.126 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.297 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 7.384 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 40.4988 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 216.464 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 5.2845 LAYER met4  ;
    ANTENNAMAXAREACAR 32.1163 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 154.972 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.621428 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 171.2800 0.0000 171.4200 0.4850 ;
    END
  END FrameStrobe[7]
  PIN FrameStrobe[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.3114 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 11.396 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 3.229 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 17.688 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 40.2213 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 215.92 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 5.2845 LAYER met4  ;
    ANTENNAMAXAREACAR 26.9138 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 132.398 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.725589 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 168.9800 0.0000 169.1200 0.4850 ;
    END
  END FrameStrobe[6]
  PIN FrameStrobe[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 54.0593 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 266.346 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 5.2845 LAYER met2  ;
    ANTENNAMAXAREACAR 25.0575 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 119.247 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.606289 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 166.6800 0.0000 166.8200 0.4850 ;
    END
  END FrameStrobe[5]
  PIN FrameStrobe[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 5.3691 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 26.3095 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.477 LAYER met2  ;
    ANTENNAMAXAREACAR 24.8201 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 117.993 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.548637 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 42.5486 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 228.8 LAYER met3  ;
    ANTENNAGATEAREA 3.18 LAYER met3  ;
    ANTENNAMAXAREACAR 50.571 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 251.756 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.601747 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 7.8126 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 42.608 LAYER met4  ;
    ANTENNAGATEAREA 5.2845 LAYER met4  ;
    ANTENNAMAXAREACAR 52.0494 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 259.819 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.853654 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 164.3800 0.0000 164.5200 0.4850 ;
    END
  END FrameStrobe[4]
  PIN FrameStrobe[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 20.6035 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 101.721 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.431 LAYER met2  ;
    ANTENNAMAXAREACAR 32.2131 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 151.47 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.662194 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 17.8946 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 97.312 LAYER met3  ;
    ANTENNAGATEAREA 2.544 LAYER met3  ;
    ANTENNAMAXAREACAR 39.2471 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 189.722 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.693641 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 28.1496 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 151.072 LAYER met4  ;
    ANTENNAGATEAREA 5.2845 LAYER met4  ;
    ANTENNAMAXAREACAR 44.5739 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 218.31 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.693641 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 162.0800 0.0000 162.2200 0.4850 ;
    END
  END FrameStrobe[3]
  PIN FrameStrobe[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 12.9373 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 62.9615 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.272 LAYER met2  ;
    ANTENNAMAXAREACAR 21.3048 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 100.184 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.527673 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 11.3728 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 61.592 LAYER met3  ;
    ANTENNAGATEAREA 1.908 LAYER met3  ;
    ANTENNAMAXAREACAR 27.2654 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 132.464 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.548637 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 44.3256 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 237.344 LAYER met4  ;
    ANTENNAGATEAREA 5.2845 LAYER met4  ;
    ANTENNAMAXAREACAR 39.6829 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 195.879 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.952201 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 159.7800 0.0000 159.9200 0.4850 ;
    END
  END FrameStrobe[2]
  PIN FrameStrobe[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.6134 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 17.906 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 15.7987 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 85.64 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.272 LAYER met3  ;
    ANTENNAMAXAREACAR 51.9951 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 254.925 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.695388 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 36.6222 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 197.2 LAYER met4  ;
    ANTENNAGATEAREA 5.2845 LAYER met4  ;
    ANTENNAMAXAREACAR 58.9252 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 292.241 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.695388 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 157.4800 0.0000 157.6200 0.4850 ;
    END
  END FrameStrobe[1]
  PIN FrameStrobe[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 43.5132 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 213.395 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 5.088 LAYER met2  ;
    ANTENNAMAXAREACAR 28.4666 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 132.793 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.614151 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 10.6968 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 57.52 LAYER met3  ;
    ANTENNAGATEAREA 5.2845 LAYER met3  ;
    ANTENNAMAXAREACAR 30.4908 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 143.678 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.614151 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 155.1800 0.0000 155.3200 0.4850 ;
    END
  END FrameStrobe[0]
  PIN FrameStrobe_O[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.9683 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.7335 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 199.8000 444.2350 199.9400 444.7200 ;
    END
  END FrameStrobe_O[19]
  PIN FrameStrobe_O[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.386 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.769 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.4 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.6 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 127.448 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 680.192 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 197.0400 444.2350 197.1800 444.7200 ;
    END
  END FrameStrobe_O[18]
  PIN FrameStrobe_O[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.7567 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.5575 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 194.7400 444.2350 194.8800 444.7200 ;
    END
  END FrameStrobe_O[17]
  PIN FrameStrobe_O[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.7163 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.4735 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 192.4400 444.2350 192.5800 444.7200 ;
    END
  END FrameStrobe_O[16]
  PIN FrameStrobe_O[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.9687 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.7355 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 190.1400 444.2350 190.2800 444.7200 ;
    END
  END FrameStrobe_O[15]
  PIN FrameStrobe_O[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.6995 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.3895 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 187.8400 444.2350 187.9800 444.7200 ;
    END
  END FrameStrobe_O[14]
  PIN FrameStrobe_O[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.6351 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.0675 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 185.0800 444.2350 185.2200 444.7200 ;
    END
  END FrameStrobe_O[13]
  PIN FrameStrobe_O[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 5.4907 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 27.3455 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 183.2400 444.2350 183.3800 444.7200 ;
    END
  END FrameStrobe_O[12]
  PIN FrameStrobe_O[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 5.7395 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 28.3535 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 180.4800 444.2350 180.6200 444.7200 ;
    END
  END FrameStrobe_O[11]
  PIN FrameStrobe_O[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 6.0983 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 30.3835 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 178.1800 444.2350 178.3200 444.7200 ;
    END
  END FrameStrobe_O[10]
  PIN FrameStrobe_O[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.1718 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.698 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 3.643 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 19.896 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 34.1886 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 183.28 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 175.8800 444.2350 176.0200 444.7200 ;
    END
  END FrameStrobe_O[9]
  PIN FrameStrobe_O[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.3041 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 11.2945 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 173.5800 444.2350 173.7200 444.7200 ;
    END
  END FrameStrobe_O[8]
  PIN FrameStrobe_O[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.3178 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.428 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.1905 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.464 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 20.7336 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 111.52 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 171.2800 444.2350 171.4200 444.7200 ;
    END
  END FrameStrobe_O[7]
  PIN FrameStrobe_O[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7448 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.563 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.366 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 7.752 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 38.3028 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 204.752 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 168.9800 444.2350 169.1200 444.7200 ;
    END
  END FrameStrobe_O[6]
  PIN FrameStrobe_O[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.9683 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.7335 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 166.6800 444.2350 166.8200 444.7200 ;
    END
  END FrameStrobe_O[5]
  PIN FrameStrobe_O[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.8493 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.1385 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 164.3800 444.2350 164.5200 444.7200 ;
    END
  END FrameStrobe_O[4]
  PIN FrameStrobe_O[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.5399 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.5915 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 162.0800 444.2350 162.2200 444.7200 ;
    END
  END FrameStrobe_O[3]
  PIN FrameStrobe_O[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.5899 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 12.8415 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 159.7800 444.2350 159.9200 444.7200 ;
    END
  END FrameStrobe_O[2]
  PIN FrameStrobe_O[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.7465 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 13.5065 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 157.4800 444.2350 157.6200 444.7200 ;
    END
  END FrameStrobe_O[1]
  PIN FrameStrobe_O[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7448 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.563 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.538 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 3.336 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 23.6148 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 126.416 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 155.1800 444.2350 155.3200 444.7200 ;
    END
  END FrameStrobe_O[0]
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;

# P/G power stripe data as pin
    PORT
      LAYER met3 ;
        RECT 5.5600 5.4300 204.6600 7.4300 ;
        RECT 5.5600 436.9500 204.6600 438.9500 ;
        RECT 5.5600 12.3400 7.5600 12.8200 ;
        RECT 5.5600 23.2200 7.5600 23.7000 ;
        RECT 5.5600 17.7800 7.5600 18.2600 ;
        RECT 5.5600 39.5400 7.5600 40.0200 ;
        RECT 5.5600 34.1000 7.5600 34.5800 ;
        RECT 5.5600 28.6600 7.5600 29.1400 ;
        RECT 5.5600 50.4200 7.5600 50.9000 ;
        RECT 5.5600 44.9800 7.5600 45.4600 ;
        RECT 5.5600 83.0600 7.5600 83.5400 ;
        RECT 5.5600 66.7400 7.5600 67.2200 ;
        RECT 5.5600 61.3000 7.5600 61.7800 ;
        RECT 5.5600 55.8600 7.5600 56.3400 ;
        RECT 5.5600 77.6200 7.5600 78.1000 ;
        RECT 5.5600 72.1800 7.5600 72.6600 ;
        RECT 5.5600 93.9400 7.5600 94.4200 ;
        RECT 5.5600 88.5000 7.5600 88.9800 ;
        RECT 5.5600 110.2600 7.5600 110.7400 ;
        RECT 5.5600 104.8200 7.5600 105.3000 ;
        RECT 5.5600 99.3800 7.5600 99.8600 ;
        RECT 5.5600 121.1400 7.5600 121.6200 ;
        RECT 5.5600 115.7000 7.5600 116.1800 ;
        RECT 5.5600 137.4600 7.5600 137.9400 ;
        RECT 5.5600 132.0200 7.5600 132.5000 ;
        RECT 5.5600 126.5800 7.5600 127.0600 ;
        RECT 5.5600 148.3400 7.5600 148.8200 ;
        RECT 5.5600 142.9000 7.5600 143.3800 ;
        RECT 5.5600 164.6600 7.5600 165.1400 ;
        RECT 5.5600 159.2200 7.5600 159.7000 ;
        RECT 5.5600 153.7800 7.5600 154.2600 ;
        RECT 5.5600 175.5400 7.5600 176.0200 ;
        RECT 5.5600 170.1000 7.5600 170.5800 ;
        RECT 5.5600 191.8600 7.5600 192.3400 ;
        RECT 5.5600 186.4200 7.5600 186.9000 ;
        RECT 5.5600 180.9800 7.5600 181.4600 ;
        RECT 5.5600 208.1800 7.5600 208.6600 ;
        RECT 5.5600 202.7400 7.5600 203.2200 ;
        RECT 5.5600 197.3000 7.5600 197.7800 ;
        RECT 5.5600 219.0600 7.5600 219.5400 ;
        RECT 5.5600 213.6200 7.5600 214.1000 ;
        RECT 202.6600 12.3400 204.6600 12.8200 ;
        RECT 202.6600 23.2200 204.6600 23.7000 ;
        RECT 202.6600 17.7800 204.6600 18.2600 ;
        RECT 202.6600 39.5400 204.6600 40.0200 ;
        RECT 202.6600 34.1000 204.6600 34.5800 ;
        RECT 202.6600 28.6600 204.6600 29.1400 ;
        RECT 202.6600 50.4200 204.6600 50.9000 ;
        RECT 202.6600 44.9800 204.6600 45.4600 ;
        RECT 202.6600 83.0600 204.6600 83.5400 ;
        RECT 202.6600 66.7400 204.6600 67.2200 ;
        RECT 202.6600 61.3000 204.6600 61.7800 ;
        RECT 202.6600 55.8600 204.6600 56.3400 ;
        RECT 202.6600 77.6200 204.6600 78.1000 ;
        RECT 202.6600 72.1800 204.6600 72.6600 ;
        RECT 202.6600 93.9400 204.6600 94.4200 ;
        RECT 202.6600 88.5000 204.6600 88.9800 ;
        RECT 202.6600 110.2600 204.6600 110.7400 ;
        RECT 202.6600 104.8200 204.6600 105.3000 ;
        RECT 202.6600 99.3800 204.6600 99.8600 ;
        RECT 202.6600 121.1400 204.6600 121.6200 ;
        RECT 202.6600 115.7000 204.6600 116.1800 ;
        RECT 202.6600 137.4600 204.6600 137.9400 ;
        RECT 202.6600 132.0200 204.6600 132.5000 ;
        RECT 202.6600 126.5800 204.6600 127.0600 ;
        RECT 202.6600 148.3400 204.6600 148.8200 ;
        RECT 202.6600 142.9000 204.6600 143.3800 ;
        RECT 202.6600 164.6600 204.6600 165.1400 ;
        RECT 202.6600 159.2200 204.6600 159.7000 ;
        RECT 202.6600 153.7800 204.6600 154.2600 ;
        RECT 202.6600 175.5400 204.6600 176.0200 ;
        RECT 202.6600 170.1000 204.6600 170.5800 ;
        RECT 202.6600 191.8600 204.6600 192.3400 ;
        RECT 202.6600 186.4200 204.6600 186.9000 ;
        RECT 202.6600 180.9800 204.6600 181.4600 ;
        RECT 202.6600 208.1800 204.6600 208.6600 ;
        RECT 202.6600 202.7400 204.6600 203.2200 ;
        RECT 202.6600 197.3000 204.6600 197.7800 ;
        RECT 202.6600 219.0600 204.6600 219.5400 ;
        RECT 202.6600 213.6200 204.6600 214.1000 ;
        RECT 5.5600 333.3000 7.5600 333.7800 ;
        RECT 5.5600 235.3800 7.5600 235.8600 ;
        RECT 5.5600 229.9400 7.5600 230.4200 ;
        RECT 5.5600 224.5000 7.5600 224.9800 ;
        RECT 5.5600 246.2600 7.5600 246.7400 ;
        RECT 5.5600 240.8200 7.5600 241.3000 ;
        RECT 5.5600 262.5800 7.5600 263.0600 ;
        RECT 5.5600 257.1400 7.5600 257.6200 ;
        RECT 5.5600 251.7000 7.5600 252.1800 ;
        RECT 5.5600 273.4600 7.5600 273.9400 ;
        RECT 5.5600 268.0200 7.5600 268.5000 ;
        RECT 5.5600 289.7800 7.5600 290.2600 ;
        RECT 5.5600 284.3400 7.5600 284.8200 ;
        RECT 5.5600 278.9000 7.5600 279.3800 ;
        RECT 5.5600 300.6600 7.5600 301.1400 ;
        RECT 5.5600 295.2200 7.5600 295.7000 ;
        RECT 5.5600 316.9800 7.5600 317.4600 ;
        RECT 5.5600 311.5400 7.5600 312.0200 ;
        RECT 5.5600 306.1000 7.5600 306.5800 ;
        RECT 5.5600 327.8600 7.5600 328.3400 ;
        RECT 5.5600 322.4200 7.5600 322.9000 ;
        RECT 5.5600 344.1800 7.5600 344.6600 ;
        RECT 5.5600 338.7400 7.5600 339.2200 ;
        RECT 5.5600 360.5000 7.5600 360.9800 ;
        RECT 5.5600 355.0600 7.5600 355.5400 ;
        RECT 5.5600 349.6200 7.5600 350.1000 ;
        RECT 5.5600 371.3800 7.5600 371.8600 ;
        RECT 5.5600 365.9400 7.5600 366.4200 ;
        RECT 5.5600 387.7000 7.5600 388.1800 ;
        RECT 5.5600 382.2600 7.5600 382.7400 ;
        RECT 5.5600 376.8200 7.5600 377.3000 ;
        RECT 5.5600 398.5800 7.5600 399.0600 ;
        RECT 5.5600 393.1400 7.5600 393.6200 ;
        RECT 5.5600 414.9000 7.5600 415.3800 ;
        RECT 5.5600 409.4600 7.5600 409.9400 ;
        RECT 5.5600 404.0200 7.5600 404.5000 ;
        RECT 5.5600 425.7800 7.5600 426.2600 ;
        RECT 5.5600 420.3400 7.5600 420.8200 ;
        RECT 5.5600 431.2200 7.5600 431.7000 ;
        RECT 202.6600 333.3000 204.6600 333.7800 ;
        RECT 202.6600 235.3800 204.6600 235.8600 ;
        RECT 202.6600 229.9400 204.6600 230.4200 ;
        RECT 202.6600 224.5000 204.6600 224.9800 ;
        RECT 202.6600 246.2600 204.6600 246.7400 ;
        RECT 202.6600 240.8200 204.6600 241.3000 ;
        RECT 202.6600 262.5800 204.6600 263.0600 ;
        RECT 202.6600 257.1400 204.6600 257.6200 ;
        RECT 202.6600 251.7000 204.6600 252.1800 ;
        RECT 202.6600 273.4600 204.6600 273.9400 ;
        RECT 202.6600 268.0200 204.6600 268.5000 ;
        RECT 202.6600 289.7800 204.6600 290.2600 ;
        RECT 202.6600 284.3400 204.6600 284.8200 ;
        RECT 202.6600 278.9000 204.6600 279.3800 ;
        RECT 202.6600 300.6600 204.6600 301.1400 ;
        RECT 202.6600 295.2200 204.6600 295.7000 ;
        RECT 202.6600 316.9800 204.6600 317.4600 ;
        RECT 202.6600 311.5400 204.6600 312.0200 ;
        RECT 202.6600 306.1000 204.6600 306.5800 ;
        RECT 202.6600 327.8600 204.6600 328.3400 ;
        RECT 202.6600 322.4200 204.6600 322.9000 ;
        RECT 202.6600 344.1800 204.6600 344.6600 ;
        RECT 202.6600 338.7400 204.6600 339.2200 ;
        RECT 202.6600 360.5000 204.6600 360.9800 ;
        RECT 202.6600 355.0600 204.6600 355.5400 ;
        RECT 202.6600 349.6200 204.6600 350.1000 ;
        RECT 202.6600 371.3800 204.6600 371.8600 ;
        RECT 202.6600 365.9400 204.6600 366.4200 ;
        RECT 202.6600 387.7000 204.6600 388.1800 ;
        RECT 202.6600 382.2600 204.6600 382.7400 ;
        RECT 202.6600 376.8200 204.6600 377.3000 ;
        RECT 202.6600 398.5800 204.6600 399.0600 ;
        RECT 202.6600 393.1400 204.6600 393.6200 ;
        RECT 202.6600 414.9000 204.6600 415.3800 ;
        RECT 202.6600 409.4600 204.6600 409.9400 ;
        RECT 202.6600 404.0200 204.6600 404.5000 ;
        RECT 202.6600 425.7800 204.6600 426.2600 ;
        RECT 202.6600 420.3400 204.6600 420.8200 ;
        RECT 202.6600 431.2200 204.6600 431.7000 ;
      LAYER met4 ;
        RECT 5.5600 5.4300 7.5600 438.9500 ;
        RECT 202.6600 5.4300 204.6600 438.9500 ;
        RECT 10.1200 5.4300 11.7200 438.9500 ;
        RECT 55.1200 5.4300 56.7200 438.9500 ;
        RECT 100.1200 5.4300 101.7200 438.9500 ;
        RECT 145.1200 5.4300 146.7200 438.9500 ;
        RECT 190.1200 5.4300 191.7200 438.9500 ;
    END
# end of P/G power stripe data as pin

  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;

# P/G power stripe data as pin
    PORT
      LAYER met3 ;
        RECT 2.5600 2.4300 207.6600 4.4300 ;
        RECT 2.5600 439.9500 207.6600 441.9500 ;
        RECT 2.5600 9.6200 4.5600 10.1000 ;
        RECT 2.5600 25.9400 4.5600 26.4200 ;
        RECT 2.5600 20.5000 4.5600 20.9800 ;
        RECT 2.5600 15.0600 4.5600 15.5400 ;
        RECT 2.5600 36.8200 4.5600 37.3000 ;
        RECT 2.5600 31.3800 4.5600 31.8600 ;
        RECT 2.5600 53.1400 4.5600 53.6200 ;
        RECT 2.5600 47.7000 4.5600 48.1800 ;
        RECT 2.5600 42.2600 4.5600 42.7400 ;
        RECT 2.5600 69.4600 4.5600 69.9400 ;
        RECT 2.5600 64.0200 4.5600 64.5000 ;
        RECT 2.5600 58.5800 4.5600 59.0600 ;
        RECT 2.5600 80.3400 4.5600 80.8200 ;
        RECT 2.5600 74.9000 4.5600 75.3800 ;
        RECT 2.5600 96.6600 4.5600 97.1400 ;
        RECT 2.5600 91.2200 4.5600 91.7000 ;
        RECT 2.5600 85.7800 4.5600 86.2600 ;
        RECT 2.5600 107.5400 4.5600 108.0200 ;
        RECT 2.5600 102.1000 4.5600 102.5800 ;
        RECT 2.5600 123.8600 4.5600 124.3400 ;
        RECT 2.5600 118.4200 4.5600 118.9000 ;
        RECT 2.5600 112.9800 4.5600 113.4600 ;
        RECT 2.5600 134.7400 4.5600 135.2200 ;
        RECT 2.5600 129.3000 4.5600 129.7800 ;
        RECT 2.5600 151.0600 4.5600 151.5400 ;
        RECT 2.5600 145.6200 4.5600 146.1000 ;
        RECT 2.5600 140.1800 4.5600 140.6600 ;
        RECT 2.5600 161.9400 4.5600 162.4200 ;
        RECT 2.5600 156.5000 4.5600 156.9800 ;
        RECT 2.5600 178.2600 4.5600 178.7400 ;
        RECT 2.5600 172.8200 4.5600 173.3000 ;
        RECT 2.5600 167.3800 4.5600 167.8600 ;
        RECT 2.5600 189.1400 4.5600 189.6200 ;
        RECT 2.5600 183.7000 4.5600 184.1800 ;
        RECT 2.5600 205.4600 4.5600 205.9400 ;
        RECT 2.5600 200.0200 4.5600 200.5000 ;
        RECT 2.5600 194.5800 4.5600 195.0600 ;
        RECT 2.5600 221.7800 4.5600 222.2600 ;
        RECT 2.5600 216.3400 4.5600 216.8200 ;
        RECT 2.5600 210.9000 4.5600 211.3800 ;
        RECT 205.6600 9.6200 207.6600 10.1000 ;
        RECT 205.6600 25.9400 207.6600 26.4200 ;
        RECT 205.6600 20.5000 207.6600 20.9800 ;
        RECT 205.6600 15.0600 207.6600 15.5400 ;
        RECT 205.6600 36.8200 207.6600 37.3000 ;
        RECT 205.6600 31.3800 207.6600 31.8600 ;
        RECT 205.6600 53.1400 207.6600 53.6200 ;
        RECT 205.6600 47.7000 207.6600 48.1800 ;
        RECT 205.6600 42.2600 207.6600 42.7400 ;
        RECT 205.6600 69.4600 207.6600 69.9400 ;
        RECT 205.6600 64.0200 207.6600 64.5000 ;
        RECT 205.6600 58.5800 207.6600 59.0600 ;
        RECT 205.6600 80.3400 207.6600 80.8200 ;
        RECT 205.6600 74.9000 207.6600 75.3800 ;
        RECT 205.6600 96.6600 207.6600 97.1400 ;
        RECT 205.6600 91.2200 207.6600 91.7000 ;
        RECT 205.6600 85.7800 207.6600 86.2600 ;
        RECT 205.6600 107.5400 207.6600 108.0200 ;
        RECT 205.6600 102.1000 207.6600 102.5800 ;
        RECT 205.6600 123.8600 207.6600 124.3400 ;
        RECT 205.6600 118.4200 207.6600 118.9000 ;
        RECT 205.6600 112.9800 207.6600 113.4600 ;
        RECT 205.6600 134.7400 207.6600 135.2200 ;
        RECT 205.6600 129.3000 207.6600 129.7800 ;
        RECT 205.6600 151.0600 207.6600 151.5400 ;
        RECT 205.6600 145.6200 207.6600 146.1000 ;
        RECT 205.6600 140.1800 207.6600 140.6600 ;
        RECT 205.6600 161.9400 207.6600 162.4200 ;
        RECT 205.6600 156.5000 207.6600 156.9800 ;
        RECT 205.6600 178.2600 207.6600 178.7400 ;
        RECT 205.6600 172.8200 207.6600 173.3000 ;
        RECT 205.6600 167.3800 207.6600 167.8600 ;
        RECT 205.6600 189.1400 207.6600 189.6200 ;
        RECT 205.6600 183.7000 207.6600 184.1800 ;
        RECT 205.6600 205.4600 207.6600 205.9400 ;
        RECT 205.6600 200.0200 207.6600 200.5000 ;
        RECT 205.6600 194.5800 207.6600 195.0600 ;
        RECT 205.6600 221.7800 207.6600 222.2600 ;
        RECT 205.6600 216.3400 207.6600 216.8200 ;
        RECT 205.6600 210.9000 207.6600 211.3800 ;
        RECT 2.5600 232.6600 4.5600 233.1400 ;
        RECT 2.5600 227.2200 4.5600 227.7000 ;
        RECT 2.5600 248.9800 4.5600 249.4600 ;
        RECT 2.5600 243.5400 4.5600 244.0200 ;
        RECT 2.5600 238.1000 4.5600 238.5800 ;
        RECT 2.5600 259.8600 4.5600 260.3400 ;
        RECT 2.5600 254.4200 4.5600 254.9000 ;
        RECT 2.5600 276.1800 4.5600 276.6600 ;
        RECT 2.5600 270.7400 4.5600 271.2200 ;
        RECT 2.5600 265.3000 4.5600 265.7800 ;
        RECT 2.5600 287.0600 4.5600 287.5400 ;
        RECT 2.5600 281.6200 4.5600 282.1000 ;
        RECT 2.5600 303.3800 4.5600 303.8600 ;
        RECT 2.5600 297.9400 4.5600 298.4200 ;
        RECT 2.5600 292.5000 4.5600 292.9800 ;
        RECT 2.5600 314.2600 4.5600 314.7400 ;
        RECT 2.5600 308.8200 4.5600 309.3000 ;
        RECT 2.5600 330.5800 4.5600 331.0600 ;
        RECT 2.5600 325.1400 4.5600 325.6200 ;
        RECT 2.5600 319.7000 4.5600 320.1800 ;
        RECT 2.5600 346.9000 4.5600 347.3800 ;
        RECT 2.5600 341.4600 4.5600 341.9400 ;
        RECT 2.5600 336.0200 4.5600 336.5000 ;
        RECT 2.5600 357.7800 4.5600 358.2600 ;
        RECT 2.5600 352.3400 4.5600 352.8200 ;
        RECT 2.5600 374.1000 4.5600 374.5800 ;
        RECT 2.5600 368.6600 4.5600 369.1400 ;
        RECT 2.5600 363.2200 4.5600 363.7000 ;
        RECT 2.5600 384.9800 4.5600 385.4600 ;
        RECT 2.5600 379.5400 4.5600 380.0200 ;
        RECT 2.5600 401.3000 4.5600 401.7800 ;
        RECT 2.5600 395.8600 4.5600 396.3400 ;
        RECT 2.5600 390.4200 4.5600 390.9000 ;
        RECT 2.5600 412.1800 4.5600 412.6600 ;
        RECT 2.5600 406.7400 4.5600 407.2200 ;
        RECT 2.5600 428.5000 4.5600 428.9800 ;
        RECT 2.5600 423.0600 4.5600 423.5400 ;
        RECT 2.5600 417.6200 4.5600 418.1000 ;
        RECT 2.5600 433.9400 4.5600 434.4200 ;
        RECT 205.6600 232.6600 207.6600 233.1400 ;
        RECT 205.6600 227.2200 207.6600 227.7000 ;
        RECT 205.6600 248.9800 207.6600 249.4600 ;
        RECT 205.6600 243.5400 207.6600 244.0200 ;
        RECT 205.6600 238.1000 207.6600 238.5800 ;
        RECT 205.6600 259.8600 207.6600 260.3400 ;
        RECT 205.6600 254.4200 207.6600 254.9000 ;
        RECT 205.6600 276.1800 207.6600 276.6600 ;
        RECT 205.6600 270.7400 207.6600 271.2200 ;
        RECT 205.6600 265.3000 207.6600 265.7800 ;
        RECT 205.6600 287.0600 207.6600 287.5400 ;
        RECT 205.6600 281.6200 207.6600 282.1000 ;
        RECT 205.6600 303.3800 207.6600 303.8600 ;
        RECT 205.6600 297.9400 207.6600 298.4200 ;
        RECT 205.6600 292.5000 207.6600 292.9800 ;
        RECT 205.6600 314.2600 207.6600 314.7400 ;
        RECT 205.6600 308.8200 207.6600 309.3000 ;
        RECT 205.6600 330.5800 207.6600 331.0600 ;
        RECT 205.6600 325.1400 207.6600 325.6200 ;
        RECT 205.6600 319.7000 207.6600 320.1800 ;
        RECT 205.6600 346.9000 207.6600 347.3800 ;
        RECT 205.6600 341.4600 207.6600 341.9400 ;
        RECT 205.6600 336.0200 207.6600 336.5000 ;
        RECT 205.6600 357.7800 207.6600 358.2600 ;
        RECT 205.6600 352.3400 207.6600 352.8200 ;
        RECT 205.6600 374.1000 207.6600 374.5800 ;
        RECT 205.6600 368.6600 207.6600 369.1400 ;
        RECT 205.6600 363.2200 207.6600 363.7000 ;
        RECT 205.6600 384.9800 207.6600 385.4600 ;
        RECT 205.6600 379.5400 207.6600 380.0200 ;
        RECT 205.6600 401.3000 207.6600 401.7800 ;
        RECT 205.6600 395.8600 207.6600 396.3400 ;
        RECT 205.6600 390.4200 207.6600 390.9000 ;
        RECT 205.6600 412.1800 207.6600 412.6600 ;
        RECT 205.6600 406.7400 207.6600 407.2200 ;
        RECT 205.6600 428.5000 207.6600 428.9800 ;
        RECT 205.6600 423.0600 207.6600 423.5400 ;
        RECT 205.6600 417.6200 207.6600 418.1000 ;
        RECT 205.6600 433.9400 207.6600 434.4200 ;
      LAYER met4 ;
        RECT 2.5600 2.4300 4.5600 441.9500 ;
        RECT 205.6600 2.4300 207.6600 441.9500 ;
        RECT 13.3200 2.4300 14.9200 441.9500 ;
        RECT 58.3200 2.4300 59.9200 441.9500 ;
        RECT 103.3200 2.4300 104.9200 441.9500 ;
        RECT 148.3200 2.4300 149.9200 441.9500 ;
        RECT 193.3200 2.4300 194.9200 441.9500 ;
    END
# end of P/G power stripe data as pin

  END VPWR
  OBS
    LAYER li1 ;
      RECT 149.5250 444.2200 210.2200 444.7200 ;
      RECT 148.6050 444.2200 149.0150 444.7200 ;
      RECT 147.2250 444.2200 148.0950 444.7200 ;
      RECT 145.8450 444.2200 146.7150 444.7200 ;
      RECT 144.4650 444.2200 145.3350 444.7200 ;
      RECT 143.0850 444.2200 143.9550 444.7200 ;
      RECT 141.7050 444.2200 142.5750 444.7200 ;
      RECT 140.3250 444.2200 141.1950 444.7200 ;
      RECT 138.9450 444.2200 139.8150 444.7200 ;
      RECT 137.5650 444.2200 138.4350 444.7200 ;
      RECT 136.1850 444.2200 137.0550 444.7200 ;
      RECT 134.8050 444.2200 135.6750 444.7200 ;
      RECT 133.4250 444.2200 134.2950 444.7200 ;
      RECT 132.0450 444.2200 132.9150 444.7200 ;
      RECT 130.6650 444.2200 131.5350 444.7200 ;
      RECT 129.2850 444.2200 130.1550 444.7200 ;
      RECT 127.9050 444.2200 128.7750 444.7200 ;
      RECT 126.5250 444.2200 127.3950 444.7200 ;
      RECT 125.6050 444.2200 126.0150 444.7200 ;
      RECT 124.2250 444.2200 125.0950 444.7200 ;
      RECT 122.8450 444.2200 123.7150 444.7200 ;
      RECT 121.4650 444.2200 122.3350 444.7200 ;
      RECT 120.0850 444.2200 120.9550 444.7200 ;
      RECT 118.7050 444.2200 119.5750 444.7200 ;
      RECT 117.3250 444.2200 118.1950 444.7200 ;
      RECT 115.9450 444.2200 116.8150 444.7200 ;
      RECT 114.5650 444.2200 115.4350 444.7200 ;
      RECT 113.1850 444.2200 114.0550 444.7200 ;
      RECT 111.8050 444.2200 112.6750 444.7200 ;
      RECT 110.4250 444.2200 111.2950 444.7200 ;
      RECT 109.0450 444.2200 109.9150 444.7200 ;
      RECT 107.6650 444.2200 108.5350 444.7200 ;
      RECT 106.2850 444.2200 107.1550 444.7200 ;
      RECT 104.9050 444.2200 105.7750 444.7200 ;
      RECT 103.5250 444.2200 104.3950 444.7200 ;
      RECT 102.6050 444.2200 103.0150 444.7200 ;
      RECT 101.2250 444.2200 102.0950 444.7200 ;
      RECT 99.8450 444.2200 100.7150 444.7200 ;
      RECT 98.4650 444.2200 99.3350 444.7200 ;
      RECT 97.0850 444.2200 97.9550 444.7200 ;
      RECT 95.7050 444.2200 96.5750 444.7200 ;
      RECT 94.3250 444.2200 95.1950 444.7200 ;
      RECT 92.9450 444.2200 93.8150 444.7200 ;
      RECT 91.5650 444.2200 92.4350 444.7200 ;
      RECT 90.1850 444.2200 91.0550 444.7200 ;
      RECT 88.8050 444.2200 89.6750 444.7200 ;
      RECT 87.4250 444.2200 88.2950 444.7200 ;
      RECT 86.0450 444.2200 86.9150 444.7200 ;
      RECT 84.6650 444.2200 85.5350 444.7200 ;
      RECT 83.2850 444.2200 84.1550 444.7200 ;
      RECT 81.9050 444.2200 82.7750 444.7200 ;
      RECT 80.5250 444.2200 81.3950 444.7200 ;
      RECT 79.6050 444.2200 80.0150 444.7200 ;
      RECT 78.2250 444.2200 79.0950 444.7200 ;
      RECT 76.8450 444.2200 77.7150 444.7200 ;
      RECT 75.4650 444.2200 76.3350 444.7200 ;
      RECT 74.0850 444.2200 74.9550 444.7200 ;
      RECT 72.7050 444.2200 73.5750 444.7200 ;
      RECT 71.3250 444.2200 72.1950 444.7200 ;
      RECT 69.9450 444.2200 70.8150 444.7200 ;
      RECT 68.5650 444.2200 69.4350 444.7200 ;
      RECT 67.1850 444.2200 68.0550 444.7200 ;
      RECT 65.8050 444.2200 66.6750 444.7200 ;
      RECT 64.4250 444.2200 65.2950 444.7200 ;
      RECT 63.0450 444.2200 63.9150 444.7200 ;
      RECT 61.6650 444.2200 62.5350 444.7200 ;
      RECT 60.2850 444.2200 61.1550 444.7200 ;
      RECT 58.9050 444.2200 59.7750 444.7200 ;
      RECT 57.5250 444.2200 58.3950 444.7200 ;
      RECT 56.6050 444.2200 57.0150 444.7200 ;
      RECT 55.2250 444.2200 56.0950 444.7200 ;
      RECT 53.8450 444.2200 54.7150 444.7200 ;
      RECT 52.4650 444.2200 53.3350 444.7200 ;
      RECT 51.0850 444.2200 51.9550 444.7200 ;
      RECT 49.7050 444.2200 50.5750 444.7200 ;
      RECT 48.3250 444.2200 49.1950 444.7200 ;
      RECT 46.9450 444.2200 47.8150 444.7200 ;
      RECT 45.5650 444.2200 46.4350 444.7200 ;
      RECT 44.1850 444.2200 45.0550 444.7200 ;
      RECT 42.8050 444.2200 43.6750 444.7200 ;
      RECT 41.4250 444.2200 42.2950 444.7200 ;
      RECT 40.0450 444.2200 40.9150 444.7200 ;
      RECT 38.6650 444.2200 39.5350 444.7200 ;
      RECT 37.2850 444.2200 38.1550 444.7200 ;
      RECT 35.9050 444.2200 36.7750 444.7200 ;
      RECT 34.5250 444.2200 35.3950 444.7200 ;
      RECT 33.6050 444.2200 34.0150 444.7200 ;
      RECT 32.2250 444.2200 33.0950 444.7200 ;
      RECT 30.8450 444.2200 31.7150 444.7200 ;
      RECT 29.4650 444.2200 30.3350 444.7200 ;
      RECT 28.0850 444.2200 28.9550 444.7200 ;
      RECT 26.7050 444.2200 27.5750 444.7200 ;
      RECT 25.3250 444.2200 26.1950 444.7200 ;
      RECT 23.9450 444.2200 24.8150 444.7200 ;
      RECT 22.5650 444.2200 23.4350 444.7200 ;
      RECT 21.1850 444.2200 22.0550 444.7200 ;
      RECT 19.8050 444.2200 20.6750 444.7200 ;
      RECT 18.4250 444.2200 19.2950 444.7200 ;
      RECT 17.0450 444.2200 17.9150 444.7200 ;
      RECT 15.6650 444.2200 16.5350 444.7200 ;
      RECT 14.2850 444.2200 15.1550 444.7200 ;
      RECT 12.9050 444.2200 13.7750 444.7200 ;
      RECT 11.5250 444.2200 12.3950 444.7200 ;
      RECT 10.6050 444.2200 11.0150 444.7200 ;
      RECT 0.0000 444.2200 10.0950 444.7200 ;
      RECT 0.0000 0.5000 210.2200 444.2200 ;
      RECT 149.5250 0.0000 210.2200 0.5000 ;
      RECT 148.6050 0.0000 149.0150 0.5000 ;
      RECT 147.2250 0.0000 148.0950 0.5000 ;
      RECT 145.8450 0.0000 146.7150 0.5000 ;
      RECT 144.4650 0.0000 145.3350 0.5000 ;
      RECT 143.0850 0.0000 143.9550 0.5000 ;
      RECT 141.7050 0.0000 142.5750 0.5000 ;
      RECT 140.3250 0.0000 141.1950 0.5000 ;
      RECT 138.9450 0.0000 139.8150 0.5000 ;
      RECT 137.5650 0.0000 138.4350 0.5000 ;
      RECT 136.1850 0.0000 137.0550 0.5000 ;
      RECT 134.8050 0.0000 135.6750 0.5000 ;
      RECT 133.4250 0.0000 134.2950 0.5000 ;
      RECT 132.0450 0.0000 132.9150 0.5000 ;
      RECT 130.6650 0.0000 131.5350 0.5000 ;
      RECT 129.2850 0.0000 130.1550 0.5000 ;
      RECT 127.9050 0.0000 128.7750 0.5000 ;
      RECT 126.5250 0.0000 127.3950 0.5000 ;
      RECT 125.6050 0.0000 126.0150 0.5000 ;
      RECT 124.2250 0.0000 125.0950 0.5000 ;
      RECT 122.8450 0.0000 123.7150 0.5000 ;
      RECT 121.4650 0.0000 122.3350 0.5000 ;
      RECT 120.0850 0.0000 120.9550 0.5000 ;
      RECT 118.7050 0.0000 119.5750 0.5000 ;
      RECT 117.3250 0.0000 118.1950 0.5000 ;
      RECT 115.9450 0.0000 116.8150 0.5000 ;
      RECT 114.5650 0.0000 115.4350 0.5000 ;
      RECT 113.1850 0.0000 114.0550 0.5000 ;
      RECT 111.8050 0.0000 112.6750 0.5000 ;
      RECT 110.4250 0.0000 111.2950 0.5000 ;
      RECT 109.0450 0.0000 109.9150 0.5000 ;
      RECT 107.6650 0.0000 108.5350 0.5000 ;
      RECT 106.2850 0.0000 107.1550 0.5000 ;
      RECT 104.9050 0.0000 105.7750 0.5000 ;
      RECT 103.5250 0.0000 104.3950 0.5000 ;
      RECT 102.6050 0.0000 103.0150 0.5000 ;
      RECT 101.2250 0.0000 102.0950 0.5000 ;
      RECT 99.8450 0.0000 100.7150 0.5000 ;
      RECT 98.4650 0.0000 99.3350 0.5000 ;
      RECT 97.0850 0.0000 97.9550 0.5000 ;
      RECT 95.7050 0.0000 96.5750 0.5000 ;
      RECT 94.3250 0.0000 95.1950 0.5000 ;
      RECT 92.9450 0.0000 93.8150 0.5000 ;
      RECT 91.5650 0.0000 92.4350 0.5000 ;
      RECT 90.1850 0.0000 91.0550 0.5000 ;
      RECT 88.8050 0.0000 89.6750 0.5000 ;
      RECT 87.4250 0.0000 88.2950 0.5000 ;
      RECT 86.0450 0.0000 86.9150 0.5000 ;
      RECT 84.6650 0.0000 85.5350 0.5000 ;
      RECT 83.2850 0.0000 84.1550 0.5000 ;
      RECT 81.9050 0.0000 82.7750 0.5000 ;
      RECT 80.5250 0.0000 81.3950 0.5000 ;
      RECT 79.6050 0.0000 80.0150 0.5000 ;
      RECT 78.2250 0.0000 79.0950 0.5000 ;
      RECT 76.8450 0.0000 77.7150 0.5000 ;
      RECT 75.4650 0.0000 76.3350 0.5000 ;
      RECT 74.0850 0.0000 74.9550 0.5000 ;
      RECT 72.7050 0.0000 73.5750 0.5000 ;
      RECT 71.3250 0.0000 72.1950 0.5000 ;
      RECT 69.9450 0.0000 70.8150 0.5000 ;
      RECT 68.5650 0.0000 69.4350 0.5000 ;
      RECT 67.1850 0.0000 68.0550 0.5000 ;
      RECT 65.8050 0.0000 66.6750 0.5000 ;
      RECT 64.4250 0.0000 65.2950 0.5000 ;
      RECT 63.0450 0.0000 63.9150 0.5000 ;
      RECT 61.6650 0.0000 62.5350 0.5000 ;
      RECT 60.2850 0.0000 61.1550 0.5000 ;
      RECT 58.9050 0.0000 59.7750 0.5000 ;
      RECT 57.5250 0.0000 58.3950 0.5000 ;
      RECT 56.6050 0.0000 57.0150 0.5000 ;
      RECT 55.2250 0.0000 56.0950 0.5000 ;
      RECT 53.8450 0.0000 54.7150 0.5000 ;
      RECT 52.4650 0.0000 53.3350 0.5000 ;
      RECT 51.0850 0.0000 51.9550 0.5000 ;
      RECT 49.7050 0.0000 50.5750 0.5000 ;
      RECT 48.3250 0.0000 49.1950 0.5000 ;
      RECT 46.9450 0.0000 47.8150 0.5000 ;
      RECT 45.5650 0.0000 46.4350 0.5000 ;
      RECT 44.1850 0.0000 45.0550 0.5000 ;
      RECT 42.8050 0.0000 43.6750 0.5000 ;
      RECT 41.4250 0.0000 42.2950 0.5000 ;
      RECT 40.0450 0.0000 40.9150 0.5000 ;
      RECT 38.6650 0.0000 39.5350 0.5000 ;
      RECT 37.2850 0.0000 38.1550 0.5000 ;
      RECT 35.9050 0.0000 36.7750 0.5000 ;
      RECT 34.5250 0.0000 35.3950 0.5000 ;
      RECT 33.6050 0.0000 34.0150 0.5000 ;
      RECT 32.2250 0.0000 33.0950 0.5000 ;
      RECT 30.8450 0.0000 31.7150 0.5000 ;
      RECT 29.4650 0.0000 30.3350 0.5000 ;
      RECT 28.0850 0.0000 28.9550 0.5000 ;
      RECT 26.7050 0.0000 27.5750 0.5000 ;
      RECT 25.3250 0.0000 26.1950 0.5000 ;
      RECT 23.9450 0.0000 24.8150 0.5000 ;
      RECT 22.5650 0.0000 23.4350 0.5000 ;
      RECT 21.1850 0.0000 22.0550 0.5000 ;
      RECT 19.8050 0.0000 20.6750 0.5000 ;
      RECT 18.4250 0.0000 19.2950 0.5000 ;
      RECT 17.0450 0.0000 17.9150 0.5000 ;
      RECT 15.6650 0.0000 16.5350 0.5000 ;
      RECT 14.2850 0.0000 15.1550 0.5000 ;
      RECT 12.9050 0.0000 13.7750 0.5000 ;
      RECT 11.5250 0.0000 12.3950 0.5000 ;
      RECT 10.6050 0.0000 11.0150 0.5000 ;
      RECT 0.0000 0.0000 10.0950 0.5000 ;
    LAYER met1 ;
      RECT 0.0000 0.0000 210.2200 444.7200 ;
    LAYER met2 ;
      RECT 200.0800 444.0950 210.2200 444.7200 ;
      RECT 197.3200 444.0950 199.6600 444.7200 ;
      RECT 195.0200 444.0950 196.9000 444.7200 ;
      RECT 192.7200 444.0950 194.6000 444.7200 ;
      RECT 190.4200 444.0950 192.3000 444.7200 ;
      RECT 188.1200 444.0950 190.0000 444.7200 ;
      RECT 185.3600 444.0950 187.7000 444.7200 ;
      RECT 183.5200 444.0950 184.9400 444.7200 ;
      RECT 180.7600 444.0950 183.1000 444.7200 ;
      RECT 178.4600 444.0950 180.3400 444.7200 ;
      RECT 176.1600 444.0950 178.0400 444.7200 ;
      RECT 173.8600 444.0950 175.7400 444.7200 ;
      RECT 171.5600 444.0950 173.4400 444.7200 ;
      RECT 169.2600 444.0950 171.1400 444.7200 ;
      RECT 166.9600 444.0950 168.8400 444.7200 ;
      RECT 164.6600 444.0950 166.5400 444.7200 ;
      RECT 162.3600 444.0950 164.2400 444.7200 ;
      RECT 160.0600 444.0950 161.9400 444.7200 ;
      RECT 157.7600 444.0950 159.6400 444.7200 ;
      RECT 155.4600 444.0950 157.3400 444.7200 ;
      RECT 0.0000 444.0950 155.0400 444.7200 ;
      RECT 0.0000 434.5600 210.2200 444.0950 ;
      RECT 0.6250 434.1400 209.5950 434.5600 ;
      RECT 0.0000 432.8600 210.2200 434.1400 ;
      RECT 0.6250 432.4400 209.5950 432.8600 ;
      RECT 0.0000 431.1600 210.2200 432.4400 ;
      RECT 0.6250 430.7400 209.5950 431.1600 ;
      RECT 0.0000 429.4600 210.2200 430.7400 ;
      RECT 0.6250 429.0400 209.5950 429.4600 ;
      RECT 0.0000 427.7600 210.2200 429.0400 ;
      RECT 0.6250 427.3400 209.5950 427.7600 ;
      RECT 0.0000 426.0600 210.2200 427.3400 ;
      RECT 0.6250 425.6400 209.5950 426.0600 ;
      RECT 0.0000 424.3600 210.2200 425.6400 ;
      RECT 0.6250 423.9400 209.5950 424.3600 ;
      RECT 0.0000 422.3200 210.2200 423.9400 ;
      RECT 0.6250 421.9000 209.5950 422.3200 ;
      RECT 0.0000 420.6200 210.2200 421.9000 ;
      RECT 0.6250 420.2000 209.5950 420.6200 ;
      RECT 0.0000 418.9200 210.2200 420.2000 ;
      RECT 0.6250 418.5000 209.5950 418.9200 ;
      RECT 0.0000 417.2200 210.2200 418.5000 ;
      RECT 0.6250 416.8000 209.5950 417.2200 ;
      RECT 0.0000 415.5200 210.2200 416.8000 ;
      RECT 0.6250 415.1000 209.5950 415.5200 ;
      RECT 0.0000 413.8200 210.2200 415.1000 ;
      RECT 0.6250 413.4000 209.5950 413.8200 ;
      RECT 0.0000 411.7800 210.2200 413.4000 ;
      RECT 0.6250 411.3600 209.5950 411.7800 ;
      RECT 0.0000 410.0800 210.2200 411.3600 ;
      RECT 0.6250 409.6600 209.5950 410.0800 ;
      RECT 0.0000 408.3800 210.2200 409.6600 ;
      RECT 0.6250 407.9600 209.5950 408.3800 ;
      RECT 0.0000 406.6800 210.2200 407.9600 ;
      RECT 0.6250 406.2600 209.5950 406.6800 ;
      RECT 0.0000 404.9800 210.2200 406.2600 ;
      RECT 0.6250 404.5600 209.5950 404.9800 ;
      RECT 0.0000 403.2800 210.2200 404.5600 ;
      RECT 0.6250 402.8600 209.5950 403.2800 ;
      RECT 0.0000 401.2400 210.2200 402.8600 ;
      RECT 0.6250 400.8200 209.5950 401.2400 ;
      RECT 0.0000 399.5400 210.2200 400.8200 ;
      RECT 0.6250 399.1200 209.5950 399.5400 ;
      RECT 0.0000 397.8400 210.2200 399.1200 ;
      RECT 0.6250 397.4200 209.5950 397.8400 ;
      RECT 0.0000 396.1400 210.2200 397.4200 ;
      RECT 0.6250 395.7200 209.5950 396.1400 ;
      RECT 0.0000 394.4400 210.2200 395.7200 ;
      RECT 0.6250 394.0200 209.5950 394.4400 ;
      RECT 0.0000 392.7400 210.2200 394.0200 ;
      RECT 0.6250 392.3200 209.5950 392.7400 ;
      RECT 0.0000 390.7000 210.2200 392.3200 ;
      RECT 0.6250 390.2800 209.5950 390.7000 ;
      RECT 0.0000 389.0000 210.2200 390.2800 ;
      RECT 0.6250 388.5800 209.5950 389.0000 ;
      RECT 0.0000 387.3000 210.2200 388.5800 ;
      RECT 0.6250 386.8800 209.5950 387.3000 ;
      RECT 0.0000 385.6000 210.2200 386.8800 ;
      RECT 0.6250 385.1800 209.5950 385.6000 ;
      RECT 0.0000 383.9000 210.2200 385.1800 ;
      RECT 0.6250 383.4800 209.5950 383.9000 ;
      RECT 0.0000 382.2000 210.2200 383.4800 ;
      RECT 0.6250 381.7800 209.5950 382.2000 ;
      RECT 0.0000 380.5000 210.2200 381.7800 ;
      RECT 0.6250 380.0800 209.5950 380.5000 ;
      RECT 0.0000 375.0600 210.2200 380.0800 ;
      RECT 0.6250 374.6400 209.5950 375.0600 ;
      RECT 0.0000 373.3600 210.2200 374.6400 ;
      RECT 0.6250 372.9400 209.5950 373.3600 ;
      RECT 0.0000 372.0000 210.2200 372.9400 ;
      RECT 0.6250 371.5800 209.5950 372.0000 ;
      RECT 0.0000 370.6400 210.2200 371.5800 ;
      RECT 0.6250 370.2200 209.5950 370.6400 ;
      RECT 0.0000 368.9400 210.2200 370.2200 ;
      RECT 0.6250 368.5200 209.5950 368.9400 ;
      RECT 0.0000 367.5800 210.2200 368.5200 ;
      RECT 0.6250 367.1600 209.5950 367.5800 ;
      RECT 0.0000 366.2200 210.2200 367.1600 ;
      RECT 0.6250 365.8000 209.5950 366.2200 ;
      RECT 0.0000 364.5200 210.2200 365.8000 ;
      RECT 0.6250 364.1000 209.5950 364.5200 ;
      RECT 0.0000 363.1600 210.2200 364.1000 ;
      RECT 0.6250 362.7400 209.5950 363.1600 ;
      RECT 0.0000 361.8000 210.2200 362.7400 ;
      RECT 0.6250 361.3800 209.5950 361.8000 ;
      RECT 0.0000 360.1000 210.2200 361.3800 ;
      RECT 0.6250 359.6800 209.5950 360.1000 ;
      RECT 0.0000 358.7400 210.2200 359.6800 ;
      RECT 0.6250 358.3200 209.5950 358.7400 ;
      RECT 0.0000 357.3800 210.2200 358.3200 ;
      RECT 0.6250 356.9600 209.5950 357.3800 ;
      RECT 0.0000 355.6800 210.2200 356.9600 ;
      RECT 0.6250 355.2600 209.5950 355.6800 ;
      RECT 0.0000 354.3200 210.2200 355.2600 ;
      RECT 0.6250 353.9000 209.5950 354.3200 ;
      RECT 0.0000 352.9600 210.2200 353.9000 ;
      RECT 0.6250 352.5400 209.5950 352.9600 ;
      RECT 0.0000 351.2600 210.2200 352.5400 ;
      RECT 0.6250 350.8400 209.5950 351.2600 ;
      RECT 0.0000 349.9000 210.2200 350.8400 ;
      RECT 0.6250 349.4800 209.5950 349.9000 ;
      RECT 0.0000 348.5400 210.2200 349.4800 ;
      RECT 0.6250 348.1200 209.5950 348.5400 ;
      RECT 0.0000 346.8400 210.2200 348.1200 ;
      RECT 0.6250 346.4200 209.5950 346.8400 ;
      RECT 0.0000 345.4800 210.2200 346.4200 ;
      RECT 0.6250 345.0600 209.5950 345.4800 ;
      RECT 0.0000 344.1200 210.2200 345.0600 ;
      RECT 0.6250 343.7000 209.5950 344.1200 ;
      RECT 0.0000 342.4200 210.2200 343.7000 ;
      RECT 0.6250 342.0000 209.5950 342.4200 ;
      RECT 0.0000 341.0600 210.2200 342.0000 ;
      RECT 0.6250 340.6400 209.5950 341.0600 ;
      RECT 0.0000 339.7000 210.2200 340.6400 ;
      RECT 0.6250 339.2800 209.5950 339.7000 ;
      RECT 0.0000 338.0000 210.2200 339.2800 ;
      RECT 0.6250 337.5800 209.5950 338.0000 ;
      RECT 0.0000 336.6400 210.2200 337.5800 ;
      RECT 0.6250 336.2200 209.5950 336.6400 ;
      RECT 0.0000 335.2800 210.2200 336.2200 ;
      RECT 0.6250 334.8600 209.5950 335.2800 ;
      RECT 0.0000 333.5800 210.2200 334.8600 ;
      RECT 0.6250 333.1600 209.5950 333.5800 ;
      RECT 0.0000 332.2200 210.2200 333.1600 ;
      RECT 0.6250 331.8000 209.5950 332.2200 ;
      RECT 0.0000 330.8600 210.2200 331.8000 ;
      RECT 0.6250 330.4400 209.5950 330.8600 ;
      RECT 0.0000 329.1600 210.2200 330.4400 ;
      RECT 0.6250 328.7400 209.5950 329.1600 ;
      RECT 0.0000 327.8000 210.2200 328.7400 ;
      RECT 0.6250 327.3800 209.5950 327.8000 ;
      RECT 0.0000 326.4400 210.2200 327.3800 ;
      RECT 0.6250 326.0200 209.5950 326.4400 ;
      RECT 0.0000 324.7400 210.2200 326.0200 ;
      RECT 0.6250 324.3200 209.5950 324.7400 ;
      RECT 0.0000 323.3800 210.2200 324.3200 ;
      RECT 0.6250 322.9600 209.5950 323.3800 ;
      RECT 0.0000 322.0200 210.2200 322.9600 ;
      RECT 0.6250 321.6000 209.5950 322.0200 ;
      RECT 0.0000 320.3200 210.2200 321.6000 ;
      RECT 0.6250 319.9000 209.5950 320.3200 ;
      RECT 0.0000 318.9600 210.2200 319.9000 ;
      RECT 0.6250 318.5400 209.5950 318.9600 ;
      RECT 0.0000 317.6000 210.2200 318.5400 ;
      RECT 0.6250 317.1800 209.5950 317.6000 ;
      RECT 0.0000 315.9000 210.2200 317.1800 ;
      RECT 0.6250 315.4800 209.5950 315.9000 ;
      RECT 0.0000 314.5400 210.2200 315.4800 ;
      RECT 0.6250 314.1200 209.5950 314.5400 ;
      RECT 0.0000 313.1800 210.2200 314.1200 ;
      RECT 0.6250 312.7600 209.5950 313.1800 ;
      RECT 0.0000 311.4800 210.2200 312.7600 ;
      RECT 0.6250 311.0600 209.5950 311.4800 ;
      RECT 0.0000 310.1200 210.2200 311.0600 ;
      RECT 0.6250 309.7000 209.5950 310.1200 ;
      RECT 0.0000 308.7600 210.2200 309.7000 ;
      RECT 0.6250 308.3400 209.5950 308.7600 ;
      RECT 0.0000 307.0600 210.2200 308.3400 ;
      RECT 0.6250 306.6400 209.5950 307.0600 ;
      RECT 0.0000 305.7000 210.2200 306.6400 ;
      RECT 0.6250 305.2800 209.5950 305.7000 ;
      RECT 0.0000 304.3400 210.2200 305.2800 ;
      RECT 0.6250 303.9200 209.5950 304.3400 ;
      RECT 0.0000 302.9800 210.2200 303.9200 ;
      RECT 0.6250 302.5600 209.5950 302.9800 ;
      RECT 0.0000 301.2800 210.2200 302.5600 ;
      RECT 0.6250 300.8600 209.5950 301.2800 ;
      RECT 0.0000 299.9200 210.2200 300.8600 ;
      RECT 0.6250 299.5000 209.5950 299.9200 ;
      RECT 0.0000 298.5600 210.2200 299.5000 ;
      RECT 0.6250 298.1400 209.5950 298.5600 ;
      RECT 0.0000 296.8600 210.2200 298.1400 ;
      RECT 0.6250 296.4400 209.5950 296.8600 ;
      RECT 0.0000 295.5000 210.2200 296.4400 ;
      RECT 0.6250 295.0800 209.5950 295.5000 ;
      RECT 0.0000 294.1400 210.2200 295.0800 ;
      RECT 0.6250 293.7200 209.5950 294.1400 ;
      RECT 0.0000 292.4400 210.2200 293.7200 ;
      RECT 0.6250 292.0200 209.5950 292.4400 ;
      RECT 0.0000 291.0800 210.2200 292.0200 ;
      RECT 0.6250 290.6600 209.5950 291.0800 ;
      RECT 0.0000 289.7200 210.2200 290.6600 ;
      RECT 0.6250 289.3000 209.5950 289.7200 ;
      RECT 0.0000 288.0200 210.2200 289.3000 ;
      RECT 0.6250 287.6000 209.5950 288.0200 ;
      RECT 0.0000 286.6600 210.2200 287.6000 ;
      RECT 0.6250 286.2400 209.5950 286.6600 ;
      RECT 0.0000 285.3000 210.2200 286.2400 ;
      RECT 0.6250 284.8800 209.5950 285.3000 ;
      RECT 0.0000 283.6000 210.2200 284.8800 ;
      RECT 0.6250 283.1800 209.5950 283.6000 ;
      RECT 0.0000 282.2400 210.2200 283.1800 ;
      RECT 0.6250 281.8200 209.5950 282.2400 ;
      RECT 0.0000 280.8800 210.2200 281.8200 ;
      RECT 0.6250 280.4600 209.5950 280.8800 ;
      RECT 0.0000 279.1800 210.2200 280.4600 ;
      RECT 0.6250 278.7600 209.5950 279.1800 ;
      RECT 0.0000 277.8200 210.2200 278.7600 ;
      RECT 0.6250 277.4000 209.5950 277.8200 ;
      RECT 0.0000 276.4600 210.2200 277.4000 ;
      RECT 0.6250 276.0400 209.5950 276.4600 ;
      RECT 0.0000 274.7600 210.2200 276.0400 ;
      RECT 0.6250 274.3400 209.5950 274.7600 ;
      RECT 0.0000 273.4000 210.2200 274.3400 ;
      RECT 0.6250 272.9800 209.5950 273.4000 ;
      RECT 0.0000 272.0400 210.2200 272.9800 ;
      RECT 0.6250 271.6200 209.5950 272.0400 ;
      RECT 0.0000 270.3400 210.2200 271.6200 ;
      RECT 0.6250 269.9200 209.5950 270.3400 ;
      RECT 0.0000 268.9800 210.2200 269.9200 ;
      RECT 0.6250 268.5600 209.5950 268.9800 ;
      RECT 0.0000 267.6200 210.2200 268.5600 ;
      RECT 0.6250 267.2000 209.5950 267.6200 ;
      RECT 0.0000 265.9200 210.2200 267.2000 ;
      RECT 0.6250 265.5000 209.5950 265.9200 ;
      RECT 0.0000 264.5600 210.2200 265.5000 ;
      RECT 0.6250 264.1400 209.5950 264.5600 ;
      RECT 0.0000 263.2000 210.2200 264.1400 ;
      RECT 0.6250 262.7800 209.5950 263.2000 ;
      RECT 0.0000 261.5000 210.2200 262.7800 ;
      RECT 0.6250 261.0800 209.5950 261.5000 ;
      RECT 0.0000 260.1400 210.2200 261.0800 ;
      RECT 0.6250 259.7200 209.5950 260.1400 ;
      RECT 0.0000 258.7800 210.2200 259.7200 ;
      RECT 0.6250 258.3600 209.5950 258.7800 ;
      RECT 0.0000 257.0800 210.2200 258.3600 ;
      RECT 0.6250 256.6600 209.5950 257.0800 ;
      RECT 0.0000 255.7200 210.2200 256.6600 ;
      RECT 0.6250 255.3000 209.5950 255.7200 ;
      RECT 0.0000 254.3600 210.2200 255.3000 ;
      RECT 0.6250 253.9400 209.5950 254.3600 ;
      RECT 0.0000 252.6600 210.2200 253.9400 ;
      RECT 0.6250 252.2400 209.5950 252.6600 ;
      RECT 0.0000 251.3000 210.2200 252.2400 ;
      RECT 0.6250 250.8800 209.5950 251.3000 ;
      RECT 0.0000 249.9400 210.2200 250.8800 ;
      RECT 0.6250 249.5200 209.5950 249.9400 ;
      RECT 0.0000 248.2400 210.2200 249.5200 ;
      RECT 0.6250 247.8200 209.5950 248.2400 ;
      RECT 0.0000 246.8800 210.2200 247.8200 ;
      RECT 0.6250 246.4600 209.5950 246.8800 ;
      RECT 0.0000 245.5200 210.2200 246.4600 ;
      RECT 0.6250 245.1000 209.5950 245.5200 ;
      RECT 0.0000 243.8200 210.2200 245.1000 ;
      RECT 0.6250 243.4000 209.5950 243.8200 ;
      RECT 0.0000 242.4600 210.2200 243.4000 ;
      RECT 0.6250 242.0400 209.5950 242.4600 ;
      RECT 0.0000 241.1000 210.2200 242.0400 ;
      RECT 0.6250 240.6800 209.5950 241.1000 ;
      RECT 0.0000 239.4000 210.2200 240.6800 ;
      RECT 0.6250 238.9800 209.5950 239.4000 ;
      RECT 0.0000 238.0400 210.2200 238.9800 ;
      RECT 0.6250 237.6200 209.5950 238.0400 ;
      RECT 0.0000 236.6800 210.2200 237.6200 ;
      RECT 0.6250 236.2600 209.5950 236.6800 ;
      RECT 0.0000 235.3200 210.2200 236.2600 ;
      RECT 0.6250 234.9000 209.5950 235.3200 ;
      RECT 0.0000 209.8200 210.2200 234.9000 ;
      RECT 0.6250 209.4000 209.5950 209.8200 ;
      RECT 0.0000 208.1200 210.2200 209.4000 ;
      RECT 0.6250 207.7000 209.5950 208.1200 ;
      RECT 0.0000 206.4200 210.2200 207.7000 ;
      RECT 0.6250 206.0000 209.5950 206.4200 ;
      RECT 0.0000 204.7200 210.2200 206.0000 ;
      RECT 0.6250 204.3000 209.5950 204.7200 ;
      RECT 0.0000 203.0200 210.2200 204.3000 ;
      RECT 0.6250 202.6000 209.5950 203.0200 ;
      RECT 0.0000 201.3200 210.2200 202.6000 ;
      RECT 0.6250 200.9000 209.5950 201.3200 ;
      RECT 0.0000 199.2800 210.2200 200.9000 ;
      RECT 0.6250 198.8600 209.5950 199.2800 ;
      RECT 0.0000 197.5800 210.2200 198.8600 ;
      RECT 0.6250 197.1600 209.5950 197.5800 ;
      RECT 0.0000 195.8800 210.2200 197.1600 ;
      RECT 0.6250 195.4600 209.5950 195.8800 ;
      RECT 0.0000 194.1800 210.2200 195.4600 ;
      RECT 0.6250 193.7600 209.5950 194.1800 ;
      RECT 0.0000 192.4800 210.2200 193.7600 ;
      RECT 0.6250 192.0600 209.5950 192.4800 ;
      RECT 0.0000 190.4400 210.2200 192.0600 ;
      RECT 0.6250 190.0200 209.5950 190.4400 ;
      RECT 0.0000 188.7400 210.2200 190.0200 ;
      RECT 0.6250 188.3200 209.5950 188.7400 ;
      RECT 0.0000 187.0400 210.2200 188.3200 ;
      RECT 0.6250 186.6200 209.5950 187.0400 ;
      RECT 0.0000 185.3400 210.2200 186.6200 ;
      RECT 0.6250 184.9200 209.5950 185.3400 ;
      RECT 0.0000 183.6400 210.2200 184.9200 ;
      RECT 0.6250 183.2200 209.5950 183.6400 ;
      RECT 0.0000 181.6000 210.2200 183.2200 ;
      RECT 0.6250 181.1800 209.5950 181.6000 ;
      RECT 0.0000 179.9000 210.2200 181.1800 ;
      RECT 0.6250 179.4800 209.5950 179.9000 ;
      RECT 0.0000 178.2000 210.2200 179.4800 ;
      RECT 0.6250 177.7800 209.5950 178.2000 ;
      RECT 0.0000 176.5000 210.2200 177.7800 ;
      RECT 0.6250 176.0800 209.5950 176.5000 ;
      RECT 0.0000 174.8000 210.2200 176.0800 ;
      RECT 0.6250 174.3800 209.5950 174.8000 ;
      RECT 0.0000 172.7600 210.2200 174.3800 ;
      RECT 0.6250 172.3400 209.5950 172.7600 ;
      RECT 0.0000 171.0600 210.2200 172.3400 ;
      RECT 0.6250 170.6400 209.5950 171.0600 ;
      RECT 0.0000 169.3600 210.2200 170.6400 ;
      RECT 0.6250 168.9400 209.5950 169.3600 ;
      RECT 0.0000 167.6600 210.2200 168.9400 ;
      RECT 0.6250 167.2400 209.5950 167.6600 ;
      RECT 0.0000 165.9600 210.2200 167.2400 ;
      RECT 0.6250 165.5400 209.5950 165.9600 ;
      RECT 0.0000 163.9200 210.2200 165.5400 ;
      RECT 0.6250 163.5000 209.5950 163.9200 ;
      RECT 0.0000 162.2200 210.2200 163.5000 ;
      RECT 0.6250 161.8000 209.5950 162.2200 ;
      RECT 0.0000 160.5200 210.2200 161.8000 ;
      RECT 0.6250 160.1000 209.5950 160.5200 ;
      RECT 0.0000 158.8200 210.2200 160.1000 ;
      RECT 0.6250 158.4000 209.5950 158.8200 ;
      RECT 0.0000 157.1200 210.2200 158.4000 ;
      RECT 0.6250 156.7000 209.5950 157.1200 ;
      RECT 0.0000 155.4200 210.2200 156.7000 ;
      RECT 0.6250 155.0000 209.5950 155.4200 ;
      RECT 0.0000 149.9800 210.2200 155.0000 ;
      RECT 0.6250 149.5600 209.5950 149.9800 ;
      RECT 0.0000 148.2800 210.2200 149.5600 ;
      RECT 0.6250 147.8600 209.5950 148.2800 ;
      RECT 0.0000 146.9200 210.2200 147.8600 ;
      RECT 0.6250 146.5000 209.5950 146.9200 ;
      RECT 0.0000 145.5600 210.2200 146.5000 ;
      RECT 0.6250 145.1400 209.5950 145.5600 ;
      RECT 0.0000 143.8600 210.2200 145.1400 ;
      RECT 0.6250 143.4400 209.5950 143.8600 ;
      RECT 0.0000 142.5000 210.2200 143.4400 ;
      RECT 0.6250 142.0800 209.5950 142.5000 ;
      RECT 0.0000 141.1400 210.2200 142.0800 ;
      RECT 0.6250 140.7200 209.5950 141.1400 ;
      RECT 0.0000 139.4400 210.2200 140.7200 ;
      RECT 0.6250 139.0200 209.5950 139.4400 ;
      RECT 0.0000 138.0800 210.2200 139.0200 ;
      RECT 0.6250 137.6600 209.5950 138.0800 ;
      RECT 0.0000 136.7200 210.2200 137.6600 ;
      RECT 0.6250 136.3000 209.5950 136.7200 ;
      RECT 0.0000 135.0200 210.2200 136.3000 ;
      RECT 0.6250 134.6000 209.5950 135.0200 ;
      RECT 0.0000 133.6600 210.2200 134.6000 ;
      RECT 0.6250 133.2400 209.5950 133.6600 ;
      RECT 0.0000 132.3000 210.2200 133.2400 ;
      RECT 0.6250 131.8800 209.5950 132.3000 ;
      RECT 0.0000 130.6000 210.2200 131.8800 ;
      RECT 0.6250 130.1800 209.5950 130.6000 ;
      RECT 0.0000 129.2400 210.2200 130.1800 ;
      RECT 0.6250 128.8200 209.5950 129.2400 ;
      RECT 0.0000 127.8800 210.2200 128.8200 ;
      RECT 0.6250 127.4600 209.5950 127.8800 ;
      RECT 0.0000 126.1800 210.2200 127.4600 ;
      RECT 0.6250 125.7600 209.5950 126.1800 ;
      RECT 0.0000 124.8200 210.2200 125.7600 ;
      RECT 0.6250 124.4000 209.5950 124.8200 ;
      RECT 0.0000 123.4600 210.2200 124.4000 ;
      RECT 0.6250 123.0400 209.5950 123.4600 ;
      RECT 0.0000 121.7600 210.2200 123.0400 ;
      RECT 0.6250 121.3400 209.5950 121.7600 ;
      RECT 0.0000 120.4000 210.2200 121.3400 ;
      RECT 0.6250 119.9800 209.5950 120.4000 ;
      RECT 0.0000 119.0400 210.2200 119.9800 ;
      RECT 0.6250 118.6200 209.5950 119.0400 ;
      RECT 0.0000 117.3400 210.2200 118.6200 ;
      RECT 0.6250 116.9200 209.5950 117.3400 ;
      RECT 0.0000 115.9800 210.2200 116.9200 ;
      RECT 0.6250 115.5600 209.5950 115.9800 ;
      RECT 0.0000 114.6200 210.2200 115.5600 ;
      RECT 0.6250 114.2000 209.5950 114.6200 ;
      RECT 0.0000 112.9200 210.2200 114.2000 ;
      RECT 0.6250 112.5000 209.5950 112.9200 ;
      RECT 0.0000 111.5600 210.2200 112.5000 ;
      RECT 0.6250 111.1400 209.5950 111.5600 ;
      RECT 0.0000 110.2000 210.2200 111.1400 ;
      RECT 0.6250 109.7800 209.5950 110.2000 ;
      RECT 0.0000 108.5000 210.2200 109.7800 ;
      RECT 0.6250 108.0800 209.5950 108.5000 ;
      RECT 0.0000 107.1400 210.2200 108.0800 ;
      RECT 0.6250 106.7200 209.5950 107.1400 ;
      RECT 0.0000 105.7800 210.2200 106.7200 ;
      RECT 0.6250 105.3600 209.5950 105.7800 ;
      RECT 0.0000 104.0800 210.2200 105.3600 ;
      RECT 0.6250 103.6600 209.5950 104.0800 ;
      RECT 0.0000 102.7200 210.2200 103.6600 ;
      RECT 0.6250 102.3000 209.5950 102.7200 ;
      RECT 0.0000 101.3600 210.2200 102.3000 ;
      RECT 0.6250 100.9400 209.5950 101.3600 ;
      RECT 0.0000 99.6600 210.2200 100.9400 ;
      RECT 0.6250 99.2400 209.5950 99.6600 ;
      RECT 0.0000 98.3000 210.2200 99.2400 ;
      RECT 0.6250 97.8800 209.5950 98.3000 ;
      RECT 0.0000 96.9400 210.2200 97.8800 ;
      RECT 0.6250 96.5200 209.5950 96.9400 ;
      RECT 0.0000 95.2400 210.2200 96.5200 ;
      RECT 0.6250 94.8200 209.5950 95.2400 ;
      RECT 0.0000 93.8800 210.2200 94.8200 ;
      RECT 0.6250 93.4600 209.5950 93.8800 ;
      RECT 0.0000 92.5200 210.2200 93.4600 ;
      RECT 0.6250 92.1000 209.5950 92.5200 ;
      RECT 0.0000 90.8200 210.2200 92.1000 ;
      RECT 0.6250 90.4000 209.5950 90.8200 ;
      RECT 0.0000 89.4600 210.2200 90.4000 ;
      RECT 0.6250 89.0400 209.5950 89.4600 ;
      RECT 0.0000 88.1000 210.2200 89.0400 ;
      RECT 0.6250 87.6800 209.5950 88.1000 ;
      RECT 0.0000 86.4000 210.2200 87.6800 ;
      RECT 0.6250 85.9800 209.5950 86.4000 ;
      RECT 0.0000 85.0400 210.2200 85.9800 ;
      RECT 0.6250 84.6200 209.5950 85.0400 ;
      RECT 0.0000 83.6800 210.2200 84.6200 ;
      RECT 0.6250 83.2600 209.5950 83.6800 ;
      RECT 0.0000 81.9800 210.2200 83.2600 ;
      RECT 0.6250 81.5600 209.5950 81.9800 ;
      RECT 0.0000 80.6200 210.2200 81.5600 ;
      RECT 0.6250 80.2000 209.5950 80.6200 ;
      RECT 0.0000 79.2600 210.2200 80.2000 ;
      RECT 0.6250 78.8400 209.5950 79.2600 ;
      RECT 0.0000 77.9000 210.2200 78.8400 ;
      RECT 0.6250 77.4800 209.5950 77.9000 ;
      RECT 0.0000 76.2000 210.2200 77.4800 ;
      RECT 0.6250 75.7800 209.5950 76.2000 ;
      RECT 0.0000 74.8400 210.2200 75.7800 ;
      RECT 0.6250 74.4200 209.5950 74.8400 ;
      RECT 0.0000 73.4800 210.2200 74.4200 ;
      RECT 0.6250 73.0600 209.5950 73.4800 ;
      RECT 0.0000 71.7800 210.2200 73.0600 ;
      RECT 0.6250 71.3600 209.5950 71.7800 ;
      RECT 0.0000 70.4200 210.2200 71.3600 ;
      RECT 0.6250 70.0000 209.5950 70.4200 ;
      RECT 0.0000 69.0600 210.2200 70.0000 ;
      RECT 0.6250 68.6400 209.5950 69.0600 ;
      RECT 0.0000 67.3600 210.2200 68.6400 ;
      RECT 0.6250 66.9400 209.5950 67.3600 ;
      RECT 0.0000 66.0000 210.2200 66.9400 ;
      RECT 0.6250 65.5800 209.5950 66.0000 ;
      RECT 0.0000 64.6400 210.2200 65.5800 ;
      RECT 0.6250 64.2200 209.5950 64.6400 ;
      RECT 0.0000 62.9400 210.2200 64.2200 ;
      RECT 0.6250 62.5200 209.5950 62.9400 ;
      RECT 0.0000 61.5800 210.2200 62.5200 ;
      RECT 0.6250 61.1600 209.5950 61.5800 ;
      RECT 0.0000 60.2200 210.2200 61.1600 ;
      RECT 0.6250 59.8000 209.5950 60.2200 ;
      RECT 0.0000 58.5200 210.2200 59.8000 ;
      RECT 0.6250 58.1000 209.5950 58.5200 ;
      RECT 0.0000 57.1600 210.2200 58.1000 ;
      RECT 0.6250 56.7400 209.5950 57.1600 ;
      RECT 0.0000 55.8000 210.2200 56.7400 ;
      RECT 0.6250 55.3800 209.5950 55.8000 ;
      RECT 0.0000 54.1000 210.2200 55.3800 ;
      RECT 0.6250 53.6800 209.5950 54.1000 ;
      RECT 0.0000 52.7400 210.2200 53.6800 ;
      RECT 0.6250 52.3200 209.5950 52.7400 ;
      RECT 0.0000 51.3800 210.2200 52.3200 ;
      RECT 0.6250 50.9600 209.5950 51.3800 ;
      RECT 0.0000 49.6800 210.2200 50.9600 ;
      RECT 0.6250 49.2600 209.5950 49.6800 ;
      RECT 0.0000 48.3200 210.2200 49.2600 ;
      RECT 0.6250 47.9000 209.5950 48.3200 ;
      RECT 0.0000 46.9600 210.2200 47.9000 ;
      RECT 0.6250 46.5400 209.5950 46.9600 ;
      RECT 0.0000 45.2600 210.2200 46.5400 ;
      RECT 0.6250 44.8400 209.5950 45.2600 ;
      RECT 0.0000 43.9000 210.2200 44.8400 ;
      RECT 0.6250 43.4800 209.5950 43.9000 ;
      RECT 0.0000 42.5400 210.2200 43.4800 ;
      RECT 0.6250 42.1200 209.5950 42.5400 ;
      RECT 0.0000 40.8400 210.2200 42.1200 ;
      RECT 0.6250 40.4200 209.5950 40.8400 ;
      RECT 0.0000 39.4800 210.2200 40.4200 ;
      RECT 0.6250 39.0600 209.5950 39.4800 ;
      RECT 0.0000 38.1200 210.2200 39.0600 ;
      RECT 0.6250 37.7000 209.5950 38.1200 ;
      RECT 0.0000 36.4200 210.2200 37.7000 ;
      RECT 0.6250 36.0000 209.5950 36.4200 ;
      RECT 0.0000 35.0600 210.2200 36.0000 ;
      RECT 0.6250 34.6400 209.5950 35.0600 ;
      RECT 0.0000 33.7000 210.2200 34.6400 ;
      RECT 0.6250 33.2800 209.5950 33.7000 ;
      RECT 0.0000 32.0000 210.2200 33.2800 ;
      RECT 0.6250 31.5800 209.5950 32.0000 ;
      RECT 0.0000 30.6400 210.2200 31.5800 ;
      RECT 0.6250 30.2200 209.5950 30.6400 ;
      RECT 0.0000 29.2800 210.2200 30.2200 ;
      RECT 0.6250 28.8600 209.5950 29.2800 ;
      RECT 0.0000 27.5800 210.2200 28.8600 ;
      RECT 0.6250 27.1600 209.5950 27.5800 ;
      RECT 0.0000 26.2200 210.2200 27.1600 ;
      RECT 0.6250 25.8000 209.5950 26.2200 ;
      RECT 0.0000 24.8600 210.2200 25.8000 ;
      RECT 0.6250 24.4400 209.5950 24.8600 ;
      RECT 0.0000 23.1600 210.2200 24.4400 ;
      RECT 0.6250 22.7400 209.5950 23.1600 ;
      RECT 0.0000 21.8000 210.2200 22.7400 ;
      RECT 0.6250 21.3800 209.5950 21.8000 ;
      RECT 0.0000 20.4400 210.2200 21.3800 ;
      RECT 0.6250 20.0200 209.5950 20.4400 ;
      RECT 0.0000 18.7400 210.2200 20.0200 ;
      RECT 0.6250 18.3200 209.5950 18.7400 ;
      RECT 0.0000 17.3800 210.2200 18.3200 ;
      RECT 0.6250 16.9600 209.5950 17.3800 ;
      RECT 0.0000 16.0200 210.2200 16.9600 ;
      RECT 0.6250 15.6000 209.5950 16.0200 ;
      RECT 0.0000 14.3200 210.2200 15.6000 ;
      RECT 0.6250 13.9000 209.5950 14.3200 ;
      RECT 0.0000 12.9600 210.2200 13.9000 ;
      RECT 0.6250 12.5400 209.5950 12.9600 ;
      RECT 0.0000 11.6000 210.2200 12.5400 ;
      RECT 0.6250 11.1800 209.5950 11.6000 ;
      RECT 0.0000 10.2400 210.2200 11.1800 ;
      RECT 0.6250 9.8200 209.5950 10.2400 ;
      RECT 0.0000 0.6250 210.2200 9.8200 ;
      RECT 200.0800 0.0000 210.2200 0.6250 ;
      RECT 197.3200 0.0000 199.6600 0.6250 ;
      RECT 195.0200 0.0000 196.9000 0.6250 ;
      RECT 192.7200 0.0000 194.6000 0.6250 ;
      RECT 190.4200 0.0000 192.3000 0.6250 ;
      RECT 188.1200 0.0000 190.0000 0.6250 ;
      RECT 185.8200 0.0000 187.7000 0.6250 ;
      RECT 183.5200 0.0000 185.4000 0.6250 ;
      RECT 181.2200 0.0000 183.1000 0.6250 ;
      RECT 178.9200 0.0000 180.8000 0.6250 ;
      RECT 176.1600 0.0000 178.5000 0.6250 ;
      RECT 173.8600 0.0000 175.7400 0.6250 ;
      RECT 171.5600 0.0000 173.4400 0.6250 ;
      RECT 169.2600 0.0000 171.1400 0.6250 ;
      RECT 166.9600 0.0000 168.8400 0.6250 ;
      RECT 164.6600 0.0000 166.5400 0.6250 ;
      RECT 162.3600 0.0000 164.2400 0.6250 ;
      RECT 160.0600 0.0000 161.9400 0.6250 ;
      RECT 157.7600 0.0000 159.6400 0.6250 ;
      RECT 155.4600 0.0000 157.3400 0.6250 ;
      RECT 0.0000 0.0000 155.0400 0.6250 ;
    LAYER met3 ;
      RECT 0.0000 442.2500 210.2200 444.7200 ;
      RECT 207.9600 439.6500 210.2200 442.2500 ;
      RECT 0.0000 439.6500 2.2600 442.2500 ;
      RECT 0.0000 439.2500 210.2200 439.6500 ;
      RECT 204.9600 436.6500 210.2200 439.2500 ;
      RECT 0.0000 436.6500 5.2600 439.2500 ;
      RECT 0.0000 434.7200 210.2200 436.6500 ;
      RECT 207.9600 433.6400 210.2200 434.7200 ;
      RECT 4.8600 433.6400 205.3600 434.7200 ;
      RECT 0.0000 433.6400 2.2600 434.7200 ;
      RECT 0.0000 432.0000 210.2200 433.6400 ;
      RECT 204.9600 430.9200 210.2200 432.0000 ;
      RECT 7.8600 430.9200 202.3600 432.0000 ;
      RECT 0.0000 430.9200 5.2600 432.0000 ;
      RECT 0.0000 429.2800 210.2200 430.9200 ;
      RECT 207.9600 428.2000 210.2200 429.2800 ;
      RECT 4.8600 428.2000 205.3600 429.2800 ;
      RECT 0.0000 428.2000 2.2600 429.2800 ;
      RECT 0.0000 426.5600 210.2200 428.2000 ;
      RECT 204.9600 425.4800 210.2200 426.5600 ;
      RECT 7.8600 425.4800 202.3600 426.5600 ;
      RECT 0.0000 425.4800 5.2600 426.5600 ;
      RECT 0.0000 423.8400 210.2200 425.4800 ;
      RECT 207.9600 422.7600 210.2200 423.8400 ;
      RECT 4.8600 422.7600 205.3600 423.8400 ;
      RECT 0.0000 422.7600 2.2600 423.8400 ;
      RECT 0.0000 421.1200 210.2200 422.7600 ;
      RECT 204.9600 420.0400 210.2200 421.1200 ;
      RECT 7.8600 420.0400 202.3600 421.1200 ;
      RECT 0.0000 420.0400 5.2600 421.1200 ;
      RECT 0.0000 418.4000 210.2200 420.0400 ;
      RECT 207.9600 417.3200 210.2200 418.4000 ;
      RECT 4.8600 417.3200 205.3600 418.4000 ;
      RECT 0.0000 417.3200 2.2600 418.4000 ;
      RECT 0.0000 415.6800 210.2200 417.3200 ;
      RECT 204.9600 414.6000 210.2200 415.6800 ;
      RECT 7.8600 414.6000 202.3600 415.6800 ;
      RECT 0.0000 414.6000 5.2600 415.6800 ;
      RECT 0.0000 412.9600 210.2200 414.6000 ;
      RECT 207.9600 411.8800 210.2200 412.9600 ;
      RECT 4.8600 411.8800 205.3600 412.9600 ;
      RECT 0.0000 411.8800 2.2600 412.9600 ;
      RECT 0.0000 410.2400 210.2200 411.8800 ;
      RECT 204.9600 409.1600 210.2200 410.2400 ;
      RECT 7.8600 409.1600 202.3600 410.2400 ;
      RECT 0.0000 409.1600 5.2600 410.2400 ;
      RECT 0.0000 407.5200 210.2200 409.1600 ;
      RECT 207.9600 406.4400 210.2200 407.5200 ;
      RECT 4.8600 406.4400 205.3600 407.5200 ;
      RECT 0.0000 406.4400 2.2600 407.5200 ;
      RECT 0.0000 404.8000 210.2200 406.4400 ;
      RECT 204.9600 403.7200 210.2200 404.8000 ;
      RECT 7.8600 403.7200 202.3600 404.8000 ;
      RECT 0.0000 403.7200 5.2600 404.8000 ;
      RECT 0.0000 402.0800 210.2200 403.7200 ;
      RECT 207.9600 401.0000 210.2200 402.0800 ;
      RECT 4.8600 401.0000 205.3600 402.0800 ;
      RECT 0.0000 401.0000 2.2600 402.0800 ;
      RECT 0.0000 399.3600 210.2200 401.0000 ;
      RECT 204.9600 398.2800 210.2200 399.3600 ;
      RECT 7.8600 398.2800 202.3600 399.3600 ;
      RECT 0.0000 398.2800 5.2600 399.3600 ;
      RECT 0.0000 396.6400 210.2200 398.2800 ;
      RECT 207.9600 395.5600 210.2200 396.6400 ;
      RECT 4.8600 395.5600 205.3600 396.6400 ;
      RECT 0.0000 395.5600 2.2600 396.6400 ;
      RECT 0.0000 393.9200 210.2200 395.5600 ;
      RECT 204.9600 392.8400 210.2200 393.9200 ;
      RECT 7.8600 392.8400 202.3600 393.9200 ;
      RECT 0.0000 392.8400 5.2600 393.9200 ;
      RECT 0.0000 391.2000 210.2200 392.8400 ;
      RECT 207.9600 390.1200 210.2200 391.2000 ;
      RECT 4.8600 390.1200 205.3600 391.2000 ;
      RECT 0.0000 390.1200 2.2600 391.2000 ;
      RECT 0.0000 388.4800 210.2200 390.1200 ;
      RECT 204.9600 387.4000 210.2200 388.4800 ;
      RECT 7.8600 387.4000 202.3600 388.4800 ;
      RECT 0.0000 387.4000 5.2600 388.4800 ;
      RECT 0.0000 385.7600 210.2200 387.4000 ;
      RECT 207.9600 384.6800 210.2200 385.7600 ;
      RECT 4.8600 384.6800 205.3600 385.7600 ;
      RECT 0.0000 384.6800 2.2600 385.7600 ;
      RECT 0.0000 383.0400 210.2200 384.6800 ;
      RECT 204.9600 381.9600 210.2200 383.0400 ;
      RECT 7.8600 381.9600 202.3600 383.0400 ;
      RECT 0.0000 381.9600 5.2600 383.0400 ;
      RECT 0.0000 380.3200 210.2200 381.9600 ;
      RECT 207.9600 379.2400 210.2200 380.3200 ;
      RECT 4.8600 379.2400 205.3600 380.3200 ;
      RECT 0.0000 379.2400 2.2600 380.3200 ;
      RECT 0.0000 377.6000 210.2200 379.2400 ;
      RECT 204.9600 376.5200 210.2200 377.6000 ;
      RECT 7.8600 376.5200 202.3600 377.6000 ;
      RECT 0.0000 376.5200 5.2600 377.6000 ;
      RECT 0.0000 374.8800 210.2200 376.5200 ;
      RECT 207.9600 373.8000 210.2200 374.8800 ;
      RECT 4.8600 373.8000 205.3600 374.8800 ;
      RECT 0.0000 373.8000 2.2600 374.8800 ;
      RECT 0.0000 372.1600 210.2200 373.8000 ;
      RECT 204.9600 371.0800 210.2200 372.1600 ;
      RECT 7.8600 371.0800 202.3600 372.1600 ;
      RECT 0.0000 371.0800 5.2600 372.1600 ;
      RECT 0.0000 369.4400 210.2200 371.0800 ;
      RECT 207.9600 368.3600 210.2200 369.4400 ;
      RECT 4.8600 368.3600 205.3600 369.4400 ;
      RECT 0.0000 368.3600 2.2600 369.4400 ;
      RECT 0.0000 366.7200 210.2200 368.3600 ;
      RECT 204.9600 365.6400 210.2200 366.7200 ;
      RECT 7.8600 365.6400 202.3600 366.7200 ;
      RECT 0.0000 365.6400 5.2600 366.7200 ;
      RECT 0.0000 364.0000 210.2200 365.6400 ;
      RECT 207.9600 362.9200 210.2200 364.0000 ;
      RECT 4.8600 362.9200 205.3600 364.0000 ;
      RECT 0.0000 362.9200 2.2600 364.0000 ;
      RECT 0.0000 361.2800 210.2200 362.9200 ;
      RECT 204.9600 360.2000 210.2200 361.2800 ;
      RECT 7.8600 360.2000 202.3600 361.2800 ;
      RECT 0.0000 360.2000 5.2600 361.2800 ;
      RECT 0.0000 358.5600 210.2200 360.2000 ;
      RECT 207.9600 357.4800 210.2200 358.5600 ;
      RECT 4.8600 357.4800 205.3600 358.5600 ;
      RECT 0.0000 357.4800 2.2600 358.5600 ;
      RECT 0.0000 355.8400 210.2200 357.4800 ;
      RECT 204.9600 354.7600 210.2200 355.8400 ;
      RECT 7.8600 354.7600 202.3600 355.8400 ;
      RECT 0.0000 354.7600 5.2600 355.8400 ;
      RECT 0.0000 353.1200 210.2200 354.7600 ;
      RECT 207.9600 352.0400 210.2200 353.1200 ;
      RECT 4.8600 352.0400 205.3600 353.1200 ;
      RECT 0.0000 352.0400 2.2600 353.1200 ;
      RECT 0.0000 350.4000 210.2200 352.0400 ;
      RECT 204.9600 349.3200 210.2200 350.4000 ;
      RECT 7.8600 349.3200 202.3600 350.4000 ;
      RECT 0.0000 349.3200 5.2600 350.4000 ;
      RECT 0.0000 347.6800 210.2200 349.3200 ;
      RECT 207.9600 346.6000 210.2200 347.6800 ;
      RECT 4.8600 346.6000 205.3600 347.6800 ;
      RECT 0.0000 346.6000 2.2600 347.6800 ;
      RECT 0.0000 344.9600 210.2200 346.6000 ;
      RECT 204.9600 343.8800 210.2200 344.9600 ;
      RECT 7.8600 343.8800 202.3600 344.9600 ;
      RECT 0.0000 343.8800 5.2600 344.9600 ;
      RECT 0.0000 342.2400 210.2200 343.8800 ;
      RECT 207.9600 341.1600 210.2200 342.2400 ;
      RECT 4.8600 341.1600 205.3600 342.2400 ;
      RECT 0.0000 341.1600 2.2600 342.2400 ;
      RECT 0.0000 339.5200 210.2200 341.1600 ;
      RECT 204.9600 338.4400 210.2200 339.5200 ;
      RECT 7.8600 338.4400 202.3600 339.5200 ;
      RECT 0.0000 338.4400 5.2600 339.5200 ;
      RECT 0.0000 336.8000 210.2200 338.4400 ;
      RECT 207.9600 335.7200 210.2200 336.8000 ;
      RECT 4.8600 335.7200 205.3600 336.8000 ;
      RECT 0.0000 335.7200 2.2600 336.8000 ;
      RECT 0.0000 334.0800 210.2200 335.7200 ;
      RECT 204.9600 333.0000 210.2200 334.0800 ;
      RECT 7.8600 333.0000 202.3600 334.0800 ;
      RECT 0.0000 333.0000 5.2600 334.0800 ;
      RECT 0.0000 331.3600 210.2200 333.0000 ;
      RECT 207.9600 330.2800 210.2200 331.3600 ;
      RECT 4.8600 330.2800 205.3600 331.3600 ;
      RECT 0.0000 330.2800 2.2600 331.3600 ;
      RECT 0.0000 328.6400 210.2200 330.2800 ;
      RECT 204.9600 327.5600 210.2200 328.6400 ;
      RECT 7.8600 327.5600 202.3600 328.6400 ;
      RECT 0.0000 327.5600 5.2600 328.6400 ;
      RECT 0.0000 325.9200 210.2200 327.5600 ;
      RECT 207.9600 324.8400 210.2200 325.9200 ;
      RECT 4.8600 324.8400 205.3600 325.9200 ;
      RECT 0.0000 324.8400 2.2600 325.9200 ;
      RECT 0.0000 323.2000 210.2200 324.8400 ;
      RECT 204.9600 322.1200 210.2200 323.2000 ;
      RECT 7.8600 322.1200 202.3600 323.2000 ;
      RECT 0.0000 322.1200 5.2600 323.2000 ;
      RECT 0.0000 320.4800 210.2200 322.1200 ;
      RECT 207.9600 319.4000 210.2200 320.4800 ;
      RECT 4.8600 319.4000 205.3600 320.4800 ;
      RECT 0.0000 319.4000 2.2600 320.4800 ;
      RECT 0.0000 317.7600 210.2200 319.4000 ;
      RECT 204.9600 316.6800 210.2200 317.7600 ;
      RECT 7.8600 316.6800 202.3600 317.7600 ;
      RECT 0.0000 316.6800 5.2600 317.7600 ;
      RECT 0.0000 315.0400 210.2200 316.6800 ;
      RECT 207.9600 313.9600 210.2200 315.0400 ;
      RECT 4.8600 313.9600 205.3600 315.0400 ;
      RECT 0.0000 313.9600 2.2600 315.0400 ;
      RECT 0.0000 312.3200 210.2200 313.9600 ;
      RECT 204.9600 311.2400 210.2200 312.3200 ;
      RECT 7.8600 311.2400 202.3600 312.3200 ;
      RECT 0.0000 311.2400 5.2600 312.3200 ;
      RECT 0.0000 309.6000 210.2200 311.2400 ;
      RECT 207.9600 308.5200 210.2200 309.6000 ;
      RECT 4.8600 308.5200 205.3600 309.6000 ;
      RECT 0.0000 308.5200 2.2600 309.6000 ;
      RECT 0.0000 306.8800 210.2200 308.5200 ;
      RECT 204.9600 305.8000 210.2200 306.8800 ;
      RECT 7.8600 305.8000 202.3600 306.8800 ;
      RECT 0.0000 305.8000 5.2600 306.8800 ;
      RECT 0.0000 304.1600 210.2200 305.8000 ;
      RECT 207.9600 303.0800 210.2200 304.1600 ;
      RECT 4.8600 303.0800 205.3600 304.1600 ;
      RECT 0.0000 303.0800 2.2600 304.1600 ;
      RECT 0.0000 301.4400 210.2200 303.0800 ;
      RECT 204.9600 300.3600 210.2200 301.4400 ;
      RECT 7.8600 300.3600 202.3600 301.4400 ;
      RECT 0.0000 300.3600 5.2600 301.4400 ;
      RECT 0.0000 298.7200 210.2200 300.3600 ;
      RECT 207.9600 297.6400 210.2200 298.7200 ;
      RECT 4.8600 297.6400 205.3600 298.7200 ;
      RECT 0.0000 297.6400 2.2600 298.7200 ;
      RECT 0.0000 296.0000 210.2200 297.6400 ;
      RECT 204.9600 294.9200 210.2200 296.0000 ;
      RECT 7.8600 294.9200 202.3600 296.0000 ;
      RECT 0.0000 294.9200 5.2600 296.0000 ;
      RECT 0.0000 293.2800 210.2200 294.9200 ;
      RECT 207.9600 292.2000 210.2200 293.2800 ;
      RECT 4.8600 292.2000 205.3600 293.2800 ;
      RECT 0.0000 292.2000 2.2600 293.2800 ;
      RECT 0.0000 290.5600 210.2200 292.2000 ;
      RECT 204.9600 289.4800 210.2200 290.5600 ;
      RECT 7.8600 289.4800 202.3600 290.5600 ;
      RECT 0.0000 289.4800 5.2600 290.5600 ;
      RECT 0.0000 287.8400 210.2200 289.4800 ;
      RECT 207.9600 286.7600 210.2200 287.8400 ;
      RECT 4.8600 286.7600 205.3600 287.8400 ;
      RECT 0.0000 286.7600 2.2600 287.8400 ;
      RECT 0.0000 285.1200 210.2200 286.7600 ;
      RECT 204.9600 284.0400 210.2200 285.1200 ;
      RECT 7.8600 284.0400 202.3600 285.1200 ;
      RECT 0.0000 284.0400 5.2600 285.1200 ;
      RECT 0.0000 282.4000 210.2200 284.0400 ;
      RECT 207.9600 281.3200 210.2200 282.4000 ;
      RECT 4.8600 281.3200 205.3600 282.4000 ;
      RECT 0.0000 281.3200 2.2600 282.4000 ;
      RECT 0.0000 279.6800 210.2200 281.3200 ;
      RECT 204.9600 278.6000 210.2200 279.6800 ;
      RECT 7.8600 278.6000 202.3600 279.6800 ;
      RECT 0.0000 278.6000 5.2600 279.6800 ;
      RECT 0.0000 276.9600 210.2200 278.6000 ;
      RECT 207.9600 275.8800 210.2200 276.9600 ;
      RECT 4.8600 275.8800 205.3600 276.9600 ;
      RECT 0.0000 275.8800 2.2600 276.9600 ;
      RECT 0.0000 274.2400 210.2200 275.8800 ;
      RECT 204.9600 273.1600 210.2200 274.2400 ;
      RECT 7.8600 273.1600 202.3600 274.2400 ;
      RECT 0.0000 273.1600 5.2600 274.2400 ;
      RECT 0.0000 271.5200 210.2200 273.1600 ;
      RECT 207.9600 270.4400 210.2200 271.5200 ;
      RECT 4.8600 270.4400 205.3600 271.5200 ;
      RECT 0.0000 270.4400 2.2600 271.5200 ;
      RECT 0.0000 268.8000 210.2200 270.4400 ;
      RECT 204.9600 267.7200 210.2200 268.8000 ;
      RECT 7.8600 267.7200 202.3600 268.8000 ;
      RECT 0.0000 267.7200 5.2600 268.8000 ;
      RECT 0.0000 266.0800 210.2200 267.7200 ;
      RECT 207.9600 265.0000 210.2200 266.0800 ;
      RECT 4.8600 265.0000 205.3600 266.0800 ;
      RECT 0.0000 265.0000 2.2600 266.0800 ;
      RECT 0.0000 263.3600 210.2200 265.0000 ;
      RECT 204.9600 262.2800 210.2200 263.3600 ;
      RECT 7.8600 262.2800 202.3600 263.3600 ;
      RECT 0.0000 262.2800 5.2600 263.3600 ;
      RECT 0.0000 260.6400 210.2200 262.2800 ;
      RECT 207.9600 259.5600 210.2200 260.6400 ;
      RECT 4.8600 259.5600 205.3600 260.6400 ;
      RECT 0.0000 259.5600 2.2600 260.6400 ;
      RECT 0.0000 257.9200 210.2200 259.5600 ;
      RECT 204.9600 256.8400 210.2200 257.9200 ;
      RECT 7.8600 256.8400 202.3600 257.9200 ;
      RECT 0.0000 256.8400 5.2600 257.9200 ;
      RECT 0.0000 255.2000 210.2200 256.8400 ;
      RECT 207.9600 254.1200 210.2200 255.2000 ;
      RECT 4.8600 254.1200 205.3600 255.2000 ;
      RECT 0.0000 254.1200 2.2600 255.2000 ;
      RECT 0.0000 252.4800 210.2200 254.1200 ;
      RECT 204.9600 251.4000 210.2200 252.4800 ;
      RECT 7.8600 251.4000 202.3600 252.4800 ;
      RECT 0.0000 251.4000 5.2600 252.4800 ;
      RECT 0.0000 249.7600 210.2200 251.4000 ;
      RECT 207.9600 248.6800 210.2200 249.7600 ;
      RECT 4.8600 248.6800 205.3600 249.7600 ;
      RECT 0.0000 248.6800 2.2600 249.7600 ;
      RECT 0.0000 247.0400 210.2200 248.6800 ;
      RECT 204.9600 245.9600 210.2200 247.0400 ;
      RECT 7.8600 245.9600 202.3600 247.0400 ;
      RECT 0.0000 245.9600 5.2600 247.0400 ;
      RECT 0.0000 244.3200 210.2200 245.9600 ;
      RECT 207.9600 243.2400 210.2200 244.3200 ;
      RECT 4.8600 243.2400 205.3600 244.3200 ;
      RECT 0.0000 243.2400 2.2600 244.3200 ;
      RECT 0.0000 241.6000 210.2200 243.2400 ;
      RECT 204.9600 240.5200 210.2200 241.6000 ;
      RECT 7.8600 240.5200 202.3600 241.6000 ;
      RECT 0.0000 240.5200 5.2600 241.6000 ;
      RECT 0.0000 238.8800 210.2200 240.5200 ;
      RECT 207.9600 237.8000 210.2200 238.8800 ;
      RECT 4.8600 237.8000 205.3600 238.8800 ;
      RECT 0.0000 237.8000 2.2600 238.8800 ;
      RECT 0.0000 236.1600 210.2200 237.8000 ;
      RECT 204.9600 235.0800 210.2200 236.1600 ;
      RECT 7.8600 235.0800 202.3600 236.1600 ;
      RECT 0.0000 235.0800 5.2600 236.1600 ;
      RECT 0.0000 233.4400 210.2200 235.0800 ;
      RECT 207.9600 232.3600 210.2200 233.4400 ;
      RECT 4.8600 232.3600 205.3600 233.4400 ;
      RECT 0.0000 232.3600 2.2600 233.4400 ;
      RECT 0.0000 230.7200 210.2200 232.3600 ;
      RECT 204.9600 229.6400 210.2200 230.7200 ;
      RECT 7.8600 229.6400 202.3600 230.7200 ;
      RECT 0.0000 229.6400 5.2600 230.7200 ;
      RECT 0.0000 228.0000 210.2200 229.6400 ;
      RECT 207.9600 226.9200 210.2200 228.0000 ;
      RECT 4.8600 226.9200 205.3600 228.0000 ;
      RECT 0.0000 226.9200 2.2600 228.0000 ;
      RECT 0.0000 225.2800 210.2200 226.9200 ;
      RECT 204.9600 224.2000 210.2200 225.2800 ;
      RECT 7.8600 224.2000 202.3600 225.2800 ;
      RECT 0.0000 224.2000 5.2600 225.2800 ;
      RECT 0.0000 222.5600 210.2200 224.2000 ;
      RECT 207.9600 221.4800 210.2200 222.5600 ;
      RECT 4.8600 221.4800 205.3600 222.5600 ;
      RECT 0.0000 221.4800 2.2600 222.5600 ;
      RECT 0.0000 219.8400 210.2200 221.4800 ;
      RECT 204.9600 218.7600 210.2200 219.8400 ;
      RECT 7.8600 218.7600 202.3600 219.8400 ;
      RECT 0.0000 218.7600 5.2600 219.8400 ;
      RECT 0.0000 217.1200 210.2200 218.7600 ;
      RECT 207.9600 216.0400 210.2200 217.1200 ;
      RECT 4.8600 216.0400 205.3600 217.1200 ;
      RECT 0.0000 216.0400 2.2600 217.1200 ;
      RECT 0.0000 214.4000 210.2200 216.0400 ;
      RECT 204.9600 213.3200 210.2200 214.4000 ;
      RECT 7.8600 213.3200 202.3600 214.4000 ;
      RECT 0.0000 213.3200 5.2600 214.4000 ;
      RECT 0.0000 211.6800 210.2200 213.3200 ;
      RECT 207.9600 210.6000 210.2200 211.6800 ;
      RECT 4.8600 210.6000 205.3600 211.6800 ;
      RECT 0.0000 210.6000 2.2600 211.6800 ;
      RECT 0.0000 208.9600 210.2200 210.6000 ;
      RECT 204.9600 207.8800 210.2200 208.9600 ;
      RECT 7.8600 207.8800 202.3600 208.9600 ;
      RECT 0.0000 207.8800 5.2600 208.9600 ;
      RECT 0.0000 206.2400 210.2200 207.8800 ;
      RECT 207.9600 205.1600 210.2200 206.2400 ;
      RECT 4.8600 205.1600 205.3600 206.2400 ;
      RECT 0.0000 205.1600 2.2600 206.2400 ;
      RECT 0.0000 203.5200 210.2200 205.1600 ;
      RECT 204.9600 202.4400 210.2200 203.5200 ;
      RECT 7.8600 202.4400 202.3600 203.5200 ;
      RECT 0.0000 202.4400 5.2600 203.5200 ;
      RECT 0.0000 200.8000 210.2200 202.4400 ;
      RECT 207.9600 199.7200 210.2200 200.8000 ;
      RECT 4.8600 199.7200 205.3600 200.8000 ;
      RECT 0.0000 199.7200 2.2600 200.8000 ;
      RECT 0.0000 198.0800 210.2200 199.7200 ;
      RECT 204.9600 197.0000 210.2200 198.0800 ;
      RECT 7.8600 197.0000 202.3600 198.0800 ;
      RECT 0.0000 197.0000 5.2600 198.0800 ;
      RECT 0.0000 195.3600 210.2200 197.0000 ;
      RECT 207.9600 194.2800 210.2200 195.3600 ;
      RECT 4.8600 194.2800 205.3600 195.3600 ;
      RECT 0.0000 194.2800 2.2600 195.3600 ;
      RECT 0.0000 192.6400 210.2200 194.2800 ;
      RECT 204.9600 191.5600 210.2200 192.6400 ;
      RECT 7.8600 191.5600 202.3600 192.6400 ;
      RECT 0.0000 191.5600 5.2600 192.6400 ;
      RECT 0.0000 189.9200 210.2200 191.5600 ;
      RECT 207.9600 188.8400 210.2200 189.9200 ;
      RECT 4.8600 188.8400 205.3600 189.9200 ;
      RECT 0.0000 188.8400 2.2600 189.9200 ;
      RECT 0.0000 187.2000 210.2200 188.8400 ;
      RECT 204.9600 186.1200 210.2200 187.2000 ;
      RECT 7.8600 186.1200 202.3600 187.2000 ;
      RECT 0.0000 186.1200 5.2600 187.2000 ;
      RECT 0.0000 184.4800 210.2200 186.1200 ;
      RECT 207.9600 183.4000 210.2200 184.4800 ;
      RECT 4.8600 183.4000 205.3600 184.4800 ;
      RECT 0.0000 183.4000 2.2600 184.4800 ;
      RECT 0.0000 181.7600 210.2200 183.4000 ;
      RECT 204.9600 180.6800 210.2200 181.7600 ;
      RECT 7.8600 180.6800 202.3600 181.7600 ;
      RECT 0.0000 180.6800 5.2600 181.7600 ;
      RECT 0.0000 179.0400 210.2200 180.6800 ;
      RECT 207.9600 177.9600 210.2200 179.0400 ;
      RECT 4.8600 177.9600 205.3600 179.0400 ;
      RECT 0.0000 177.9600 2.2600 179.0400 ;
      RECT 0.0000 176.3200 210.2200 177.9600 ;
      RECT 204.9600 175.2400 210.2200 176.3200 ;
      RECT 7.8600 175.2400 202.3600 176.3200 ;
      RECT 0.0000 175.2400 5.2600 176.3200 ;
      RECT 0.0000 173.6000 210.2200 175.2400 ;
      RECT 207.9600 172.5200 210.2200 173.6000 ;
      RECT 4.8600 172.5200 205.3600 173.6000 ;
      RECT 0.0000 172.5200 2.2600 173.6000 ;
      RECT 0.0000 170.8800 210.2200 172.5200 ;
      RECT 204.9600 169.8000 210.2200 170.8800 ;
      RECT 7.8600 169.8000 202.3600 170.8800 ;
      RECT 0.0000 169.8000 5.2600 170.8800 ;
      RECT 0.0000 168.1600 210.2200 169.8000 ;
      RECT 207.9600 167.0800 210.2200 168.1600 ;
      RECT 4.8600 167.0800 205.3600 168.1600 ;
      RECT 0.0000 167.0800 2.2600 168.1600 ;
      RECT 0.0000 165.4400 210.2200 167.0800 ;
      RECT 204.9600 164.3600 210.2200 165.4400 ;
      RECT 7.8600 164.3600 202.3600 165.4400 ;
      RECT 0.0000 164.3600 5.2600 165.4400 ;
      RECT 0.0000 162.7200 210.2200 164.3600 ;
      RECT 207.9600 161.6400 210.2200 162.7200 ;
      RECT 4.8600 161.6400 205.3600 162.7200 ;
      RECT 0.0000 161.6400 2.2600 162.7200 ;
      RECT 0.0000 160.0000 210.2200 161.6400 ;
      RECT 204.9600 158.9200 210.2200 160.0000 ;
      RECT 7.8600 158.9200 202.3600 160.0000 ;
      RECT 0.0000 158.9200 5.2600 160.0000 ;
      RECT 0.0000 157.2800 210.2200 158.9200 ;
      RECT 207.9600 156.2000 210.2200 157.2800 ;
      RECT 4.8600 156.2000 205.3600 157.2800 ;
      RECT 0.0000 156.2000 2.2600 157.2800 ;
      RECT 0.0000 154.5600 210.2200 156.2000 ;
      RECT 204.9600 153.4800 210.2200 154.5600 ;
      RECT 7.8600 153.4800 202.3600 154.5600 ;
      RECT 0.0000 153.4800 5.2600 154.5600 ;
      RECT 0.0000 151.8400 210.2200 153.4800 ;
      RECT 207.9600 150.7600 210.2200 151.8400 ;
      RECT 4.8600 150.7600 205.3600 151.8400 ;
      RECT 0.0000 150.7600 2.2600 151.8400 ;
      RECT 0.0000 149.1200 210.2200 150.7600 ;
      RECT 204.9600 148.0400 210.2200 149.1200 ;
      RECT 7.8600 148.0400 202.3600 149.1200 ;
      RECT 0.0000 148.0400 5.2600 149.1200 ;
      RECT 0.0000 146.4000 210.2200 148.0400 ;
      RECT 207.9600 145.3200 210.2200 146.4000 ;
      RECT 4.8600 145.3200 205.3600 146.4000 ;
      RECT 0.0000 145.3200 2.2600 146.4000 ;
      RECT 0.0000 143.6800 210.2200 145.3200 ;
      RECT 204.9600 142.6000 210.2200 143.6800 ;
      RECT 7.8600 142.6000 202.3600 143.6800 ;
      RECT 0.0000 142.6000 5.2600 143.6800 ;
      RECT 0.0000 140.9600 210.2200 142.6000 ;
      RECT 207.9600 139.8800 210.2200 140.9600 ;
      RECT 4.8600 139.8800 205.3600 140.9600 ;
      RECT 0.0000 139.8800 2.2600 140.9600 ;
      RECT 0.0000 138.2400 210.2200 139.8800 ;
      RECT 204.9600 137.1600 210.2200 138.2400 ;
      RECT 7.8600 137.1600 202.3600 138.2400 ;
      RECT 0.0000 137.1600 5.2600 138.2400 ;
      RECT 0.0000 135.5200 210.2200 137.1600 ;
      RECT 207.9600 134.4400 210.2200 135.5200 ;
      RECT 4.8600 134.4400 205.3600 135.5200 ;
      RECT 0.0000 134.4400 2.2600 135.5200 ;
      RECT 0.0000 132.8000 210.2200 134.4400 ;
      RECT 204.9600 131.7200 210.2200 132.8000 ;
      RECT 7.8600 131.7200 202.3600 132.8000 ;
      RECT 0.0000 131.7200 5.2600 132.8000 ;
      RECT 0.0000 130.0800 210.2200 131.7200 ;
      RECT 207.9600 129.0000 210.2200 130.0800 ;
      RECT 4.8600 129.0000 205.3600 130.0800 ;
      RECT 0.0000 129.0000 2.2600 130.0800 ;
      RECT 0.0000 127.3600 210.2200 129.0000 ;
      RECT 204.9600 126.2800 210.2200 127.3600 ;
      RECT 7.8600 126.2800 202.3600 127.3600 ;
      RECT 0.0000 126.2800 5.2600 127.3600 ;
      RECT 0.0000 124.6400 210.2200 126.2800 ;
      RECT 207.9600 123.5600 210.2200 124.6400 ;
      RECT 4.8600 123.5600 205.3600 124.6400 ;
      RECT 0.0000 123.5600 2.2600 124.6400 ;
      RECT 0.0000 121.9200 210.2200 123.5600 ;
      RECT 204.9600 120.8400 210.2200 121.9200 ;
      RECT 7.8600 120.8400 202.3600 121.9200 ;
      RECT 0.0000 120.8400 5.2600 121.9200 ;
      RECT 0.0000 119.2000 210.2200 120.8400 ;
      RECT 207.9600 118.1200 210.2200 119.2000 ;
      RECT 4.8600 118.1200 205.3600 119.2000 ;
      RECT 0.0000 118.1200 2.2600 119.2000 ;
      RECT 0.0000 116.4800 210.2200 118.1200 ;
      RECT 204.9600 115.4000 210.2200 116.4800 ;
      RECT 7.8600 115.4000 202.3600 116.4800 ;
      RECT 0.0000 115.4000 5.2600 116.4800 ;
      RECT 0.0000 113.7600 210.2200 115.4000 ;
      RECT 207.9600 112.6800 210.2200 113.7600 ;
      RECT 4.8600 112.6800 205.3600 113.7600 ;
      RECT 0.0000 112.6800 2.2600 113.7600 ;
      RECT 0.0000 111.0400 210.2200 112.6800 ;
      RECT 204.9600 109.9600 210.2200 111.0400 ;
      RECT 7.8600 109.9600 202.3600 111.0400 ;
      RECT 0.0000 109.9600 5.2600 111.0400 ;
      RECT 0.0000 108.3200 210.2200 109.9600 ;
      RECT 207.9600 107.2400 210.2200 108.3200 ;
      RECT 4.8600 107.2400 205.3600 108.3200 ;
      RECT 0.0000 107.2400 2.2600 108.3200 ;
      RECT 0.0000 105.6000 210.2200 107.2400 ;
      RECT 204.9600 104.5200 210.2200 105.6000 ;
      RECT 7.8600 104.5200 202.3600 105.6000 ;
      RECT 0.0000 104.5200 5.2600 105.6000 ;
      RECT 0.0000 102.8800 210.2200 104.5200 ;
      RECT 207.9600 101.8000 210.2200 102.8800 ;
      RECT 4.8600 101.8000 205.3600 102.8800 ;
      RECT 0.0000 101.8000 2.2600 102.8800 ;
      RECT 0.0000 100.1600 210.2200 101.8000 ;
      RECT 204.9600 99.0800 210.2200 100.1600 ;
      RECT 7.8600 99.0800 202.3600 100.1600 ;
      RECT 0.0000 99.0800 5.2600 100.1600 ;
      RECT 0.0000 97.4400 210.2200 99.0800 ;
      RECT 207.9600 96.3600 210.2200 97.4400 ;
      RECT 4.8600 96.3600 205.3600 97.4400 ;
      RECT 0.0000 96.3600 2.2600 97.4400 ;
      RECT 0.0000 94.7200 210.2200 96.3600 ;
      RECT 204.9600 93.6400 210.2200 94.7200 ;
      RECT 7.8600 93.6400 202.3600 94.7200 ;
      RECT 0.0000 93.6400 5.2600 94.7200 ;
      RECT 0.0000 92.0000 210.2200 93.6400 ;
      RECT 207.9600 90.9200 210.2200 92.0000 ;
      RECT 4.8600 90.9200 205.3600 92.0000 ;
      RECT 0.0000 90.9200 2.2600 92.0000 ;
      RECT 0.0000 89.2800 210.2200 90.9200 ;
      RECT 204.9600 88.2000 210.2200 89.2800 ;
      RECT 7.8600 88.2000 202.3600 89.2800 ;
      RECT 0.0000 88.2000 5.2600 89.2800 ;
      RECT 0.0000 86.5600 210.2200 88.2000 ;
      RECT 207.9600 85.4800 210.2200 86.5600 ;
      RECT 4.8600 85.4800 205.3600 86.5600 ;
      RECT 0.0000 85.4800 2.2600 86.5600 ;
      RECT 0.0000 83.8400 210.2200 85.4800 ;
      RECT 204.9600 82.7600 210.2200 83.8400 ;
      RECT 7.8600 82.7600 202.3600 83.8400 ;
      RECT 0.0000 82.7600 5.2600 83.8400 ;
      RECT 0.0000 81.1200 210.2200 82.7600 ;
      RECT 207.9600 80.0400 210.2200 81.1200 ;
      RECT 4.8600 80.0400 205.3600 81.1200 ;
      RECT 0.0000 80.0400 2.2600 81.1200 ;
      RECT 0.0000 78.4000 210.2200 80.0400 ;
      RECT 204.9600 77.3200 210.2200 78.4000 ;
      RECT 7.8600 77.3200 202.3600 78.4000 ;
      RECT 0.0000 77.3200 5.2600 78.4000 ;
      RECT 0.0000 75.6800 210.2200 77.3200 ;
      RECT 207.9600 74.6000 210.2200 75.6800 ;
      RECT 4.8600 74.6000 205.3600 75.6800 ;
      RECT 0.0000 74.6000 2.2600 75.6800 ;
      RECT 0.0000 72.9600 210.2200 74.6000 ;
      RECT 204.9600 71.8800 210.2200 72.9600 ;
      RECT 7.8600 71.8800 202.3600 72.9600 ;
      RECT 0.0000 71.8800 5.2600 72.9600 ;
      RECT 0.0000 70.2400 210.2200 71.8800 ;
      RECT 207.9600 69.1600 210.2200 70.2400 ;
      RECT 4.8600 69.1600 205.3600 70.2400 ;
      RECT 0.0000 69.1600 2.2600 70.2400 ;
      RECT 0.0000 67.5200 210.2200 69.1600 ;
      RECT 204.9600 66.4400 210.2200 67.5200 ;
      RECT 7.8600 66.4400 202.3600 67.5200 ;
      RECT 0.0000 66.4400 5.2600 67.5200 ;
      RECT 0.0000 64.8000 210.2200 66.4400 ;
      RECT 207.9600 63.7200 210.2200 64.8000 ;
      RECT 4.8600 63.7200 205.3600 64.8000 ;
      RECT 0.0000 63.7200 2.2600 64.8000 ;
      RECT 0.0000 62.0800 210.2200 63.7200 ;
      RECT 204.9600 61.0000 210.2200 62.0800 ;
      RECT 7.8600 61.0000 202.3600 62.0800 ;
      RECT 0.0000 61.0000 5.2600 62.0800 ;
      RECT 0.0000 59.3600 210.2200 61.0000 ;
      RECT 207.9600 58.2800 210.2200 59.3600 ;
      RECT 4.8600 58.2800 205.3600 59.3600 ;
      RECT 0.0000 58.2800 2.2600 59.3600 ;
      RECT 0.0000 56.6400 210.2200 58.2800 ;
      RECT 204.9600 55.5600 210.2200 56.6400 ;
      RECT 7.8600 55.5600 202.3600 56.6400 ;
      RECT 0.0000 55.5600 5.2600 56.6400 ;
      RECT 0.0000 53.9200 210.2200 55.5600 ;
      RECT 207.9600 52.8400 210.2200 53.9200 ;
      RECT 4.8600 52.8400 205.3600 53.9200 ;
      RECT 0.0000 52.8400 2.2600 53.9200 ;
      RECT 0.0000 51.2000 210.2200 52.8400 ;
      RECT 204.9600 50.1200 210.2200 51.2000 ;
      RECT 7.8600 50.1200 202.3600 51.2000 ;
      RECT 0.0000 50.1200 5.2600 51.2000 ;
      RECT 0.0000 48.4800 210.2200 50.1200 ;
      RECT 207.9600 47.4000 210.2200 48.4800 ;
      RECT 4.8600 47.4000 205.3600 48.4800 ;
      RECT 0.0000 47.4000 2.2600 48.4800 ;
      RECT 0.0000 45.7600 210.2200 47.4000 ;
      RECT 204.9600 44.6800 210.2200 45.7600 ;
      RECT 7.8600 44.6800 202.3600 45.7600 ;
      RECT 0.0000 44.6800 5.2600 45.7600 ;
      RECT 0.0000 43.0400 210.2200 44.6800 ;
      RECT 207.9600 41.9600 210.2200 43.0400 ;
      RECT 4.8600 41.9600 205.3600 43.0400 ;
      RECT 0.0000 41.9600 2.2600 43.0400 ;
      RECT 0.0000 40.3200 210.2200 41.9600 ;
      RECT 204.9600 39.2400 210.2200 40.3200 ;
      RECT 7.8600 39.2400 202.3600 40.3200 ;
      RECT 0.0000 39.2400 5.2600 40.3200 ;
      RECT 0.0000 37.6000 210.2200 39.2400 ;
      RECT 207.9600 36.5200 210.2200 37.6000 ;
      RECT 4.8600 36.5200 205.3600 37.6000 ;
      RECT 0.0000 36.5200 2.2600 37.6000 ;
      RECT 0.0000 34.8800 210.2200 36.5200 ;
      RECT 204.9600 33.8000 210.2200 34.8800 ;
      RECT 7.8600 33.8000 202.3600 34.8800 ;
      RECT 0.0000 33.8000 5.2600 34.8800 ;
      RECT 0.0000 32.1600 210.2200 33.8000 ;
      RECT 207.9600 31.0800 210.2200 32.1600 ;
      RECT 4.8600 31.0800 205.3600 32.1600 ;
      RECT 0.0000 31.0800 2.2600 32.1600 ;
      RECT 0.0000 29.4400 210.2200 31.0800 ;
      RECT 204.9600 28.3600 210.2200 29.4400 ;
      RECT 7.8600 28.3600 202.3600 29.4400 ;
      RECT 0.0000 28.3600 5.2600 29.4400 ;
      RECT 0.0000 26.7200 210.2200 28.3600 ;
      RECT 207.9600 25.6400 210.2200 26.7200 ;
      RECT 4.8600 25.6400 205.3600 26.7200 ;
      RECT 0.0000 25.6400 2.2600 26.7200 ;
      RECT 0.0000 24.0000 210.2200 25.6400 ;
      RECT 204.9600 22.9200 210.2200 24.0000 ;
      RECT 7.8600 22.9200 202.3600 24.0000 ;
      RECT 0.0000 22.9200 5.2600 24.0000 ;
      RECT 0.0000 21.2800 210.2200 22.9200 ;
      RECT 207.9600 20.2000 210.2200 21.2800 ;
      RECT 4.8600 20.2000 205.3600 21.2800 ;
      RECT 0.0000 20.2000 2.2600 21.2800 ;
      RECT 0.0000 18.5600 210.2200 20.2000 ;
      RECT 204.9600 17.4800 210.2200 18.5600 ;
      RECT 7.8600 17.4800 202.3600 18.5600 ;
      RECT 0.0000 17.4800 5.2600 18.5600 ;
      RECT 0.0000 15.8400 210.2200 17.4800 ;
      RECT 207.9600 14.7600 210.2200 15.8400 ;
      RECT 4.8600 14.7600 205.3600 15.8400 ;
      RECT 0.0000 14.7600 2.2600 15.8400 ;
      RECT 0.0000 13.1200 210.2200 14.7600 ;
      RECT 204.9600 12.0400 210.2200 13.1200 ;
      RECT 7.8600 12.0400 202.3600 13.1200 ;
      RECT 0.0000 12.0400 5.2600 13.1200 ;
      RECT 0.0000 10.4000 210.2200 12.0400 ;
      RECT 207.9600 9.3200 210.2200 10.4000 ;
      RECT 4.8600 9.3200 205.3600 10.4000 ;
      RECT 0.0000 9.3200 2.2600 10.4000 ;
      RECT 0.0000 7.7300 210.2200 9.3200 ;
      RECT 204.9600 5.1300 210.2200 7.7300 ;
      RECT 0.0000 5.1300 5.2600 7.7300 ;
      RECT 0.0000 4.7300 210.2200 5.1300 ;
      RECT 207.9600 2.1300 210.2200 4.7300 ;
      RECT 0.0000 2.1300 2.2600 4.7300 ;
      RECT 0.0000 0.0000 210.2200 2.1300 ;
    LAYER met4 ;
      RECT 0.0000 442.2500 210.2200 444.7200 ;
      RECT 195.2200 439.2500 205.3600 442.2500 ;
      RECT 150.2200 439.2500 193.0200 442.2500 ;
      RECT 105.2200 439.2500 148.0200 442.2500 ;
      RECT 60.2200 439.2500 103.0200 442.2500 ;
      RECT 15.2200 439.2500 58.0200 442.2500 ;
      RECT 4.8600 439.2500 13.0200 442.2500 ;
      RECT 204.9600 5.1300 205.3600 439.2500 ;
      RECT 195.2200 5.1300 202.3600 439.2500 ;
      RECT 192.0200 5.1300 193.0200 439.2500 ;
      RECT 150.2200 5.1300 189.8200 439.2500 ;
      RECT 147.0200 5.1300 148.0200 439.2500 ;
      RECT 105.2200 5.1300 144.8200 439.2500 ;
      RECT 102.0200 5.1300 103.0200 439.2500 ;
      RECT 60.2200 5.1300 99.8200 439.2500 ;
      RECT 57.0200 5.1300 58.0200 439.2500 ;
      RECT 15.2200 5.1300 54.8200 439.2500 ;
      RECT 12.0200 5.1300 13.0200 439.2500 ;
      RECT 7.8600 5.1300 9.8200 439.2500 ;
      RECT 4.8600 5.1300 5.2600 439.2500 ;
      RECT 207.9600 2.1300 210.2200 442.2500 ;
      RECT 195.2200 2.1300 205.3600 5.1300 ;
      RECT 150.2200 2.1300 193.0200 5.1300 ;
      RECT 105.2200 2.1300 148.0200 5.1300 ;
      RECT 60.2200 2.1300 103.0200 5.1300 ;
      RECT 15.2200 2.1300 58.0200 5.1300 ;
      RECT 4.8600 2.1300 13.0200 5.1300 ;
      RECT 0.0000 2.1300 2.2600 442.2500 ;
      RECT 0.0000 1.1000 210.2200 2.1300 ;
      RECT 90.1500 0.0000 210.2200 1.1000 ;
      RECT 0.0000 0.0000 89.2500 1.1000 ;
  END
END DSP

END LIBRARY
