magic
tech sky130B
magscale 1 2
timestamp 1707688321
<< pwell >>
rect -76 -26 256 2026
<< mvnnmos >>
rect 0 0 180 2000
<< mvndiff >>
rect -50 0 0 2000
rect 180 0 230 2000
<< poly >>
rect 0 2000 180 2032
rect 0 -32 180 0
<< locali >>
rect -45 -4 -11 1966
rect 191 -4 225 1966
use DFL1sd_CDNS_52468879185709  DFL1sd_CDNS_52468879185709_0
timestamp 1707688321
transform -1 0 0 0 1 0
box -26 -26 79 2026
use DFL1sd_CDNS_52468879185709  DFL1sd_CDNS_52468879185709_1
timestamp 1707688321
transform 1 0 180 0 1 0
box -26 -26 79 2026
<< labels >>
flabel comment s -28 981 -28 981 0 FreeSans 300 0 0 0 S
flabel comment s 208 981 208 981 0 FreeSans 300 0 0 0 D
<< properties >>
string GDS_END 86613718
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 86612768
<< end >>
