magic
tech sky130B
magscale 1 2
timestamp 1707688321
<< locali >>
rect 66 2732 168 2798
rect 227 2699 293 2797
rect 222 2672 293 2699
rect 222 2638 264 2672
rect 99 2372 133 2410
rect 474 2372 508 2410
rect 12 1840 46 1878
rect 650 1840 684 1878
rect 702 1484 808 1516
rect 736 1450 774 1484
rect 99 1367 137 1401
rect 65 1282 171 1367
rect 378 918 412 1450
rect 528 1416 630 1450
rect 842 1416 876 2699
rect 1378 1450 1412 1556
rect 2001 1450 2035 1556
rect 188 846 222 884
rect 398 884 412 918
rect 364 846 412 884
rect 398 812 412 846
rect 460 1382 630 1416
rect 704 1382 876 1416
rect 1138 1416 1412 1450
rect 1764 1416 2035 1450
rect 460 918 494 1382
rect 704 1348 806 1382
rect 1138 1348 1172 1416
rect 1764 1348 1798 1416
rect 1648 1282 1798 1348
rect 460 884 474 918
rect 460 846 508 884
rect 460 812 474 846
rect 1764 917 1798 1282
rect 650 846 684 884
rect 932 845 966 883
rect 1764 883 1769 917
rect 1764 845 1803 883
rect 826 770 860 808
rect 1206 770 1240 808
rect 1492 770 1526 808
rect 1764 811 1769 845
rect 1403 308 1437 346
rect 1668 308 1702 346
rect 1316 150 1350 188
rect 1764 99 1798 811
rect 238 49 242 66
rect 272 15 310 49
rect 558 32 596 66
rect 238 0 242 15
rect 524 0 528 32
rect 1832 0 1934 66
rect 66 -37 168 0
rect 100 -71 138 -37
<< viali >>
rect 99 2410 133 2444
rect 99 2338 133 2372
rect 474 2410 508 2444
rect 474 2338 508 2372
rect 12 1878 46 1912
rect 12 1806 46 1840
rect 650 1878 684 1912
rect 650 1806 684 1840
rect 702 1450 736 1484
rect 774 1450 808 1484
rect 65 1367 99 1401
rect 137 1367 171 1401
rect 188 884 222 918
rect 188 812 222 846
rect 364 884 398 918
rect 364 812 398 846
rect 474 884 508 918
rect 474 812 508 846
rect 650 884 684 918
rect 650 812 684 846
rect 932 883 966 917
rect 826 808 860 842
rect 932 811 966 845
rect 1769 883 1803 917
rect 826 736 860 770
rect 1206 808 1240 842
rect 1206 736 1240 770
rect 1492 808 1526 842
rect 1492 736 1526 770
rect 1769 811 1803 845
rect 1403 346 1437 380
rect 1403 274 1437 308
rect 1668 346 1702 380
rect 1668 274 1702 308
rect 1316 188 1350 222
rect 1316 116 1350 150
rect 238 15 272 49
rect 310 15 344 49
rect 524 32 558 66
rect 596 32 630 66
rect 66 -71 100 -37
rect 138 -71 172 -37
<< metal1 >>
rect 93 2444 139 2456
rect 93 2410 99 2444
rect 133 2410 139 2444
rect 93 2378 139 2410
rect 468 2444 514 2456
rect 468 2410 474 2444
rect 508 2410 514 2444
tri 139 2378 164 2403 sw
tri 443 2378 468 2403 se
rect 468 2378 514 2410
rect 93 2372 514 2378
rect 93 2338 99 2372
rect 133 2338 474 2372
rect 508 2338 514 2372
rect 93 2326 514 2338
rect 0 2096 29 2298
rect 205 2096 286 2298
rect 843 2096 942 2298
rect 2038 2110 2067 2298
rect 0 2022 942 2096
rect 0 1912 58 1918
rect 0 1878 12 1912
rect 46 1878 58 1912
rect 638 1912 696 1918
tri 58 1878 74 1894 sw
rect 638 1878 650 1912
rect 684 1878 696 1912
rect 0 1871 74 1878
tri 74 1871 81 1878 sw
rect 0 1846 81 1871
tri 81 1846 106 1871 sw
tri 613 1846 638 1871 se
rect 0 1840 58 1846
rect 0 1806 12 1840
rect 46 1806 58 1840
rect 0 1800 58 1806
rect 205 1800 286 1846
rect 638 1840 696 1878
tri 696 1846 721 1871 sw
rect 638 1806 650 1840
rect 684 1806 696 1840
rect 638 1800 696 1806
rect 843 1800 936 1846
rect 2052 1800 2082 1846
rect 0 1772 2082 1800
rect 0 1570 29 1772
rect 205 1570 286 1772
rect 843 1570 936 1772
rect 2184 1570 2214 1772
rect 690 1484 820 1490
rect 690 1450 702 1484
rect 736 1450 774 1484
rect 808 1450 820 1484
tri 665 1407 690 1432 se
rect 690 1407 820 1450
rect 53 1401 820 1407
rect 53 1367 65 1401
rect 99 1367 137 1401
rect 171 1367 820 1401
rect 53 1361 820 1367
rect 0 1026 29 1228
rect 410 1026 462 1228
rect 1252 1026 1333 1228
rect 1685 1026 1795 1228
rect 1971 1026 2000 1228
rect 0 998 2000 1026
rect 0 952 29 998
rect 410 952 462 998
rect 1252 952 1333 998
rect 1685 952 1795 998
rect 1971 952 2000 998
rect 176 918 234 924
rect 176 884 188 918
rect 222 884 234 918
rect 176 846 234 884
rect 352 918 410 924
rect 352 884 364 918
rect 398 884 410 918
tri 234 853 259 878 nw
tri 327 853 352 878 ne
rect 176 812 188 846
rect 222 812 234 846
rect 176 806 234 812
rect 352 846 410 884
rect 352 812 364 846
rect 398 812 410 846
rect 352 806 410 812
rect 462 918 520 924
rect 462 884 474 918
rect 508 884 520 918
rect 462 846 520 884
rect 638 918 696 924
rect 638 884 650 918
rect 684 884 696 918
tri 520 853 545 878 nw
tri 613 853 638 878 ne
rect 462 812 474 846
rect 508 812 520 846
rect 462 806 520 812
rect 638 846 696 884
rect 920 917 1815 923
rect 920 883 932 917
rect 966 895 1769 917
rect 966 883 991 895
tri 991 883 1003 895 nw
tri 1732 883 1744 895 ne
rect 1744 883 1769 895
rect 1803 883 1815 917
rect 638 812 650 846
rect 684 812 696 846
rect 638 806 696 812
rect 814 842 872 848
rect 814 808 826 842
rect 860 808 872 842
tri 789 776 814 801 se
rect 0 730 29 776
rect 410 730 462 776
rect 814 770 872 808
rect 920 845 978 883
tri 978 870 991 883 nw
tri 1744 870 1757 883 ne
rect 920 811 932 845
rect 966 811 978 845
rect 920 805 978 811
rect 1194 842 1252 848
rect 1194 808 1206 842
rect 1240 808 1252 842
tri 872 776 897 801 sw
tri 1169 776 1194 801 se
rect 1194 776 1252 808
rect 1480 842 1538 848
rect 1480 808 1492 842
rect 1526 808 1538 842
tri 1252 776 1277 801 sw
tri 1455 776 1480 801 se
rect 814 736 826 770
rect 860 736 872 770
rect 814 730 872 736
rect 1194 770 1333 776
rect 1194 736 1206 770
rect 1240 736 1333 770
rect 1194 730 1333 736
rect 1480 770 1538 808
rect 1757 845 1815 883
rect 1757 811 1769 845
rect 1803 811 1815 845
rect 1757 805 1815 811
tri 1538 776 1563 801 sw
rect 1480 736 1492 770
rect 1526 736 1538 770
rect 1480 730 1538 736
rect 1685 730 1795 776
rect 1971 730 2000 776
rect 0 702 2000 730
rect -2335 622 -2133 642
rect -2105 622 -2059 642
rect -1792 616 -1607 642
rect 0 500 29 702
rect 410 500 462 702
rect 1252 500 1333 702
rect 1685 500 1795 702
rect 1971 500 2000 702
rect 0 420 2000 472
tri 985 395 1010 420 ne
tri 1246 395 1271 420 nw
rect 1397 380 1443 392
rect 1397 346 1403 380
rect 1437 346 1443 380
tri 1372 314 1397 339 se
rect 1397 314 1443 346
rect 1662 380 1708 392
rect 1662 346 1668 380
rect 1702 346 1708 380
tri 1443 314 1468 339 sw
tri 1637 314 1662 339 se
rect 1662 314 1708 346
tri 1708 314 1733 339 sw
rect 0 308 2000 314
rect 0 274 1403 308
rect 1437 274 1668 308
rect 1702 274 2000 308
rect 0 262 2000 274
rect 0 222 2000 234
rect 0 188 1316 222
rect 1350 188 2000 222
rect 0 182 2000 188
tri 1285 157 1310 182 ne
rect 1310 150 1356 182
tri 1356 157 1381 182 nw
tri 36 119 42 125 se
rect 42 119 454 125
tri 454 119 460 125 sw
tri 33 116 36 119 se
rect 36 116 460 119
tri 460 116 463 119 sw
rect 1310 116 1316 150
rect 1350 116 1356 150
tri 1 84 33 116 se
rect 33 104 463 116
tri 463 104 475 116 sw
rect 1310 104 1356 116
rect 33 97 475 104
rect 33 84 42 97
tri 42 84 55 97 nw
tri 441 84 454 97 ne
rect 454 84 475 97
tri -5 78 1 84 se
rect 1 78 36 84
tri 36 78 42 84 nw
tri 454 78 460 84 ne
rect 460 78 475 84
tri 475 78 501 104 sw
tri -17 66 -5 78 se
rect -5 66 24 78
tri 24 66 36 78 nw
tri 460 66 472 78 ne
rect 472 66 636 78
tri -22 61 -17 66 se
rect -17 61 19 66
tri 19 61 24 66 nw
tri 472 61 477 66 ne
rect 477 61 524 66
tri -34 49 -22 61 se
rect -22 49 7 61
tri 7 49 19 61 nw
tri 220 49 232 61 se
rect 232 49 350 61
tri -40 43 -34 49 se
rect -34 43 1 49
tri 1 43 7 49 nw
tri 214 43 220 49 se
rect 220 43 238 49
tri -47 36 -40 43 se
rect -40 36 -6 43
tri -6 36 1 43 nw
tri 207 36 214 43 se
rect 214 36 238 43
rect -75 31 -11 36
tri -11 31 -6 36 nw
tri 202 31 207 36 se
rect 207 31 238 36
rect -75 30 -12 31
tri -12 30 -11 31 nw
tri 28 30 29 31 se
rect 29 30 238 31
rect -75 15 -27 30
tri -27 15 -12 30 nw
tri 13 15 28 30 se
rect 28 15 238 30
rect 272 15 310 49
rect 344 15 350 49
tri 477 32 506 61 ne
rect 506 32 524 61
rect 558 32 596 66
rect 630 32 636 66
tri 506 20 518 32 ne
rect 518 20 636 32
rect -75 8 -34 15
tri -34 8 -27 15 nw
tri 6 8 13 15 se
rect 13 8 350 15
tri 1 3 6 8 se
rect 6 3 350 8
tri -12 -10 1 3 se
rect 1 -10 29 3
tri 29 -10 42 3 nw
tri -27 -25 -12 -10 se
rect -12 -25 14 -10
tri 14 -25 29 -10 nw
tri -31 -29 -27 -25 se
rect -27 -29 10 -25
tri 10 -29 14 -25 nw
rect -75 -37 2 -29
tri 2 -37 10 -29 nw
rect 60 -37 182 -25
rect -75 -57 -18 -37
tri -18 -57 2 -37 nw
rect 60 -71 66 -37
rect 100 -71 138 -37
rect 172 -71 182 -37
rect 60 -82 182 -71
tri 182 -82 239 -25 sw
rect 60 -83 239 -82
tri 239 -83 240 -82 sw
tri 194 -128 239 -83 ne
rect 239 -88 240 -83
tri 240 -88 245 -83 sw
rect 239 -128 245 -88
tri 245 -128 285 -88 sw
tri 1761 -128 1801 -88 se
rect 1801 -120 2147 -88
tri 239 -174 285 -128 ne
tri 285 -134 291 -128 sw
tri 1755 -134 1761 -128 se
rect 1761 -134 1801 -128
tri 1801 -134 1815 -120 nw
rect 285 -174 291 -134
tri 291 -174 331 -134 sw
tri 1715 -174 1755 -134 se
rect 1755 -174 1761 -134
tri 1761 -174 1801 -134 nw
tri 285 -206 317 -174 ne
rect 317 -206 1729 -174
tri 1729 -206 1761 -174 nw
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_0
timestamp 1707688321
transform 0 1 66 -1 0 -37
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_1
timestamp 1707688321
transform 0 1 238 -1 0 49
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_2
timestamp 1707688321
transform 0 1 524 -1 0 66
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_3
timestamp 1707688321
transform -1 0 222 0 1 812
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_4
timestamp 1707688321
transform -1 0 1803 0 1 811
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_5
timestamp 1707688321
transform -1 0 966 0 1 811
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_6
timestamp 1707688321
transform -1 0 860 0 1 736
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_7
timestamp 1707688321
transform -1 0 1240 0 1 736
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_8
timestamp 1707688321
transform -1 0 1526 0 1 736
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_9
timestamp 1707688321
transform 1 0 12 0 -1 1912
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_10
timestamp 1707688321
transform 1 0 650 0 -1 1912
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_11
timestamp 1707688321
transform 1 0 364 0 1 812
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_12
timestamp 1707688321
transform 1 0 474 0 1 812
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_13
timestamp 1707688321
transform 1 0 650 0 1 812
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_0
timestamp 1707688321
transform 0 -1 508 1 0 2338
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_1
timestamp 1707688321
transform 0 -1 133 1 0 2338
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_2
timestamp 1707688321
transform 0 -1 1702 1 0 274
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_3
timestamp 1707688321
transform 0 -1 1437 1 0 274
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_4
timestamp 1707688321
transform 0 -1 1350 1 0 116
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_5
timestamp 1707688321
transform 1 0 65 0 1 1367
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_6
timestamp 1707688321
transform 1 0 702 0 1 1450
box 0 0 1 1
use sky130_fd_io__sio_hotswap_dly  sky130_fd_io__sio_hotswap_dly_0
timestamp 1707688321
transform -1 0 2302 0 1 1522
box 88 -936 4685 922
use sky130_fd_io__sio_hvsbt_inv_x1  sky130_fd_io__sio_hvsbt_inv_x1_0
timestamp 1707688321
transform -1 0 1971 0 -1 1369
box -107 21 267 1369
use sky130_fd_io__sio_hvsbt_inv_x1  sky130_fd_io__sio_hvsbt_inv_x1_1
timestamp 1707688321
transform -1 0 1509 0 -1 1369
box -107 21 267 1369
use sky130_fd_io__sio_hvsbt_inv_x1  sky130_fd_io__sio_hvsbt_inv_x1_2
timestamp 1707688321
transform 1 0 1509 0 -1 1369
box -107 21 267 1369
use sky130_fd_io__sio_hvsbt_inv_x1  sky130_fd_io__sio_hvsbt_inv_x1_3
timestamp 1707688321
transform 1 0 29 0 1 1429
box -107 21 267 1369
use sky130_fd_io__sio_hvsbt_inv_x1  sky130_fd_io__sio_hvsbt_inv_x1_4
timestamp 1707688321
transform 1 0 667 0 1 1429
box -107 21 267 1369
use sky130_fd_io__sio_hvsbt_nand2  sky130_fd_io__sio_hvsbt_nand2_0
timestamp 1707688321
transform -1 0 667 0 1 1429
box -107 21 459 1369
use sky130_fd_io__sio_hvsbt_nand2  sky130_fd_io__sio_hvsbt_nand2_1
timestamp 1707688321
transform -1 0 843 0 -1 1369
box -107 21 459 1369
use sky130_fd_io__sio_hvsbt_nand2  sky130_fd_io__sio_hvsbt_nand2_2
timestamp 1707688321
transform 1 0 29 0 -1 1369
box -107 21 459 1369
use sky130_fd_io__sio_hvsbt_nor  sky130_fd_io__sio_hvsbt_nor_0
timestamp 1707688321
transform 1 0 843 0 -1 1369
box -107 21 487 1369
<< labels >>
flabel metal1 s -2105 622 -2059 642 0 FreeSans 200 180 0 0 vgnd
port 1 nsew
flabel metal1 s 916 1800 936 1846 0 FreeSans 200 180 0 0 vgnd
port 1 nsew
flabel metal1 s 2052 1800 2082 1846 0 FreeSans 200 180 0 0 vgnd
port 1 nsew
flabel metal1 s -2335 622 -2133 642 0 FreeSans 200 180 0 0 vgnd
port 1 nsew
flabel metal1 s 2184 1570 2214 1772 0 FreeSans 300 180 0 0 vgnd
port 1 nsew
flabel metal1 s 916 1570 936 1772 0 FreeSans 200 180 0 0 vgnd
port 1 nsew
flabel metal1 s -1792 616 -1607 642 0 FreeSans 200 180 0 0 vcc_io
port 2 nsew
flabel metal1 s 916 2022 942 2298 0 FreeSans 200 180 0 0 vcc_io
port 2 nsew
flabel metal1 s 2038 2110 2067 2298 0 FreeSans 200 180 0 0 vcc_io
port 2 nsew
flabel metal1 s 1848 2070 1848 2070 0 FreeSans 100 0 0 0 enhs_dly_h
flabel metal1 s 1954 420 2000 472 0 FreeSans 200 0 0 0 exiths_h
port 3 nsew
flabel metal1 s 0 420 46 472 0 FreeSans 200 0 0 0 exiths_h
port 3 nsew
flabel metal1 s 0 262 46 314 0 FreeSans 200 0 0 0 enhs_h_n
port 4 nsew
flabel metal1 s 1954 262 2000 314 0 FreeSans 200 0 0 0 enhs_h_n
port 4 nsew
flabel metal1 s 1954 182 2000 234 0 FreeSans 200 0 0 0 enhs_h
port 5 nsew
flabel metal1 s 0 182 46 234 0 FreeSans 200 0 0 0 enhs_h
port 5 nsew
flabel metal1 s 0 952 29 998 0 FreeSans 200 0 0 0 vgnd
port 1 nsew
flabel metal1 s 0 1800 29 1846 0 FreeSans 200 0 0 0 vgnd
port 1 nsew
flabel metal1 s 2199 1671 2199 1671 0 FreeSans 200 0 0 0 vgnd
flabel metal1 s 0 1570 29 1772 0 FreeSans 200 0 0 0 vgnd
port 1 nsew
flabel metal1 s 0 1026 29 1228 0 FreeSans 200 0 0 0 vgnd
port 1 nsew
flabel metal1 s 1971 1026 2000 1228 0 FreeSans 200 0 0 0 vgnd
port 1 nsew
flabel metal1 s 1971 500 2000 776 0 FreeSans 200 0 0 0 vcc_io
port 2 nsew
flabel metal1 s 0 500 29 776 0 FreeSans 200 0 0 0 vcc_io
port 2 nsew
flabel metal1 s 2053 2204 2053 2204 0 FreeSans 200 0 0 0 vcc_io
flabel metal1 s 2045 -120 2147 -88 0 FreeSans 200 0 0 0 od_h
port 6 nsew
flabel metal1 s -75 -57 -33 -29 0 FreeSans 200 0 0 0 forcehi_h<1>
port 7 nsew
flabel metal1 s -75 8 -36 36 0 FreeSans 200 0 0 0 en_h
port 8 nsew
flabel metal1 s 1971 952 2000 998 0 FreeSans 200 0 0 0 vgnd
port 1 nsew
flabel locali s 1284 1435 1284 1435 0 FreeSans 200 0 0 0 enhs_dly_h_n
flabel locali s 66 2732 168 2798 0 FreeSans 200 0 0 0 dishs_h
port 10 nsew
flabel locali s 1832 0 1934 66 0 FreeSans 200 0 0 0 enhs_lat_h_n
port 11 nsew
flabel locali s 227 2736 293 2797 0 FreeSans 200 0 0 0 dishs_h_n
port 12 nsew
<< properties >>
string GDS_END 88554750
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 88544216
<< end >>
