magic
tech sky130A
magscale 1 2
timestamp 1707688321
<< nwell >>
rect -266 -66 219 216
<< mvpmos >>
rect 0 0 100 150
<< mvpdiff >>
rect -50 0 0 150
rect 100 114 153 150
rect 100 80 111 114
rect 145 80 153 114
rect 100 46 153 80
rect 100 12 111 46
rect 145 12 153 46
rect 100 0 153 12
<< mvpdiffc >>
rect 111 80 145 114
rect 111 12 145 46
<< poly >>
rect 0 150 100 182
rect 0 -32 100 0
<< locali >>
rect -113 -4 -11 142
rect 111 114 145 130
rect 111 46 145 80
rect 111 -4 145 12
use DFL1sd_CDNS_5246887918546  DFL1sd_CDNS_5246887918546_0
timestamp 1707688321
transform 1 0 100 0 1 0
box 0 0 1 1
use hvDFTPL1s_CDNS_52468879185912  hvDFTPL1s_CDNS_52468879185912_0
timestamp 1707688321
transform -1 0 0 0 1 0
box -36 -36 236 186
<< labels >>
flabel comment s -62 69 -62 69 0 FreeSans 300 0 0 0 S
flabel comment s 128 63 128 63 0 FreeSans 300 0 0 0 D
<< properties >>
string GDS_END 80654564
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 80653546
<< end >>
