magic
tech sky130A
magscale 1 2
timestamp 1707688321
<< nwell >>
rect -38 261 1326 582
<< pwell >>
rect 1 21 1215 203
rect 30 -17 64 21
<< scnmos >>
rect 79 47 109 177
rect 267 47 297 177
rect 351 47 381 177
rect 435 47 465 177
rect 519 47 549 177
rect 603 47 633 177
rect 687 47 717 177
rect 771 47 801 177
rect 855 47 885 177
rect 939 47 969 177
rect 1023 47 1053 177
rect 1107 47 1137 177
<< scpmoshvt >>
rect 79 297 109 497
rect 267 297 297 497
rect 351 297 381 497
rect 435 297 465 497
rect 519 297 549 497
rect 603 297 633 497
rect 687 297 717 497
rect 771 297 801 497
rect 855 297 885 497
rect 939 297 969 497
rect 1023 297 1053 497
rect 1107 297 1137 497
<< ndiff >>
rect 27 165 79 177
rect 27 131 35 165
rect 69 131 79 165
rect 27 97 79 131
rect 27 63 35 97
rect 69 63 79 97
rect 27 47 79 63
rect 109 165 161 177
rect 109 131 119 165
rect 153 131 161 165
rect 109 97 161 131
rect 109 63 119 97
rect 153 63 161 97
rect 109 47 161 63
rect 215 165 267 177
rect 215 131 223 165
rect 257 131 267 165
rect 215 97 267 131
rect 215 63 223 97
rect 257 63 267 97
rect 215 47 267 63
rect 297 97 351 177
rect 297 63 307 97
rect 341 63 351 97
rect 297 47 351 63
rect 381 165 435 177
rect 381 131 391 165
rect 425 131 435 165
rect 381 97 435 131
rect 381 63 391 97
rect 425 63 435 97
rect 381 47 435 63
rect 465 97 519 177
rect 465 63 475 97
rect 509 63 519 97
rect 465 47 519 63
rect 549 165 603 177
rect 549 131 559 165
rect 593 131 603 165
rect 549 97 603 131
rect 549 63 559 97
rect 593 63 603 97
rect 549 47 603 63
rect 633 97 687 177
rect 633 63 643 97
rect 677 63 687 97
rect 633 47 687 63
rect 717 165 771 177
rect 717 131 727 165
rect 761 131 771 165
rect 717 97 771 131
rect 717 63 727 97
rect 761 63 771 97
rect 717 47 771 63
rect 801 97 855 177
rect 801 63 811 97
rect 845 63 855 97
rect 801 47 855 63
rect 885 165 939 177
rect 885 131 895 165
rect 929 131 939 165
rect 885 97 939 131
rect 885 63 895 97
rect 929 63 939 97
rect 885 47 939 63
rect 969 97 1023 177
rect 969 63 979 97
rect 1013 63 1023 97
rect 969 47 1023 63
rect 1053 165 1107 177
rect 1053 131 1063 165
rect 1097 131 1107 165
rect 1053 97 1107 131
rect 1053 63 1063 97
rect 1097 63 1107 97
rect 1053 47 1107 63
rect 1137 97 1189 177
rect 1137 63 1147 97
rect 1181 63 1189 97
rect 1137 47 1189 63
<< pdiff >>
rect 27 485 79 497
rect 27 451 35 485
rect 69 451 79 485
rect 27 417 79 451
rect 27 383 35 417
rect 69 383 79 417
rect 27 349 79 383
rect 27 315 35 349
rect 69 315 79 349
rect 27 297 79 315
rect 109 479 161 497
rect 109 445 119 479
rect 153 445 161 479
rect 109 411 161 445
rect 109 377 119 411
rect 153 377 161 411
rect 109 343 161 377
rect 109 309 119 343
rect 153 309 161 343
rect 109 297 161 309
rect 215 479 267 497
rect 215 445 223 479
rect 257 445 267 479
rect 215 411 267 445
rect 215 377 223 411
rect 257 377 267 411
rect 215 343 267 377
rect 215 309 223 343
rect 257 309 267 343
rect 215 297 267 309
rect 297 485 351 497
rect 297 451 307 485
rect 341 451 351 485
rect 297 417 351 451
rect 297 383 307 417
rect 341 383 351 417
rect 297 297 351 383
rect 381 479 435 497
rect 381 445 391 479
rect 425 445 435 479
rect 381 411 435 445
rect 381 377 391 411
rect 425 377 435 411
rect 381 343 435 377
rect 381 309 391 343
rect 425 309 435 343
rect 381 297 435 309
rect 465 485 519 497
rect 465 451 475 485
rect 509 451 519 485
rect 465 417 519 451
rect 465 383 475 417
rect 509 383 519 417
rect 465 297 519 383
rect 549 479 603 497
rect 549 445 559 479
rect 593 445 603 479
rect 549 411 603 445
rect 549 377 559 411
rect 593 377 603 411
rect 549 343 603 377
rect 549 309 559 343
rect 593 309 603 343
rect 549 297 603 309
rect 633 485 687 497
rect 633 451 643 485
rect 677 451 687 485
rect 633 417 687 451
rect 633 383 643 417
rect 677 383 687 417
rect 633 297 687 383
rect 717 479 771 497
rect 717 445 727 479
rect 761 445 771 479
rect 717 411 771 445
rect 717 377 727 411
rect 761 377 771 411
rect 717 343 771 377
rect 717 309 727 343
rect 761 309 771 343
rect 717 297 771 309
rect 801 485 855 497
rect 801 451 811 485
rect 845 451 855 485
rect 801 417 855 451
rect 801 383 811 417
rect 845 383 855 417
rect 801 297 855 383
rect 885 479 939 497
rect 885 445 895 479
rect 929 445 939 479
rect 885 411 939 445
rect 885 377 895 411
rect 929 377 939 411
rect 885 343 939 377
rect 885 309 895 343
rect 929 309 939 343
rect 885 297 939 309
rect 969 485 1023 497
rect 969 451 979 485
rect 1013 451 1023 485
rect 969 417 1023 451
rect 969 383 979 417
rect 1013 383 1023 417
rect 969 297 1023 383
rect 1053 479 1107 497
rect 1053 445 1063 479
rect 1097 445 1107 479
rect 1053 411 1107 445
rect 1053 377 1063 411
rect 1097 377 1107 411
rect 1053 343 1107 377
rect 1053 309 1063 343
rect 1097 309 1107 343
rect 1053 297 1107 309
rect 1137 485 1189 497
rect 1137 451 1147 485
rect 1181 451 1189 485
rect 1137 417 1189 451
rect 1137 383 1147 417
rect 1181 383 1189 417
rect 1137 297 1189 383
<< ndiffc >>
rect 35 131 69 165
rect 35 63 69 97
rect 119 131 153 165
rect 119 63 153 97
rect 223 131 257 165
rect 223 63 257 97
rect 307 63 341 97
rect 391 131 425 165
rect 391 63 425 97
rect 475 63 509 97
rect 559 131 593 165
rect 559 63 593 97
rect 643 63 677 97
rect 727 131 761 165
rect 727 63 761 97
rect 811 63 845 97
rect 895 131 929 165
rect 895 63 929 97
rect 979 63 1013 97
rect 1063 131 1097 165
rect 1063 63 1097 97
rect 1147 63 1181 97
<< pdiffc >>
rect 35 451 69 485
rect 35 383 69 417
rect 35 315 69 349
rect 119 445 153 479
rect 119 377 153 411
rect 119 309 153 343
rect 223 445 257 479
rect 223 377 257 411
rect 223 309 257 343
rect 307 451 341 485
rect 307 383 341 417
rect 391 445 425 479
rect 391 377 425 411
rect 391 309 425 343
rect 475 451 509 485
rect 475 383 509 417
rect 559 445 593 479
rect 559 377 593 411
rect 559 309 593 343
rect 643 451 677 485
rect 643 383 677 417
rect 727 445 761 479
rect 727 377 761 411
rect 727 309 761 343
rect 811 451 845 485
rect 811 383 845 417
rect 895 445 929 479
rect 895 377 929 411
rect 895 309 929 343
rect 979 451 1013 485
rect 979 383 1013 417
rect 1063 445 1097 479
rect 1063 377 1097 411
rect 1063 309 1097 343
rect 1147 451 1181 485
rect 1147 383 1181 417
<< poly >>
rect 79 497 109 523
rect 267 497 297 523
rect 351 497 381 523
rect 435 497 465 523
rect 519 497 549 523
rect 603 497 633 523
rect 687 497 717 523
rect 771 497 801 523
rect 855 497 885 523
rect 939 497 969 523
rect 1023 497 1053 523
rect 1107 497 1137 523
rect 79 265 109 297
rect 21 249 109 265
rect 21 215 38 249
rect 72 215 109 249
rect 21 199 109 215
rect 79 177 109 199
rect 267 259 297 297
rect 351 259 381 297
rect 435 259 465 297
rect 267 249 465 259
rect 267 215 307 249
rect 341 215 375 249
rect 409 215 465 249
rect 267 205 465 215
rect 267 177 297 205
rect 351 177 381 205
rect 435 177 465 205
rect 519 259 549 297
rect 603 259 633 297
rect 687 259 717 297
rect 771 259 801 297
rect 855 259 885 297
rect 939 259 969 297
rect 1023 259 1053 297
rect 1107 259 1137 297
rect 519 249 1137 259
rect 519 215 543 249
rect 577 215 611 249
rect 645 215 679 249
rect 713 215 747 249
rect 781 215 815 249
rect 849 215 883 249
rect 917 215 951 249
rect 985 215 1019 249
rect 1053 215 1087 249
rect 1121 215 1137 249
rect 519 205 1137 215
rect 519 177 549 205
rect 603 177 633 205
rect 687 177 717 205
rect 771 177 801 205
rect 855 177 885 205
rect 939 177 969 205
rect 1023 177 1053 205
rect 1107 177 1137 205
rect 79 21 109 47
rect 267 21 297 47
rect 351 21 381 47
rect 435 21 465 47
rect 519 21 549 47
rect 603 21 633 47
rect 687 21 717 47
rect 771 21 801 47
rect 855 21 885 47
rect 939 21 969 47
rect 1023 21 1053 47
rect 1107 21 1137 47
<< polycont >>
rect 38 215 72 249
rect 307 215 341 249
rect 375 215 409 249
rect 543 215 577 249
rect 611 215 645 249
rect 679 215 713 249
rect 747 215 781 249
rect 815 215 849 249
rect 883 215 917 249
rect 951 215 985 249
rect 1019 215 1053 249
rect 1087 215 1121 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1288 561
rect 35 485 69 527
rect 35 417 69 451
rect 35 349 69 383
rect 35 289 69 315
rect 103 479 169 493
rect 103 445 119 479
rect 153 445 169 479
rect 103 411 169 445
rect 103 377 119 411
rect 153 377 169 411
rect 103 343 169 377
rect 103 309 119 343
rect 153 309 169 343
rect 135 255 169 309
rect 207 479 273 493
rect 207 445 223 479
rect 257 445 273 479
rect 207 411 273 445
rect 207 377 223 411
rect 257 377 273 411
rect 207 343 273 377
rect 307 485 341 527
rect 307 417 341 451
rect 307 357 341 383
rect 375 479 441 493
rect 375 445 391 479
rect 425 445 441 479
rect 375 411 441 445
rect 375 377 391 411
rect 425 377 441 411
rect 207 309 223 343
rect 257 323 273 343
rect 375 343 441 377
rect 475 485 509 527
rect 475 417 509 451
rect 475 357 509 383
rect 543 479 609 493
rect 543 445 559 479
rect 593 445 609 479
rect 543 411 609 445
rect 543 377 559 411
rect 593 377 609 411
rect 375 323 391 343
rect 257 309 391 323
rect 425 323 441 343
rect 543 343 609 377
rect 643 485 677 527
rect 643 417 677 451
rect 643 367 677 383
rect 711 479 777 493
rect 711 445 727 479
rect 761 445 777 479
rect 711 411 777 445
rect 711 377 727 411
rect 761 377 777 411
rect 425 309 509 323
rect 207 289 509 309
rect 543 309 559 343
rect 593 323 609 343
rect 711 343 777 377
rect 811 485 845 527
rect 811 417 845 451
rect 811 367 845 383
rect 879 479 945 493
rect 879 445 895 479
rect 929 445 945 479
rect 879 411 945 445
rect 879 377 895 411
rect 929 377 945 411
rect 711 323 727 343
rect 593 309 727 323
rect 761 323 777 343
rect 879 343 945 377
rect 979 485 1013 527
rect 979 417 1013 451
rect 979 367 1013 383
rect 1047 479 1113 493
rect 1047 445 1063 479
rect 1097 445 1113 479
rect 1047 411 1113 445
rect 1047 377 1063 411
rect 1097 377 1113 411
rect 879 323 895 343
rect 761 309 895 323
rect 929 323 945 343
rect 1047 343 1113 377
rect 1147 485 1181 527
rect 1147 417 1181 451
rect 1147 367 1181 383
rect 1047 323 1063 343
rect 929 309 1063 323
rect 1097 323 1113 343
rect 1097 309 1271 323
rect 543 289 1271 309
rect 475 255 509 289
rect 17 249 101 255
rect 17 215 38 249
rect 72 215 101 249
rect 135 249 441 255
rect 135 215 307 249
rect 341 215 375 249
rect 409 215 441 249
rect 475 249 1152 255
rect 475 215 543 249
rect 577 215 611 249
rect 645 215 679 249
rect 713 215 747 249
rect 781 215 815 249
rect 849 215 883 249
rect 917 215 951 249
rect 985 215 1019 249
rect 1053 215 1087 249
rect 1121 215 1152 249
rect 135 181 169 215
rect 475 181 509 215
rect 1194 181 1271 289
rect 35 165 69 181
rect 35 97 69 131
rect 35 17 69 63
rect 103 165 169 181
rect 103 131 119 165
rect 153 131 169 165
rect 103 97 169 131
rect 103 63 119 97
rect 153 63 169 97
rect 103 52 169 63
rect 207 165 509 181
rect 207 131 223 165
rect 257 147 391 165
rect 257 131 273 147
rect 207 97 273 131
rect 375 131 391 147
rect 425 147 509 165
rect 543 165 1271 181
rect 425 131 441 147
rect 207 63 223 97
rect 257 63 273 97
rect 207 52 273 63
rect 307 97 341 113
rect 307 17 341 63
rect 375 97 441 131
rect 543 131 559 165
rect 593 147 727 165
rect 593 131 609 147
rect 375 63 391 97
rect 425 63 441 97
rect 375 52 441 63
rect 475 97 509 113
rect 475 17 509 63
rect 543 97 609 131
rect 711 131 727 147
rect 761 147 895 165
rect 761 131 777 147
rect 543 63 559 97
rect 593 63 609 97
rect 543 52 609 63
rect 643 97 677 113
rect 643 17 677 63
rect 711 97 777 131
rect 879 131 895 147
rect 929 147 1063 165
rect 929 131 945 147
rect 711 63 727 97
rect 761 63 777 97
rect 711 52 777 63
rect 811 97 845 113
rect 811 17 845 63
rect 879 97 945 131
rect 1047 131 1063 147
rect 1097 147 1271 165
rect 1097 131 1113 147
rect 879 63 895 97
rect 929 63 945 97
rect 879 52 945 63
rect 979 97 1013 113
rect 979 17 1013 63
rect 1047 97 1113 131
rect 1047 63 1063 97
rect 1097 63 1113 97
rect 1047 52 1113 63
rect 1147 97 1181 113
rect 1147 17 1181 63
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1288 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 1225 527 1259 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
rect 1225 -17 1259 17
<< metal1 >>
rect 0 561 1288 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1288 561
rect 0 496 1288 527
rect 0 17 1288 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1288 17
rect 0 -48 1288 -17
<< labels >>
flabel locali s 30 221 64 255 0 FreeSans 200 0 0 0 A
port 1 nsew signal input
flabel locali s 1225 221 1259 255 0 FreeSans 200 0 0 0 Y
port 6 nsew signal output
flabel locali s 1225 289 1259 323 0 FreeSans 200 0 0 0 Y
port 6 nsew signal output
flabel pwell s 30 -17 64 17 0 FreeSans 200 0 0 0 VNB
port 3 nsew ground bidirectional
flabel nwell s 30 527 64 561 0 FreeSans 200 0 0 0 VPB
port 4 nsew power bidirectional
flabel metal1 s 30 -17 64 17 0 FreeSans 200 0 0 0 VGND
port 2 nsew ground bidirectional abutment
flabel metal1 s 30 527 64 561 0 FreeSans 200 0 0 0 VPWR
port 5 nsew power bidirectional abutment
rlabel comment s 0 0 0 0 4 bufinv_8
rlabel metal1 s 0 -48 1288 48 1 VGND
port 2 nsew ground bidirectional abutment
rlabel metal1 s 0 496 1288 592 1 VPWR
port 5 nsew power bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 1288 544
string GDS_END 3224762
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_START 3214610
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string path 0.000 0.000 32.200 0.000 
<< end >>
