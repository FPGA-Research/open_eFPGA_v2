magic
tech sky130A
timestamp 1707688321
<< metal1 >>
rect 0 0 3 154
rect 157 0 160 154
<< via1 >>
rect 3 0 157 154
<< metal2 >>
rect 0 0 3 154
rect 157 0 160 154
<< properties >>
string GDS_END 86913194
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 86911462
<< end >>
