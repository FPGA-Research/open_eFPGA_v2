magic
tech sky130A
timestamp 1707688321
<< metal1 >>
rect 0 0 3 90
rect 221 0 224 90
<< via1 >>
rect 3 0 221 90
<< metal2 >>
rect 0 0 3 90
rect 221 0 224 90
<< properties >>
string GDS_END 86905458
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 86903982
<< end >>
