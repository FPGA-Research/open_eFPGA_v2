magic
tech sky130B
magscale 1 2
timestamp 1707688321
use sky130_fd_pr__dfl1sd2__example_55959141808521  sky130_fd_pr__dfl1sd2__example_55959141808521_0
timestamp 1707688321
transform 1 0 100 0 1 0
box 0 0 1 1
use sky130_fd_pr__dfl1sd2__example_55959141808521  sky130_fd_pr__dfl1sd2__example_55959141808521_1
timestamp 1707688321
transform 1 0 256 0 1 0
box 0 0 1 1
use sky130_fd_pr__dfl1sd2__example_55959141808521  sky130_fd_pr__dfl1sd2__example_55959141808521_2
timestamp 1707688321
transform 1 0 412 0 1 0
box 0 0 1 1
use sky130_fd_pr__dfl1sd2__example_55959141808521  sky130_fd_pr__dfl1sd2__example_55959141808521_3
timestamp 1707688321
transform 1 0 568 0 1 0
box 0 0 1 1
use sky130_fd_pr__dfl1sd__example_55959141808520  sky130_fd_pr__dfl1sd__example_55959141808520_0
timestamp 1707688321
transform -1 0 0 0 1 0
box 0 0 1 1
use sky130_fd_pr__dfl1sd__example_55959141808520  sky130_fd_pr__dfl1sd__example_55959141808520_1
timestamp 1707688321
transform 1 0 724 0 1 0
box 0 0 1 1
<< properties >>
string GDS_END 63732174
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 63729188
<< end >>
