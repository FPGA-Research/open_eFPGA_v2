magic
tech sky130B
magscale 1 2
timestamp 1707688321
<< pwell >>
rect 1176 1289 1197 1338
<< obsli1 >>
rect 0 2272 2282 2338
rect 0 2166 66 2272
rect 100 2202 2181 2236
rect 0 2132 1080 2166
rect 0 2026 66 2132
rect 1114 2096 1168 2202
rect 2216 2166 2282 2272
rect 1202 2132 2282 2166
rect 100 2062 2181 2096
rect 0 1992 1080 2026
rect 0 1886 66 1992
rect 1114 1956 1168 2062
rect 2216 2026 2282 2132
rect 1202 1992 2282 2026
rect 100 1922 2181 1956
rect 0 1852 1080 1886
rect 0 1746 66 1852
rect 1114 1816 1168 1922
rect 2216 1886 2282 1992
rect 1202 1852 2282 1886
rect 100 1782 2181 1816
rect 0 1712 1080 1746
rect 0 1606 66 1712
rect 1114 1676 1168 1782
rect 2216 1746 2282 1852
rect 1202 1712 2282 1746
rect 100 1642 2181 1676
rect 0 1572 1080 1606
rect 0 1466 66 1572
rect 1114 1536 1168 1642
rect 2216 1606 2282 1712
rect 1202 1572 2282 1606
rect 100 1502 2181 1536
rect 0 1432 1080 1466
rect 0 1326 66 1432
rect 1114 1396 1168 1502
rect 2216 1466 2282 1572
rect 1202 1432 2282 1466
rect 100 1362 2181 1396
rect 0 1292 1080 1326
rect 0 1186 66 1292
rect 1114 1256 1168 1362
rect 2216 1326 2282 1432
rect 1202 1292 2282 1326
rect 100 1222 2181 1256
rect 0 1152 1080 1186
rect 0 1046 66 1152
rect 1114 1116 1168 1222
rect 2216 1186 2282 1292
rect 1202 1152 2282 1186
rect 100 1082 2181 1116
rect 0 1012 1080 1046
rect 0 906 66 1012
rect 1114 976 1168 1082
rect 2216 1046 2282 1152
rect 1202 1012 2282 1046
rect 100 942 2181 976
rect 0 872 1080 906
rect 0 766 66 872
rect 1114 836 1168 942
rect 2216 906 2282 1012
rect 1202 872 2282 906
rect 100 802 2181 836
rect 0 732 1080 766
rect 0 626 66 732
rect 1114 696 1168 802
rect 2216 766 2282 872
rect 1202 732 2282 766
rect 100 662 2181 696
rect 0 592 1080 626
rect 0 486 66 592
rect 1114 556 1168 662
rect 2216 626 2282 732
rect 1202 592 2282 626
rect 100 522 2181 556
rect 0 452 1080 486
rect 0 346 66 452
rect 1114 416 1168 522
rect 2216 486 2282 592
rect 1202 452 2282 486
rect 100 382 2181 416
rect 0 312 1080 346
rect 0 206 66 312
rect 1114 276 1168 382
rect 2216 346 2282 452
rect 1202 312 2282 346
rect 100 242 2181 276
rect 0 172 1080 206
rect 0 66 66 172
rect 1114 136 1168 242
rect 2216 206 2282 312
rect 1202 172 2282 206
rect 100 102 2181 136
rect 2216 66 2282 172
rect 0 0 2282 66
<< obsm1 >>
rect 0 2272 2282 2338
rect 0 66 66 2272
rect 100 1201 128 2244
rect 156 1229 184 2272
rect 212 1201 240 2244
rect 268 1229 296 2272
rect 324 1201 352 2244
rect 380 1229 408 2272
rect 436 1201 464 2244
rect 492 1229 520 2272
rect 548 1201 576 2244
rect 604 1229 632 2272
rect 660 1201 688 2244
rect 716 1229 744 2272
rect 772 1201 800 2244
rect 828 1229 856 2272
rect 884 1201 912 2244
rect 940 1229 968 2272
rect 996 1201 1024 2244
rect 1052 1229 1080 2272
rect 1114 1201 1168 2244
rect 1202 1229 1230 2272
rect 1258 1201 1286 2244
rect 1314 1229 1342 2272
rect 1370 1201 1398 2244
rect 1426 1229 1454 2272
rect 1482 1201 1510 2244
rect 1538 1229 1566 2272
rect 1594 1201 1622 2244
rect 1650 1229 1678 2272
rect 1706 1201 1734 2244
rect 1762 1229 1790 2272
rect 1818 1201 1846 2244
rect 1874 1229 1902 2272
rect 1930 1201 1958 2244
rect 1986 1229 2014 2272
rect 2042 1201 2070 2244
rect 2098 1229 2126 2272
rect 2154 1201 2182 2244
rect 100 1137 2182 1201
rect 100 94 128 1137
rect 156 66 184 1109
rect 212 94 240 1137
rect 268 66 296 1109
rect 324 94 352 1137
rect 380 66 408 1109
rect 436 94 464 1137
rect 492 66 520 1109
rect 548 94 576 1137
rect 604 66 632 1109
rect 660 94 688 1137
rect 716 66 744 1109
rect 772 94 800 1137
rect 828 66 856 1109
rect 884 94 912 1137
rect 940 66 968 1109
rect 996 94 1024 1137
rect 1052 66 1080 1109
rect 1114 94 1168 1137
rect 1202 66 1230 1109
rect 1258 94 1286 1137
rect 1314 66 1342 1109
rect 1370 94 1398 1137
rect 1426 66 1454 1109
rect 1482 94 1510 1137
rect 1538 66 1566 1109
rect 1594 94 1622 1137
rect 1650 66 1678 1109
rect 1706 94 1734 1137
rect 1762 66 1790 1109
rect 1818 94 1846 1137
rect 1874 66 1902 1109
rect 1930 94 1958 1137
rect 1986 66 2014 1109
rect 2042 94 2070 1137
rect 2098 66 2126 1109
rect 2154 94 2182 1137
rect 2216 66 2282 2272
rect 0 0 2282 66
<< metal2 >>
rect 0 2272 1086 2338
rect 0 2188 66 2272
rect 1114 2244 1168 2338
rect 1196 2272 2282 2338
rect 94 2216 2188 2244
rect 0 2160 1086 2188
rect 0 2076 66 2160
rect 1114 2132 1168 2216
rect 2216 2188 2282 2272
rect 1196 2160 2282 2188
rect 94 2104 2188 2132
rect 0 2048 1086 2076
rect 0 1964 66 2048
rect 1114 2020 1168 2104
rect 2216 2076 2282 2160
rect 1196 2048 2282 2076
rect 94 1992 2188 2020
rect 0 1936 1086 1964
rect 0 1852 66 1936
rect 1114 1908 1168 1992
rect 2216 1964 2282 2048
rect 1196 1936 2282 1964
rect 94 1880 2188 1908
rect 0 1824 1086 1852
rect 0 1740 66 1824
rect 1114 1796 1168 1880
rect 2216 1852 2282 1936
rect 1196 1824 2282 1852
rect 94 1768 2188 1796
rect 0 1712 1086 1740
rect 0 1628 66 1712
rect 1114 1684 1168 1768
rect 2216 1740 2282 1824
rect 1196 1712 2282 1740
rect 94 1656 2188 1684
rect 0 1600 1086 1628
rect 0 1516 66 1600
rect 1114 1572 1168 1656
rect 2216 1628 2282 1712
rect 1196 1600 2282 1628
rect 94 1544 2188 1572
rect 0 1488 1086 1516
rect 0 1404 66 1488
rect 1114 1460 1168 1544
rect 2216 1516 2282 1600
rect 1196 1488 2282 1516
rect 94 1432 2188 1460
rect 0 1376 1086 1404
rect 0 1292 66 1376
rect 1114 1348 1168 1432
rect 2216 1404 2282 1488
rect 1196 1376 2282 1404
rect 94 1320 2188 1348
rect 0 1264 1086 1292
rect 0 1224 66 1264
rect 1114 1196 1168 1320
rect 2216 1292 2282 1376
rect 1196 1264 2282 1292
rect 2216 1224 2282 1264
rect 0 1142 2282 1196
rect 0 1074 66 1114
rect 0 1046 1086 1074
rect 0 962 66 1046
rect 1114 1018 1168 1142
rect 2216 1074 2282 1114
rect 1196 1046 2282 1074
rect 94 990 2188 1018
rect 0 934 1086 962
rect 0 850 66 934
rect 1114 906 1168 990
rect 2216 962 2282 1046
rect 1196 934 2282 962
rect 94 878 2188 906
rect 0 822 1086 850
rect 0 738 66 822
rect 1114 794 1168 878
rect 2216 850 2282 934
rect 1196 822 2282 850
rect 94 766 2188 794
rect 0 710 1086 738
rect 0 626 66 710
rect 1114 682 1168 766
rect 2216 738 2282 822
rect 1196 710 2282 738
rect 94 654 2188 682
rect 0 598 1086 626
rect 0 514 66 598
rect 1114 570 1168 654
rect 2216 626 2282 710
rect 1196 598 2282 626
rect 94 542 2188 570
rect 0 486 1086 514
rect 0 402 66 486
rect 1114 458 1168 542
rect 2216 514 2282 598
rect 1196 486 2282 514
rect 94 430 2188 458
rect 0 374 1086 402
rect 0 290 66 374
rect 1114 346 1168 430
rect 2216 402 2282 486
rect 1196 374 2282 402
rect 94 318 2188 346
rect 0 262 1086 290
rect 0 178 66 262
rect 1114 234 1168 318
rect 2216 290 2282 374
rect 1196 262 2282 290
rect 94 206 2188 234
rect 0 150 1086 178
rect 0 66 66 150
rect 1114 122 1168 206
rect 2216 178 2282 262
rect 1196 150 2282 178
rect 94 94 2188 122
rect 0 0 1086 66
rect 1114 0 1168 94
rect 2216 66 2282 150
rect 1196 0 2282 66
<< metal3 >>
rect 0 0 2282 2338
<< labels >>
rlabel metal2 s 2216 2188 2282 2272 6 C0
port 1 nsew
rlabel metal2 s 2216 2076 2282 2160 6 C0
port 1 nsew
rlabel metal2 s 2216 1964 2282 2048 6 C0
port 1 nsew
rlabel metal2 s 2216 1852 2282 1936 6 C0
port 1 nsew
rlabel metal2 s 2216 1740 2282 1824 6 C0
port 1 nsew
rlabel metal2 s 2216 1628 2282 1712 6 C0
port 1 nsew
rlabel metal2 s 2216 1516 2282 1600 6 C0
port 1 nsew
rlabel metal2 s 2216 1404 2282 1488 6 C0
port 1 nsew
rlabel metal2 s 2216 1292 2282 1376 6 C0
port 1 nsew
rlabel metal2 s 2216 1224 2282 1264 6 C0
port 1 nsew
rlabel metal2 s 2216 1074 2282 1114 6 C0
port 1 nsew
rlabel metal2 s 2216 962 2282 1046 6 C0
port 1 nsew
rlabel metal2 s 2216 850 2282 934 6 C0
port 1 nsew
rlabel metal2 s 2216 738 2282 822 6 C0
port 1 nsew
rlabel metal2 s 2216 626 2282 710 6 C0
port 1 nsew
rlabel metal2 s 2216 514 2282 598 6 C0
port 1 nsew
rlabel metal2 s 2216 402 2282 486 6 C0
port 1 nsew
rlabel metal2 s 2216 290 2282 374 6 C0
port 1 nsew
rlabel metal2 s 2216 178 2282 262 6 C0
port 1 nsew
rlabel metal2 s 2216 66 2282 150 6 C0
port 1 nsew
rlabel metal2 s 1196 2272 2282 2338 6 C0
port 1 nsew
rlabel metal2 s 1196 2160 2282 2188 6 C0
port 1 nsew
rlabel metal2 s 1196 2048 2282 2076 6 C0
port 1 nsew
rlabel metal2 s 1196 1936 2282 1964 6 C0
port 1 nsew
rlabel metal2 s 1196 1824 2282 1852 6 C0
port 1 nsew
rlabel metal2 s 1196 1712 2282 1740 6 C0
port 1 nsew
rlabel metal2 s 1196 1600 2282 1628 6 C0
port 1 nsew
rlabel metal2 s 1196 1488 2282 1516 6 C0
port 1 nsew
rlabel metal2 s 1196 1376 2282 1404 6 C0
port 1 nsew
rlabel metal2 s 1196 1264 2282 1292 6 C0
port 1 nsew
rlabel metal2 s 1196 1046 2282 1074 6 C0
port 1 nsew
rlabel metal2 s 1196 934 2282 962 6 C0
port 1 nsew
rlabel metal2 s 1196 822 2282 850 6 C0
port 1 nsew
rlabel metal2 s 1196 710 2282 738 6 C0
port 1 nsew
rlabel metal2 s 1196 598 2282 626 6 C0
port 1 nsew
rlabel metal2 s 1196 486 2282 514 6 C0
port 1 nsew
rlabel metal2 s 1196 374 2282 402 6 C0
port 1 nsew
rlabel metal2 s 1196 262 2282 290 6 C0
port 1 nsew
rlabel metal2 s 1196 150 2282 178 6 C0
port 1 nsew
rlabel metal2 s 1196 0 2282 66 6 C0
port 1 nsew
rlabel metal2 s 0 2272 1086 2338 6 C0
port 1 nsew
rlabel metal2 s 0 2188 66 2272 6 C0
port 1 nsew
rlabel metal2 s 0 2160 1086 2188 6 C0
port 1 nsew
rlabel metal2 s 0 2076 66 2160 6 C0
port 1 nsew
rlabel metal2 s 0 2048 1086 2076 6 C0
port 1 nsew
rlabel metal2 s 0 1964 66 2048 6 C0
port 1 nsew
rlabel metal2 s 0 1936 1086 1964 6 C0
port 1 nsew
rlabel metal2 s 0 1852 66 1936 6 C0
port 1 nsew
rlabel metal2 s 0 1824 1086 1852 6 C0
port 1 nsew
rlabel metal2 s 0 1740 66 1824 6 C0
port 1 nsew
rlabel metal2 s 0 1712 1086 1740 6 C0
port 1 nsew
rlabel metal2 s 0 1628 66 1712 6 C0
port 1 nsew
rlabel metal2 s 0 1600 1086 1628 6 C0
port 1 nsew
rlabel metal2 s 0 1516 66 1600 6 C0
port 1 nsew
rlabel metal2 s 0 1488 1086 1516 6 C0
port 1 nsew
rlabel metal2 s 0 1404 66 1488 6 C0
port 1 nsew
rlabel metal2 s 0 1376 1086 1404 6 C0
port 1 nsew
rlabel metal2 s 0 1292 66 1376 6 C0
port 1 nsew
rlabel metal2 s 0 1264 1086 1292 6 C0
port 1 nsew
rlabel metal2 s 0 1224 66 1264 6 C0
port 1 nsew
rlabel metal2 s 0 1074 66 1114 6 C0
port 1 nsew
rlabel metal2 s 0 1046 1086 1074 6 C0
port 1 nsew
rlabel metal2 s 0 962 66 1046 6 C0
port 1 nsew
rlabel metal2 s 0 934 1086 962 6 C0
port 1 nsew
rlabel metal2 s 0 850 66 934 6 C0
port 1 nsew
rlabel metal2 s 0 822 1086 850 6 C0
port 1 nsew
rlabel metal2 s 0 738 66 822 6 C0
port 1 nsew
rlabel metal2 s 0 710 1086 738 6 C0
port 1 nsew
rlabel metal2 s 0 626 66 710 6 C0
port 1 nsew
rlabel metal2 s 0 598 1086 626 6 C0
port 1 nsew
rlabel metal2 s 0 514 66 598 6 C0
port 1 nsew
rlabel metal2 s 0 486 1086 514 6 C0
port 1 nsew
rlabel metal2 s 0 402 66 486 6 C0
port 1 nsew
rlabel metal2 s 0 374 1086 402 6 C0
port 1 nsew
rlabel metal2 s 0 290 66 374 6 C0
port 1 nsew
rlabel metal2 s 0 262 1086 290 6 C0
port 1 nsew
rlabel metal2 s 0 178 66 262 6 C0
port 1 nsew
rlabel metal2 s 0 150 1086 178 6 C0
port 1 nsew
rlabel metal2 s 0 66 66 150 6 C0
port 1 nsew
rlabel metal2 s 0 0 1086 66 6 C0
port 1 nsew
rlabel metal2 s 1114 2244 1168 2338 6 C1
port 2 nsew
rlabel metal2 s 1114 2132 1168 2216 6 C1
port 2 nsew
rlabel metal2 s 1114 2020 1168 2104 6 C1
port 2 nsew
rlabel metal2 s 1114 1908 1168 1992 6 C1
port 2 nsew
rlabel metal2 s 1114 1796 1168 1880 6 C1
port 2 nsew
rlabel metal2 s 1114 1684 1168 1768 6 C1
port 2 nsew
rlabel metal2 s 1114 1572 1168 1656 6 C1
port 2 nsew
rlabel metal2 s 1114 1460 1168 1544 6 C1
port 2 nsew
rlabel metal2 s 1114 1348 1168 1432 6 C1
port 2 nsew
rlabel metal2 s 1114 1196 1168 1320 6 C1
port 2 nsew
rlabel metal2 s 1114 1018 1168 1142 6 C1
port 2 nsew
rlabel metal2 s 1114 906 1168 990 6 C1
port 2 nsew
rlabel metal2 s 1114 794 1168 878 6 C1
port 2 nsew
rlabel metal2 s 1114 682 1168 766 6 C1
port 2 nsew
rlabel metal2 s 1114 570 1168 654 6 C1
port 2 nsew
rlabel metal2 s 1114 458 1168 542 6 C1
port 2 nsew
rlabel metal2 s 1114 346 1168 430 6 C1
port 2 nsew
rlabel metal2 s 1114 234 1168 318 6 C1
port 2 nsew
rlabel metal2 s 1114 122 1168 206 6 C1
port 2 nsew
rlabel metal2 s 1114 0 1168 94 6 C1
port 2 nsew
rlabel metal2 s 94 2216 2188 2244 6 C1
port 2 nsew
rlabel metal2 s 94 2104 2188 2132 6 C1
port 2 nsew
rlabel metal2 s 94 1992 2188 2020 6 C1
port 2 nsew
rlabel metal2 s 94 1880 2188 1908 6 C1
port 2 nsew
rlabel metal2 s 94 1768 2188 1796 6 C1
port 2 nsew
rlabel metal2 s 94 1656 2188 1684 6 C1
port 2 nsew
rlabel metal2 s 94 1544 2188 1572 6 C1
port 2 nsew
rlabel metal2 s 94 1432 2188 1460 6 C1
port 2 nsew
rlabel metal2 s 94 1320 2188 1348 6 C1
port 2 nsew
rlabel metal2 s 94 990 2188 1018 6 C1
port 2 nsew
rlabel metal2 s 94 878 2188 906 6 C1
port 2 nsew
rlabel metal2 s 94 766 2188 794 6 C1
port 2 nsew
rlabel metal2 s 94 654 2188 682 6 C1
port 2 nsew
rlabel metal2 s 94 542 2188 570 6 C1
port 2 nsew
rlabel metal2 s 94 430 2188 458 6 C1
port 2 nsew
rlabel metal2 s 94 318 2188 346 6 C1
port 2 nsew
rlabel metal2 s 94 206 2188 234 6 C1
port 2 nsew
rlabel metal2 s 94 94 2188 122 6 C1
port 2 nsew
rlabel metal2 s 0 1142 2282 1196 6 C1
port 2 nsew
rlabel metal3 s 0 0 2282 2338 6 MET3
port 4 nsew
rlabel pwell s 1176 1289 1197 1338 6 SUB
port 3 nsew
<< properties >>
string FIXED_BBOX 0 0 2282 2338
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 678284
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_pr/gds/sky130_fd_pr.gds
string GDS_START 627998
string device primitive
<< end >>
