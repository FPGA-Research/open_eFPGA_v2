magic
tech sky130B
magscale 1 2
timestamp 1707688321
<< dnwell >>
rect 147 7540 2857 8764
rect 26 34 2857 7540
<< nwell >>
rect -59 7249 2937 7419
rect -59 2201 111 7249
rect 2577 2201 2937 7249
rect -59 2031 2937 2201
rect -59 -9 111 2031
rect 694 1504 1994 2031
rect 2577 -46 2937 2031
<< pwell >>
rect 29 7479 2706 7567
rect 171 7079 2517 7167
rect 171 2349 259 7079
rect 2429 2349 2517 7079
rect 171 2261 2517 2349
<< mvpsubdiff >>
rect 55 7540 2680 7541
rect 55 7506 89 7540
rect 123 7506 157 7540
rect 191 7506 225 7540
rect 259 7506 293 7540
rect 327 7506 361 7540
rect 395 7506 429 7540
rect 463 7506 497 7540
rect 531 7506 565 7540
rect 599 7506 633 7540
rect 667 7506 701 7540
rect 735 7506 769 7540
rect 803 7506 837 7540
rect 871 7506 905 7540
rect 939 7506 973 7540
rect 1007 7506 1041 7540
rect 1075 7506 1109 7540
rect 1143 7506 1177 7540
rect 1211 7506 1245 7540
rect 1279 7506 1313 7540
rect 1347 7506 1381 7540
rect 1415 7506 1449 7540
rect 1483 7506 1517 7540
rect 1551 7506 1585 7540
rect 1619 7506 1653 7540
rect 1687 7506 1721 7540
rect 1755 7506 1789 7540
rect 1823 7506 1857 7540
rect 1891 7506 1925 7540
rect 1959 7506 1993 7540
rect 2027 7506 2061 7540
rect 2095 7506 2129 7540
rect 2163 7506 2197 7540
rect 2231 7506 2265 7540
rect 2299 7506 2333 7540
rect 2367 7506 2401 7540
rect 2435 7506 2469 7540
rect 2503 7506 2537 7540
rect 2571 7506 2605 7540
rect 2639 7506 2680 7540
rect 55 7505 2680 7506
rect 197 7140 2491 7141
rect 197 7106 231 7140
rect 265 7106 299 7140
rect 333 7106 367 7140
rect 401 7106 435 7140
rect 469 7106 503 7140
rect 537 7106 571 7140
rect 605 7106 639 7140
rect 673 7106 707 7140
rect 741 7106 775 7140
rect 809 7106 843 7140
rect 877 7106 911 7140
rect 945 7106 979 7140
rect 1013 7106 1047 7140
rect 1081 7106 1115 7140
rect 1149 7106 1183 7140
rect 1217 7106 1251 7140
rect 1285 7106 1319 7140
rect 1353 7106 1387 7140
rect 1421 7106 1455 7140
rect 1489 7106 1523 7140
rect 1557 7106 1591 7140
rect 1625 7106 1659 7140
rect 1693 7106 1727 7140
rect 1761 7106 1795 7140
rect 1829 7106 1863 7140
rect 1897 7106 1931 7140
rect 1965 7106 1999 7140
rect 2033 7106 2067 7140
rect 2101 7106 2135 7140
rect 2169 7106 2203 7140
rect 2237 7106 2271 7140
rect 2305 7106 2339 7140
rect 2373 7107 2491 7140
rect 2373 7106 2456 7107
rect 197 7105 2456 7106
rect 197 7047 233 7105
rect 2455 7073 2456 7105
rect 2490 7073 2491 7107
rect 197 7013 198 7047
rect 232 7013 233 7047
rect 197 6979 233 7013
rect 2455 7039 2491 7073
rect 2455 7005 2456 7039
rect 2490 7005 2491 7039
rect 197 6945 198 6979
rect 232 6945 233 6979
rect 197 6911 233 6945
rect 197 6877 198 6911
rect 232 6877 233 6911
rect 197 6843 233 6877
rect 197 6809 198 6843
rect 232 6809 233 6843
rect 197 6775 233 6809
rect 197 6741 198 6775
rect 232 6741 233 6775
rect 197 6707 233 6741
rect 197 6673 198 6707
rect 232 6673 233 6707
rect 197 6639 233 6673
rect 197 6605 198 6639
rect 232 6605 233 6639
rect 197 6571 233 6605
rect 197 6537 198 6571
rect 232 6537 233 6571
rect 197 6503 233 6537
rect 197 6469 198 6503
rect 232 6469 233 6503
rect 197 6435 233 6469
rect 197 6401 198 6435
rect 232 6401 233 6435
rect 197 6367 233 6401
rect 197 6333 198 6367
rect 232 6333 233 6367
rect 197 6299 233 6333
rect 197 6265 198 6299
rect 232 6265 233 6299
rect 197 6231 233 6265
rect 197 6197 198 6231
rect 232 6197 233 6231
rect 197 6163 233 6197
rect 197 6129 198 6163
rect 232 6129 233 6163
rect 197 6095 233 6129
rect 197 6061 198 6095
rect 232 6061 233 6095
rect 197 6027 233 6061
rect 197 5993 198 6027
rect 232 5993 233 6027
rect 197 5959 233 5993
rect 197 5925 198 5959
rect 232 5925 233 5959
rect 197 5891 233 5925
rect 2455 6971 2491 7005
rect 2455 6937 2456 6971
rect 2490 6937 2491 6971
rect 2455 6903 2491 6937
rect 2455 6869 2456 6903
rect 2490 6869 2491 6903
rect 2455 6835 2491 6869
rect 2455 6801 2456 6835
rect 2490 6801 2491 6835
rect 2455 6767 2491 6801
rect 2455 6733 2456 6767
rect 2490 6733 2491 6767
rect 2455 6699 2491 6733
rect 2455 6665 2456 6699
rect 2490 6665 2491 6699
rect 2455 6631 2491 6665
rect 2455 6597 2456 6631
rect 2490 6597 2491 6631
rect 2455 6563 2491 6597
rect 2455 6529 2456 6563
rect 2490 6529 2491 6563
rect 2455 6495 2491 6529
rect 2455 6461 2456 6495
rect 2490 6461 2491 6495
rect 2455 6427 2491 6461
rect 2455 6393 2456 6427
rect 2490 6393 2491 6427
rect 2455 6359 2491 6393
rect 2455 6325 2456 6359
rect 2490 6325 2491 6359
rect 2455 6291 2491 6325
rect 2455 6257 2456 6291
rect 2490 6257 2491 6291
rect 2455 6223 2491 6257
rect 2455 6189 2456 6223
rect 2490 6189 2491 6223
rect 2455 6155 2491 6189
rect 2455 6121 2456 6155
rect 2490 6121 2491 6155
rect 2455 6087 2491 6121
rect 2455 6053 2456 6087
rect 2490 6053 2491 6087
rect 2455 6019 2491 6053
rect 2455 5985 2456 6019
rect 2490 5985 2491 6019
rect 2455 5951 2491 5985
rect 197 5857 198 5891
rect 232 5857 233 5891
rect 2455 5917 2456 5951
rect 2490 5917 2491 5951
rect 2455 5883 2491 5917
rect 197 5823 233 5857
rect 197 5789 198 5823
rect 232 5789 233 5823
rect 2455 5849 2456 5883
rect 2490 5849 2491 5883
rect 2455 5815 2491 5849
rect 197 5755 233 5789
rect 197 5721 198 5755
rect 232 5721 233 5755
rect 197 5687 233 5721
rect 197 5653 198 5687
rect 232 5653 233 5687
rect 197 5619 233 5653
rect 197 5585 198 5619
rect 232 5585 233 5619
rect 197 5551 233 5585
rect 197 5517 198 5551
rect 232 5517 233 5551
rect 197 5483 233 5517
rect 197 5449 198 5483
rect 232 5449 233 5483
rect 197 5415 233 5449
rect 197 5381 198 5415
rect 232 5381 233 5415
rect 197 5347 233 5381
rect 197 5313 198 5347
rect 232 5313 233 5347
rect 197 5279 233 5313
rect 197 5245 198 5279
rect 232 5245 233 5279
rect 197 5211 233 5245
rect 197 5177 198 5211
rect 232 5177 233 5211
rect 197 5143 233 5177
rect 197 5109 198 5143
rect 232 5109 233 5143
rect 197 5075 233 5109
rect 197 5041 198 5075
rect 232 5041 233 5075
rect 197 5007 233 5041
rect 197 4973 198 5007
rect 232 4973 233 5007
rect 197 4939 233 4973
rect 197 4905 198 4939
rect 232 4905 233 4939
rect 197 4871 233 4905
rect 197 4837 198 4871
rect 232 4837 233 4871
rect 197 4803 233 4837
rect 197 4769 198 4803
rect 232 4769 233 4803
rect 197 4735 233 4769
rect 197 4701 198 4735
rect 232 4701 233 4735
rect 2455 5781 2456 5815
rect 2490 5781 2491 5815
rect 2455 5747 2491 5781
rect 2455 5713 2456 5747
rect 2490 5713 2491 5747
rect 2455 5679 2491 5713
rect 2455 5645 2456 5679
rect 2490 5645 2491 5679
rect 2455 5611 2491 5645
rect 2455 5577 2456 5611
rect 2490 5577 2491 5611
rect 2455 5543 2491 5577
rect 2455 5509 2456 5543
rect 2490 5509 2491 5543
rect 2455 5475 2491 5509
rect 2455 5441 2456 5475
rect 2490 5441 2491 5475
rect 2455 5407 2491 5441
rect 2455 5373 2456 5407
rect 2490 5373 2491 5407
rect 2455 5339 2491 5373
rect 2455 5305 2456 5339
rect 2490 5305 2491 5339
rect 2455 5271 2491 5305
rect 2455 5237 2456 5271
rect 2490 5237 2491 5271
rect 2455 5203 2491 5237
rect 2455 5169 2456 5203
rect 2490 5169 2491 5203
rect 2455 5135 2491 5169
rect 2455 5101 2456 5135
rect 2490 5101 2491 5135
rect 2455 5067 2491 5101
rect 2455 5033 2456 5067
rect 2490 5033 2491 5067
rect 2455 4999 2491 5033
rect 2455 4965 2456 4999
rect 2490 4965 2491 4999
rect 2455 4931 2491 4965
rect 2455 4897 2456 4931
rect 2490 4897 2491 4931
rect 2455 4863 2491 4897
rect 2455 4829 2456 4863
rect 2490 4829 2491 4863
rect 2455 4795 2491 4829
rect 2455 4761 2456 4795
rect 2490 4761 2491 4795
rect 197 4667 233 4701
rect 2455 4727 2491 4761
rect 2455 4693 2456 4727
rect 2490 4693 2491 4727
rect 197 4633 198 4667
rect 232 4633 233 4667
rect 197 4599 233 4633
rect 2455 4659 2491 4693
rect 2455 4625 2456 4659
rect 2490 4625 2491 4659
rect 197 4565 198 4599
rect 232 4565 233 4599
rect 197 4531 233 4565
rect 197 4497 198 4531
rect 232 4497 233 4531
rect 197 4463 233 4497
rect 197 4429 198 4463
rect 232 4429 233 4463
rect 197 4395 233 4429
rect 197 4361 198 4395
rect 232 4361 233 4395
rect 197 4327 233 4361
rect 197 4293 198 4327
rect 232 4293 233 4327
rect 197 4259 233 4293
rect 197 4225 198 4259
rect 232 4225 233 4259
rect 197 4191 233 4225
rect 197 4157 198 4191
rect 232 4157 233 4191
rect 197 4123 233 4157
rect 197 4089 198 4123
rect 232 4089 233 4123
rect 197 4055 233 4089
rect 197 4021 198 4055
rect 232 4021 233 4055
rect 197 3987 233 4021
rect 197 3953 198 3987
rect 232 3953 233 3987
rect 197 3919 233 3953
rect 197 3885 198 3919
rect 232 3885 233 3919
rect 197 3851 233 3885
rect 197 3817 198 3851
rect 232 3817 233 3851
rect 197 3783 233 3817
rect 197 3749 198 3783
rect 232 3749 233 3783
rect 197 3715 233 3749
rect 197 3681 198 3715
rect 232 3681 233 3715
rect 197 3647 233 3681
rect 197 3613 198 3647
rect 232 3613 233 3647
rect 197 3579 233 3613
rect 197 3545 198 3579
rect 232 3545 233 3579
rect 197 3511 233 3545
rect 2455 4591 2491 4625
rect 2455 4557 2456 4591
rect 2490 4557 2491 4591
rect 2455 4523 2491 4557
rect 2455 4489 2456 4523
rect 2490 4489 2491 4523
rect 2455 4455 2491 4489
rect 2455 4421 2456 4455
rect 2490 4421 2491 4455
rect 2455 4387 2491 4421
rect 2455 4353 2456 4387
rect 2490 4353 2491 4387
rect 2455 4319 2491 4353
rect 2455 4285 2456 4319
rect 2490 4285 2491 4319
rect 2455 4251 2491 4285
rect 2455 4217 2456 4251
rect 2490 4217 2491 4251
rect 2455 4183 2491 4217
rect 2455 4149 2456 4183
rect 2490 4149 2491 4183
rect 2455 4115 2491 4149
rect 2455 4081 2456 4115
rect 2490 4081 2491 4115
rect 2455 4047 2491 4081
rect 2455 4013 2456 4047
rect 2490 4013 2491 4047
rect 2455 3979 2491 4013
rect 2455 3945 2456 3979
rect 2490 3945 2491 3979
rect 2455 3911 2491 3945
rect 2455 3877 2456 3911
rect 2490 3877 2491 3911
rect 2455 3843 2491 3877
rect 2455 3809 2456 3843
rect 2490 3809 2491 3843
rect 2455 3775 2491 3809
rect 2455 3741 2456 3775
rect 2490 3741 2491 3775
rect 2455 3707 2491 3741
rect 2455 3673 2456 3707
rect 2490 3673 2491 3707
rect 2455 3639 2491 3673
rect 2455 3605 2456 3639
rect 2490 3605 2491 3639
rect 2455 3571 2491 3605
rect 2455 3537 2456 3571
rect 2490 3537 2491 3571
rect 197 3477 198 3511
rect 232 3477 233 3511
rect 2455 3503 2491 3537
rect 197 3443 233 3477
rect 197 3409 198 3443
rect 232 3409 233 3443
rect 2455 3469 2456 3503
rect 2490 3469 2491 3503
rect 2455 3435 2491 3469
rect 197 3375 233 3409
rect 197 3341 198 3375
rect 232 3341 233 3375
rect 197 3307 233 3341
rect 197 3273 198 3307
rect 232 3273 233 3307
rect 197 3239 233 3273
rect 197 3205 198 3239
rect 232 3205 233 3239
rect 197 3171 233 3205
rect 197 3137 198 3171
rect 232 3137 233 3171
rect 197 3103 233 3137
rect 197 3069 198 3103
rect 232 3069 233 3103
rect 197 3035 233 3069
rect 197 3001 198 3035
rect 232 3001 233 3035
rect 197 2967 233 3001
rect 197 2933 198 2967
rect 232 2933 233 2967
rect 197 2899 233 2933
rect 197 2865 198 2899
rect 232 2865 233 2899
rect 197 2831 233 2865
rect 197 2797 198 2831
rect 232 2797 233 2831
rect 197 2763 233 2797
rect 197 2729 198 2763
rect 232 2729 233 2763
rect 197 2695 233 2729
rect 197 2661 198 2695
rect 232 2661 233 2695
rect 197 2627 233 2661
rect 197 2593 198 2627
rect 232 2593 233 2627
rect 197 2559 233 2593
rect 197 2525 198 2559
rect 232 2525 233 2559
rect 197 2491 233 2525
rect 197 2457 198 2491
rect 232 2457 233 2491
rect 197 2423 233 2457
rect 197 2389 198 2423
rect 232 2389 233 2423
rect 197 2355 233 2389
rect 197 2321 198 2355
rect 232 2323 233 2355
rect 2455 3401 2456 3435
rect 2490 3401 2491 3435
rect 2455 3367 2491 3401
rect 2455 3333 2456 3367
rect 2490 3333 2491 3367
rect 2455 3299 2491 3333
rect 2455 3265 2456 3299
rect 2490 3265 2491 3299
rect 2455 3231 2491 3265
rect 2455 3197 2456 3231
rect 2490 3197 2491 3231
rect 2455 3163 2491 3197
rect 2455 3129 2456 3163
rect 2490 3129 2491 3163
rect 2455 3095 2491 3129
rect 2455 3061 2456 3095
rect 2490 3061 2491 3095
rect 2455 3027 2491 3061
rect 2455 2993 2456 3027
rect 2490 2993 2491 3027
rect 2455 2959 2491 2993
rect 2455 2925 2456 2959
rect 2490 2925 2491 2959
rect 2455 2891 2491 2925
rect 2455 2857 2456 2891
rect 2490 2857 2491 2891
rect 2455 2823 2491 2857
rect 2455 2789 2456 2823
rect 2490 2789 2491 2823
rect 2455 2755 2491 2789
rect 2455 2721 2456 2755
rect 2490 2721 2491 2755
rect 2455 2687 2491 2721
rect 2455 2653 2456 2687
rect 2490 2653 2491 2687
rect 2455 2619 2491 2653
rect 2455 2585 2456 2619
rect 2490 2585 2491 2619
rect 2455 2551 2491 2585
rect 2455 2517 2456 2551
rect 2490 2517 2491 2551
rect 2455 2483 2491 2517
rect 2455 2449 2456 2483
rect 2490 2449 2491 2483
rect 2455 2323 2491 2449
rect 232 2322 2491 2323
rect 232 2321 315 2322
rect 197 2288 315 2321
rect 349 2288 383 2322
rect 417 2288 451 2322
rect 485 2288 519 2322
rect 553 2288 587 2322
rect 621 2288 655 2322
rect 689 2288 723 2322
rect 757 2288 791 2322
rect 825 2288 859 2322
rect 893 2288 927 2322
rect 961 2288 995 2322
rect 1029 2288 1063 2322
rect 1097 2288 1131 2322
rect 1165 2288 1199 2322
rect 1233 2288 1267 2322
rect 1301 2288 1335 2322
rect 1369 2288 1403 2322
rect 1437 2288 1471 2322
rect 1505 2288 1539 2322
rect 1573 2288 1607 2322
rect 1641 2288 1675 2322
rect 1709 2288 1743 2322
rect 1777 2288 1811 2322
rect 1845 2288 1879 2322
rect 1913 2288 1947 2322
rect 1981 2288 2015 2322
rect 2049 2288 2083 2322
rect 2117 2288 2151 2322
rect 2185 2288 2219 2322
rect 2253 2288 2287 2322
rect 2321 2288 2355 2322
rect 2389 2288 2423 2322
rect 2457 2288 2491 2322
rect 197 2287 2491 2288
<< mvnsubdiff >>
rect 8 7351 2680 7352
rect 8 7317 85 7351
rect 119 7317 187 7351
rect 221 7317 255 7351
rect 289 7317 323 7351
rect 357 7317 391 7351
rect 425 7317 459 7351
rect 493 7317 527 7351
rect 561 7317 595 7351
rect 629 7317 663 7351
rect 697 7317 731 7351
rect 765 7317 799 7351
rect 833 7317 867 7351
rect 901 7317 935 7351
rect 969 7317 1003 7351
rect 1037 7317 1071 7351
rect 1105 7317 1139 7351
rect 1173 7317 1207 7351
rect 1241 7317 1275 7351
rect 1309 7317 1343 7351
rect 1377 7317 1411 7351
rect 1445 7317 1479 7351
rect 1513 7317 1547 7351
rect 1581 7317 1615 7351
rect 1649 7317 1683 7351
rect 1717 7317 1751 7351
rect 1785 7317 1819 7351
rect 1853 7317 1887 7351
rect 1921 7317 1955 7351
rect 1989 7317 2023 7351
rect 2057 7317 2091 7351
rect 2125 7317 2159 7351
rect 2193 7317 2227 7351
rect 2261 7317 2295 7351
rect 2329 7317 2363 7351
rect 2397 7317 2431 7351
rect 2465 7317 2499 7351
rect 2533 7317 2567 7351
rect 2601 7317 2680 7351
rect 8 7316 2680 7317
rect 8 7256 44 7316
rect 8 7222 9 7256
rect 43 7222 44 7256
rect 8 7188 44 7222
rect 8 7154 9 7188
rect 43 7154 44 7188
rect 8 7120 44 7154
rect 2644 7282 2680 7316
rect 2644 7248 2645 7282
rect 2679 7248 2680 7282
rect 2644 7214 2680 7248
rect 2644 7180 2645 7214
rect 2679 7180 2680 7214
rect 2644 7146 2680 7180
rect 8 7086 9 7120
rect 43 7086 44 7120
rect 8 7052 44 7086
rect 8 7018 9 7052
rect 43 7018 44 7052
rect 8 6984 44 7018
rect 8 6950 9 6984
rect 43 6950 44 6984
rect 8 6916 44 6950
rect 8 6882 9 6916
rect 43 6882 44 6916
rect 8 6848 44 6882
rect 8 6814 9 6848
rect 43 6814 44 6848
rect 8 6780 44 6814
rect 8 6746 9 6780
rect 43 6746 44 6780
rect 8 6712 44 6746
rect 8 6678 9 6712
rect 43 6678 44 6712
rect 8 6644 44 6678
rect 8 6610 9 6644
rect 43 6610 44 6644
rect 8 6576 44 6610
rect 8 6542 9 6576
rect 43 6542 44 6576
rect 8 6508 44 6542
rect 8 6474 9 6508
rect 43 6474 44 6508
rect 8 6440 44 6474
rect 8 6406 9 6440
rect 43 6406 44 6440
rect 8 6372 44 6406
rect 8 6338 9 6372
rect 43 6338 44 6372
rect 8 6304 44 6338
rect 8 6270 9 6304
rect 43 6270 44 6304
rect 8 6236 44 6270
rect 8 6202 9 6236
rect 43 6202 44 6236
rect 8 6168 44 6202
rect 8 6134 9 6168
rect 43 6134 44 6168
rect 8 6100 44 6134
rect 8 6066 9 6100
rect 43 6066 44 6100
rect 8 6032 44 6066
rect 8 5998 9 6032
rect 43 5998 44 6032
rect 8 5964 44 5998
rect 8 5930 9 5964
rect 43 5930 44 5964
rect 8 5896 44 5930
rect 8 5862 9 5896
rect 43 5862 44 5896
rect 8 5828 44 5862
rect 8 5794 9 5828
rect 43 5794 44 5828
rect 8 5760 44 5794
rect 8 5726 9 5760
rect 43 5726 44 5760
rect 8 5692 44 5726
rect 8 5658 9 5692
rect 43 5658 44 5692
rect 8 5624 44 5658
rect 8 5590 9 5624
rect 43 5590 44 5624
rect 8 5556 44 5590
rect 8 5522 9 5556
rect 43 5522 44 5556
rect 8 5488 44 5522
rect 8 5454 9 5488
rect 43 5454 44 5488
rect 8 5420 44 5454
rect 8 5386 9 5420
rect 43 5386 44 5420
rect 8 5352 44 5386
rect 8 5318 9 5352
rect 43 5318 44 5352
rect 8 5284 44 5318
rect 8 5250 9 5284
rect 43 5250 44 5284
rect 8 5216 44 5250
rect 8 5182 9 5216
rect 43 5182 44 5216
rect 8 5148 44 5182
rect 8 5114 9 5148
rect 43 5114 44 5148
rect 8 5080 44 5114
rect 8 5046 9 5080
rect 43 5046 44 5080
rect 8 5012 44 5046
rect 8 4978 9 5012
rect 43 4978 44 5012
rect 8 4944 44 4978
rect 8 4910 9 4944
rect 43 4910 44 4944
rect 8 4876 44 4910
rect 8 4842 9 4876
rect 43 4842 44 4876
rect 8 4808 44 4842
rect 8 4774 9 4808
rect 43 4774 44 4808
rect 8 4740 44 4774
rect 8 4706 9 4740
rect 43 4706 44 4740
rect 8 4672 44 4706
rect 8 4638 9 4672
rect 43 4638 44 4672
rect 8 4604 44 4638
rect 8 4570 9 4604
rect 43 4570 44 4604
rect 8 4536 44 4570
rect 8 4502 9 4536
rect 43 4502 44 4536
rect 8 4468 44 4502
rect 8 4434 9 4468
rect 43 4434 44 4468
rect 8 4400 44 4434
rect 8 4366 9 4400
rect 43 4366 44 4400
rect 8 4332 44 4366
rect 8 4298 9 4332
rect 43 4298 44 4332
rect 8 4264 44 4298
rect 8 4230 9 4264
rect 43 4230 44 4264
rect 8 4196 44 4230
rect 8 4162 9 4196
rect 43 4162 44 4196
rect 8 4128 44 4162
rect 8 4094 9 4128
rect 43 4094 44 4128
rect 8 4060 44 4094
rect 8 4026 9 4060
rect 43 4026 44 4060
rect 8 3992 44 4026
rect 8 3958 9 3992
rect 43 3958 44 3992
rect 8 3924 44 3958
rect 8 3890 9 3924
rect 43 3890 44 3924
rect 8 3856 44 3890
rect 8 3822 9 3856
rect 43 3822 44 3856
rect 8 3788 44 3822
rect 8 3754 9 3788
rect 43 3754 44 3788
rect 8 3720 44 3754
rect 8 3686 9 3720
rect 43 3686 44 3720
rect 8 3652 44 3686
rect 8 3618 9 3652
rect 43 3618 44 3652
rect 8 3584 44 3618
rect 8 3550 9 3584
rect 43 3550 44 3584
rect 8 3516 44 3550
rect 8 3482 9 3516
rect 43 3482 44 3516
rect 8 3448 44 3482
rect 8 3414 9 3448
rect 43 3414 44 3448
rect 8 3380 44 3414
rect 8 3346 9 3380
rect 43 3346 44 3380
rect 8 3312 44 3346
rect 8 3278 9 3312
rect 43 3278 44 3312
rect 8 3244 44 3278
rect 8 3210 9 3244
rect 43 3210 44 3244
rect 8 3176 44 3210
rect 8 3142 9 3176
rect 43 3142 44 3176
rect 8 3108 44 3142
rect 8 3074 9 3108
rect 43 3074 44 3108
rect 8 3040 44 3074
rect 8 3006 9 3040
rect 43 3006 44 3040
rect 8 2972 44 3006
rect 8 2938 9 2972
rect 43 2938 44 2972
rect 8 2904 44 2938
rect 8 2870 9 2904
rect 43 2870 44 2904
rect 8 2836 44 2870
rect 8 2802 9 2836
rect 43 2802 44 2836
rect 8 2768 44 2802
rect 8 2734 9 2768
rect 43 2734 44 2768
rect 8 2700 44 2734
rect 8 2666 9 2700
rect 43 2666 44 2700
rect 8 2632 44 2666
rect 8 2598 9 2632
rect 43 2598 44 2632
rect 8 2564 44 2598
rect 8 2530 9 2564
rect 43 2530 44 2564
rect 8 2496 44 2530
rect 8 2462 9 2496
rect 43 2462 44 2496
rect 8 2428 44 2462
rect 8 2394 9 2428
rect 43 2394 44 2428
rect 8 2360 44 2394
rect 8 2326 9 2360
rect 43 2326 44 2360
rect 8 2292 44 2326
rect 8 2258 9 2292
rect 43 2258 44 2292
rect 2644 7112 2645 7146
rect 2679 7112 2680 7146
rect 2644 7078 2680 7112
rect 2644 7044 2645 7078
rect 2679 7044 2680 7078
rect 2644 7010 2680 7044
rect 2644 6976 2645 7010
rect 2679 6976 2680 7010
rect 2644 6942 2680 6976
rect 2644 6908 2645 6942
rect 2679 6908 2680 6942
rect 2644 6874 2680 6908
rect 2644 6840 2645 6874
rect 2679 6840 2680 6874
rect 2644 6806 2680 6840
rect 2644 6772 2645 6806
rect 2679 6772 2680 6806
rect 2644 6738 2680 6772
rect 2644 6704 2645 6738
rect 2679 6704 2680 6738
rect 2644 6670 2680 6704
rect 2644 6636 2645 6670
rect 2679 6636 2680 6670
rect 2644 6602 2680 6636
rect 2644 6568 2645 6602
rect 2679 6568 2680 6602
rect 2644 6534 2680 6568
rect 2644 6500 2645 6534
rect 2679 6500 2680 6534
rect 2644 6466 2680 6500
rect 2644 6432 2645 6466
rect 2679 6432 2680 6466
rect 2644 6398 2680 6432
rect 2644 6364 2645 6398
rect 2679 6364 2680 6398
rect 2644 6330 2680 6364
rect 2644 6296 2645 6330
rect 2679 6296 2680 6330
rect 2644 6262 2680 6296
rect 2644 6228 2645 6262
rect 2679 6228 2680 6262
rect 2644 6194 2680 6228
rect 2644 6160 2645 6194
rect 2679 6160 2680 6194
rect 2644 6126 2680 6160
rect 2644 6092 2645 6126
rect 2679 6092 2680 6126
rect 2644 6058 2680 6092
rect 2644 6024 2645 6058
rect 2679 6024 2680 6058
rect 2644 5990 2680 6024
rect 2644 5956 2645 5990
rect 2679 5956 2680 5990
rect 2644 5922 2680 5956
rect 2644 5888 2645 5922
rect 2679 5888 2680 5922
rect 2644 5854 2680 5888
rect 2644 5820 2645 5854
rect 2679 5820 2680 5854
rect 2644 5786 2680 5820
rect 2644 5752 2645 5786
rect 2679 5752 2680 5786
rect 2644 5718 2680 5752
rect 2644 5684 2645 5718
rect 2679 5684 2680 5718
rect 2644 5650 2680 5684
rect 2644 5616 2645 5650
rect 2679 5616 2680 5650
rect 2644 5582 2680 5616
rect 2644 5548 2645 5582
rect 2679 5548 2680 5582
rect 2644 5514 2680 5548
rect 2644 5480 2645 5514
rect 2679 5480 2680 5514
rect 2644 5446 2680 5480
rect 2644 5412 2645 5446
rect 2679 5412 2680 5446
rect 2644 5378 2680 5412
rect 2644 5344 2645 5378
rect 2679 5344 2680 5378
rect 2644 5310 2680 5344
rect 2644 5276 2645 5310
rect 2679 5276 2680 5310
rect 2644 5242 2680 5276
rect 2644 5208 2645 5242
rect 2679 5208 2680 5242
rect 2644 5174 2680 5208
rect 2644 5140 2645 5174
rect 2679 5140 2680 5174
rect 2644 5106 2680 5140
rect 2644 5072 2645 5106
rect 2679 5072 2680 5106
rect 2644 5038 2680 5072
rect 2644 5004 2645 5038
rect 2679 5004 2680 5038
rect 2644 4970 2680 5004
rect 2644 4936 2645 4970
rect 2679 4936 2680 4970
rect 2644 4902 2680 4936
rect 2644 4868 2645 4902
rect 2679 4868 2680 4902
rect 2644 4834 2680 4868
rect 2644 4800 2645 4834
rect 2679 4800 2680 4834
rect 2644 4766 2680 4800
rect 2644 4732 2645 4766
rect 2679 4732 2680 4766
rect 2644 4698 2680 4732
rect 2644 4664 2645 4698
rect 2679 4664 2680 4698
rect 2644 4630 2680 4664
rect 2644 4596 2645 4630
rect 2679 4596 2680 4630
rect 2644 4562 2680 4596
rect 2644 4528 2645 4562
rect 2679 4528 2680 4562
rect 2644 4494 2680 4528
rect 2644 4460 2645 4494
rect 2679 4460 2680 4494
rect 2644 4426 2680 4460
rect 2644 4392 2645 4426
rect 2679 4392 2680 4426
rect 2644 4358 2680 4392
rect 2644 4324 2645 4358
rect 2679 4324 2680 4358
rect 2644 4290 2680 4324
rect 2644 4256 2645 4290
rect 2679 4256 2680 4290
rect 2644 4222 2680 4256
rect 2644 4188 2645 4222
rect 2679 4188 2680 4222
rect 2644 4154 2680 4188
rect 2644 4120 2645 4154
rect 2679 4120 2680 4154
rect 2644 4086 2680 4120
rect 2644 4052 2645 4086
rect 2679 4052 2680 4086
rect 2644 4018 2680 4052
rect 2644 3984 2645 4018
rect 2679 3984 2680 4018
rect 2644 3950 2680 3984
rect 2644 3916 2645 3950
rect 2679 3916 2680 3950
rect 2644 3882 2680 3916
rect 2644 3848 2645 3882
rect 2679 3848 2680 3882
rect 2644 3814 2680 3848
rect 2644 3780 2645 3814
rect 2679 3780 2680 3814
rect 2644 3746 2680 3780
rect 2644 3712 2645 3746
rect 2679 3712 2680 3746
rect 2644 3678 2680 3712
rect 2644 3644 2645 3678
rect 2679 3644 2680 3678
rect 2644 3610 2680 3644
rect 2644 3576 2645 3610
rect 2679 3576 2680 3610
rect 2644 3542 2680 3576
rect 2644 3508 2645 3542
rect 2679 3508 2680 3542
rect 2644 3474 2680 3508
rect 2644 3440 2645 3474
rect 2679 3440 2680 3474
rect 2644 3406 2680 3440
rect 2644 3372 2645 3406
rect 2679 3372 2680 3406
rect 2644 3338 2680 3372
rect 2644 3304 2645 3338
rect 2679 3304 2680 3338
rect 2644 3270 2680 3304
rect 2644 3236 2645 3270
rect 2679 3236 2680 3270
rect 2644 3202 2680 3236
rect 2644 3168 2645 3202
rect 2679 3168 2680 3202
rect 2644 3134 2680 3168
rect 2644 3100 2645 3134
rect 2679 3100 2680 3134
rect 2644 3066 2680 3100
rect 2644 3032 2645 3066
rect 2679 3032 2680 3066
rect 2644 2998 2680 3032
rect 2644 2964 2645 2998
rect 2679 2964 2680 2998
rect 2644 2930 2680 2964
rect 2644 2896 2645 2930
rect 2679 2896 2680 2930
rect 2644 2862 2680 2896
rect 2644 2828 2645 2862
rect 2679 2828 2680 2862
rect 2644 2794 2680 2828
rect 2644 2760 2645 2794
rect 2679 2760 2680 2794
rect 2644 2726 2680 2760
rect 2644 2692 2645 2726
rect 2679 2692 2680 2726
rect 2644 2658 2680 2692
rect 2644 2624 2645 2658
rect 2679 2624 2680 2658
rect 2644 2590 2680 2624
rect 2644 2556 2645 2590
rect 2679 2556 2680 2590
rect 2644 2522 2680 2556
rect 2644 2488 2645 2522
rect 2679 2488 2680 2522
rect 2644 2454 2680 2488
rect 2644 2420 2645 2454
rect 2679 2420 2680 2454
rect 2644 2386 2680 2420
rect 2644 2352 2645 2386
rect 2679 2352 2680 2386
rect 2644 2318 2680 2352
rect 8 2224 44 2258
rect 8 2190 9 2224
rect 43 2190 44 2224
rect 8 2156 44 2190
rect 8 2122 9 2156
rect 43 2134 44 2156
rect 2644 2284 2645 2318
rect 2679 2284 2680 2318
rect 2644 2250 2680 2284
rect 2644 2216 2645 2250
rect 2679 2216 2680 2250
rect 2644 2182 2680 2216
rect 2644 2148 2645 2182
rect 2679 2148 2680 2182
rect 2644 2134 2680 2148
rect 43 2133 2680 2134
rect 43 2122 128 2133
rect 8 2099 128 2122
rect 162 2099 196 2133
rect 230 2099 264 2133
rect 298 2099 332 2133
rect 366 2099 400 2133
rect 434 2099 468 2133
rect 502 2099 536 2133
rect 570 2099 604 2133
rect 638 2099 672 2133
rect 706 2099 740 2133
rect 774 2099 808 2133
rect 842 2099 876 2133
rect 910 2099 944 2133
rect 978 2099 1012 2133
rect 1046 2099 1080 2133
rect 1114 2099 1148 2133
rect 1182 2099 1216 2133
rect 1250 2099 1284 2133
rect 1318 2099 1352 2133
rect 1386 2099 1420 2133
rect 1454 2099 1488 2133
rect 1522 2099 1556 2133
rect 1590 2099 1624 2133
rect 1658 2099 1692 2133
rect 1726 2099 1760 2133
rect 1794 2099 1828 2133
rect 1862 2099 1896 2133
rect 1930 2099 1964 2133
rect 1998 2099 2032 2133
rect 2066 2099 2100 2133
rect 2134 2099 2168 2133
rect 2202 2099 2236 2133
rect 2270 2099 2304 2133
rect 2338 2099 2372 2133
rect 2406 2099 2440 2133
rect 2474 2099 2508 2133
rect 2542 2099 2576 2133
rect 2610 2114 2680 2133
rect 2610 2099 2645 2114
rect 8 2098 2645 2099
rect 8 2088 44 2098
rect 8 2054 9 2088
rect 43 2054 44 2088
rect 2644 2080 2645 2098
rect 2679 2080 2680 2114
rect 8 2020 44 2054
rect 8 1986 9 2020
rect 43 1986 44 2020
rect 8 1952 44 1986
rect 8 1918 9 1952
rect 43 1918 44 1952
rect 2644 2046 2680 2080
rect 2644 2012 2645 2046
rect 2679 2012 2680 2046
rect 2644 1978 2680 2012
rect 2644 1944 2645 1978
rect 2679 1944 2680 1978
rect 8 1884 44 1918
rect 8 1850 9 1884
rect 43 1850 44 1884
rect 8 1816 44 1850
rect 8 1782 9 1816
rect 43 1782 44 1816
rect 8 1748 44 1782
rect 8 1714 9 1748
rect 43 1714 44 1748
rect 8 1680 44 1714
rect 8 1646 9 1680
rect 43 1646 44 1680
rect 8 1612 44 1646
rect 8 1578 9 1612
rect 43 1578 44 1612
rect 8 1544 44 1578
rect 8 1510 9 1544
rect 43 1510 44 1544
rect 8 1476 44 1510
rect 8 1442 9 1476
rect 43 1442 44 1476
rect 8 1408 44 1442
rect 8 1374 9 1408
rect 43 1374 44 1408
rect 8 1340 44 1374
rect 8 1306 9 1340
rect 43 1306 44 1340
rect 8 1272 44 1306
rect 8 1238 9 1272
rect 43 1238 44 1272
rect 8 1204 44 1238
rect 8 1170 9 1204
rect 43 1170 44 1204
rect 8 1136 44 1170
rect 8 1102 9 1136
rect 43 1102 44 1136
rect 8 1068 44 1102
rect 8 1034 9 1068
rect 43 1034 44 1068
rect 8 1000 44 1034
rect 8 966 9 1000
rect 43 966 44 1000
rect 8 932 44 966
rect 8 898 9 932
rect 43 898 44 932
rect 8 864 44 898
rect 8 830 9 864
rect 43 830 44 864
rect 8 796 44 830
rect 8 762 9 796
rect 43 762 44 796
rect 8 728 44 762
rect 8 694 9 728
rect 43 694 44 728
rect 8 660 44 694
rect 8 626 9 660
rect 43 626 44 660
rect 8 592 44 626
rect 8 558 9 592
rect 43 558 44 592
rect 8 524 44 558
rect 2644 1910 2680 1944
rect 2644 1876 2645 1910
rect 2679 1876 2680 1910
rect 2644 1842 2680 1876
rect 2644 1808 2645 1842
rect 2679 1808 2680 1842
rect 2644 1774 2680 1808
rect 2644 1740 2645 1774
rect 2679 1740 2680 1774
rect 2644 1706 2680 1740
rect 2644 1672 2645 1706
rect 2679 1672 2680 1706
rect 2644 1638 2680 1672
rect 2644 1604 2645 1638
rect 2679 1604 2680 1638
rect 2644 1570 2680 1604
rect 2644 1536 2645 1570
rect 2679 1536 2680 1570
rect 2644 1502 2680 1536
rect 2644 1468 2645 1502
rect 2679 1468 2680 1502
rect 2644 1434 2680 1468
rect 2644 1400 2645 1434
rect 2679 1400 2680 1434
rect 2644 1366 2680 1400
rect 2644 1332 2645 1366
rect 2679 1332 2680 1366
rect 2644 1298 2680 1332
rect 2644 1264 2645 1298
rect 2679 1264 2680 1298
rect 2644 1230 2680 1264
rect 2644 1196 2645 1230
rect 2679 1196 2680 1230
rect 2644 1162 2680 1196
rect 2644 1128 2645 1162
rect 2679 1128 2680 1162
rect 2644 1094 2680 1128
rect 2644 1060 2645 1094
rect 2679 1060 2680 1094
rect 2644 1026 2680 1060
rect 2644 992 2645 1026
rect 2679 992 2680 1026
rect 2644 958 2680 992
rect 2644 924 2645 958
rect 2679 924 2680 958
rect 2644 890 2680 924
rect 2644 856 2645 890
rect 2679 856 2680 890
rect 2644 822 2680 856
rect 2644 788 2645 822
rect 2679 788 2680 822
rect 2644 754 2680 788
rect 2644 720 2645 754
rect 2679 720 2680 754
rect 2644 686 2680 720
rect 2644 652 2645 686
rect 2679 652 2680 686
rect 2644 618 2680 652
rect 2644 584 2645 618
rect 2679 584 2680 618
rect 2644 550 2680 584
rect 8 490 9 524
rect 43 490 44 524
rect 8 329 44 490
rect 8 295 9 329
rect 43 295 44 329
rect 8 261 44 295
rect 8 227 9 261
rect 43 227 44 261
rect 8 193 44 227
rect 8 159 9 193
rect 43 159 44 193
rect 8 125 44 159
rect 2644 516 2645 550
rect 2679 516 2680 550
rect 2644 482 2680 516
rect 2644 448 2645 482
rect 2679 448 2680 482
rect 2644 414 2680 448
rect 2644 380 2645 414
rect 2679 380 2680 414
rect 2644 346 2680 380
rect 2644 312 2645 346
rect 2679 312 2680 346
rect 2644 278 2680 312
rect 2644 244 2645 278
rect 2679 244 2680 278
rect 2644 210 2680 244
rect 2644 176 2645 210
rect 2679 176 2680 210
rect 8 91 9 125
rect 43 91 44 125
rect 8 57 44 91
rect 2644 142 2680 176
rect 2644 108 2645 142
rect 2679 108 2680 142
rect 2644 57 2680 108
<< mvpsubdiffcont >>
rect 89 7506 123 7540
rect 157 7506 191 7540
rect 225 7506 259 7540
rect 293 7506 327 7540
rect 361 7506 395 7540
rect 429 7506 463 7540
rect 497 7506 531 7540
rect 565 7506 599 7540
rect 633 7506 667 7540
rect 701 7506 735 7540
rect 769 7506 803 7540
rect 837 7506 871 7540
rect 905 7506 939 7540
rect 973 7506 1007 7540
rect 1041 7506 1075 7540
rect 1109 7506 1143 7540
rect 1177 7506 1211 7540
rect 1245 7506 1279 7540
rect 1313 7506 1347 7540
rect 1381 7506 1415 7540
rect 1449 7506 1483 7540
rect 1517 7506 1551 7540
rect 1585 7506 1619 7540
rect 1653 7506 1687 7540
rect 1721 7506 1755 7540
rect 1789 7506 1823 7540
rect 1857 7506 1891 7540
rect 1925 7506 1959 7540
rect 1993 7506 2027 7540
rect 2061 7506 2095 7540
rect 2129 7506 2163 7540
rect 2197 7506 2231 7540
rect 2265 7506 2299 7540
rect 2333 7506 2367 7540
rect 2401 7506 2435 7540
rect 2469 7506 2503 7540
rect 2537 7506 2571 7540
rect 2605 7506 2639 7540
rect 231 7106 265 7140
rect 299 7106 333 7140
rect 367 7106 401 7140
rect 435 7106 469 7140
rect 503 7106 537 7140
rect 571 7106 605 7140
rect 639 7106 673 7140
rect 707 7106 741 7140
rect 775 7106 809 7140
rect 843 7106 877 7140
rect 911 7106 945 7140
rect 979 7106 1013 7140
rect 1047 7106 1081 7140
rect 1115 7106 1149 7140
rect 1183 7106 1217 7140
rect 1251 7106 1285 7140
rect 1319 7106 1353 7140
rect 1387 7106 1421 7140
rect 1455 7106 1489 7140
rect 1523 7106 1557 7140
rect 1591 7106 1625 7140
rect 1659 7106 1693 7140
rect 1727 7106 1761 7140
rect 1795 7106 1829 7140
rect 1863 7106 1897 7140
rect 1931 7106 1965 7140
rect 1999 7106 2033 7140
rect 2067 7106 2101 7140
rect 2135 7106 2169 7140
rect 2203 7106 2237 7140
rect 2271 7106 2305 7140
rect 2339 7106 2373 7140
rect 2456 7073 2490 7107
rect 198 7013 232 7047
rect 2456 7005 2490 7039
rect 198 6945 232 6979
rect 198 6877 232 6911
rect 198 6809 232 6843
rect 198 6741 232 6775
rect 198 6673 232 6707
rect 198 6605 232 6639
rect 198 6537 232 6571
rect 198 6469 232 6503
rect 198 6401 232 6435
rect 198 6333 232 6367
rect 198 6265 232 6299
rect 198 6197 232 6231
rect 198 6129 232 6163
rect 198 6061 232 6095
rect 198 5993 232 6027
rect 198 5925 232 5959
rect 2456 6937 2490 6971
rect 2456 6869 2490 6903
rect 2456 6801 2490 6835
rect 2456 6733 2490 6767
rect 2456 6665 2490 6699
rect 2456 6597 2490 6631
rect 2456 6529 2490 6563
rect 2456 6461 2490 6495
rect 2456 6393 2490 6427
rect 2456 6325 2490 6359
rect 2456 6257 2490 6291
rect 2456 6189 2490 6223
rect 2456 6121 2490 6155
rect 2456 6053 2490 6087
rect 2456 5985 2490 6019
rect 198 5857 232 5891
rect 2456 5917 2490 5951
rect 198 5789 232 5823
rect 2456 5849 2490 5883
rect 198 5721 232 5755
rect 198 5653 232 5687
rect 198 5585 232 5619
rect 198 5517 232 5551
rect 198 5449 232 5483
rect 198 5381 232 5415
rect 198 5313 232 5347
rect 198 5245 232 5279
rect 198 5177 232 5211
rect 198 5109 232 5143
rect 198 5041 232 5075
rect 198 4973 232 5007
rect 198 4905 232 4939
rect 198 4837 232 4871
rect 198 4769 232 4803
rect 198 4701 232 4735
rect 2456 5781 2490 5815
rect 2456 5713 2490 5747
rect 2456 5645 2490 5679
rect 2456 5577 2490 5611
rect 2456 5509 2490 5543
rect 2456 5441 2490 5475
rect 2456 5373 2490 5407
rect 2456 5305 2490 5339
rect 2456 5237 2490 5271
rect 2456 5169 2490 5203
rect 2456 5101 2490 5135
rect 2456 5033 2490 5067
rect 2456 4965 2490 4999
rect 2456 4897 2490 4931
rect 2456 4829 2490 4863
rect 2456 4761 2490 4795
rect 2456 4693 2490 4727
rect 198 4633 232 4667
rect 2456 4625 2490 4659
rect 198 4565 232 4599
rect 198 4497 232 4531
rect 198 4429 232 4463
rect 198 4361 232 4395
rect 198 4293 232 4327
rect 198 4225 232 4259
rect 198 4157 232 4191
rect 198 4089 232 4123
rect 198 4021 232 4055
rect 198 3953 232 3987
rect 198 3885 232 3919
rect 198 3817 232 3851
rect 198 3749 232 3783
rect 198 3681 232 3715
rect 198 3613 232 3647
rect 198 3545 232 3579
rect 2456 4557 2490 4591
rect 2456 4489 2490 4523
rect 2456 4421 2490 4455
rect 2456 4353 2490 4387
rect 2456 4285 2490 4319
rect 2456 4217 2490 4251
rect 2456 4149 2490 4183
rect 2456 4081 2490 4115
rect 2456 4013 2490 4047
rect 2456 3945 2490 3979
rect 2456 3877 2490 3911
rect 2456 3809 2490 3843
rect 2456 3741 2490 3775
rect 2456 3673 2490 3707
rect 2456 3605 2490 3639
rect 2456 3537 2490 3571
rect 198 3477 232 3511
rect 198 3409 232 3443
rect 2456 3469 2490 3503
rect 198 3341 232 3375
rect 198 3273 232 3307
rect 198 3205 232 3239
rect 198 3137 232 3171
rect 198 3069 232 3103
rect 198 3001 232 3035
rect 198 2933 232 2967
rect 198 2865 232 2899
rect 198 2797 232 2831
rect 198 2729 232 2763
rect 198 2661 232 2695
rect 198 2593 232 2627
rect 198 2525 232 2559
rect 198 2457 232 2491
rect 198 2389 232 2423
rect 198 2321 232 2355
rect 2456 3401 2490 3435
rect 2456 3333 2490 3367
rect 2456 3265 2490 3299
rect 2456 3197 2490 3231
rect 2456 3129 2490 3163
rect 2456 3061 2490 3095
rect 2456 2993 2490 3027
rect 2456 2925 2490 2959
rect 2456 2857 2490 2891
rect 2456 2789 2490 2823
rect 2456 2721 2490 2755
rect 2456 2653 2490 2687
rect 2456 2585 2490 2619
rect 2456 2517 2490 2551
rect 2456 2449 2490 2483
rect 315 2288 349 2322
rect 383 2288 417 2322
rect 451 2288 485 2322
rect 519 2288 553 2322
rect 587 2288 621 2322
rect 655 2288 689 2322
rect 723 2288 757 2322
rect 791 2288 825 2322
rect 859 2288 893 2322
rect 927 2288 961 2322
rect 995 2288 1029 2322
rect 1063 2288 1097 2322
rect 1131 2288 1165 2322
rect 1199 2288 1233 2322
rect 1267 2288 1301 2322
rect 1335 2288 1369 2322
rect 1403 2288 1437 2322
rect 1471 2288 1505 2322
rect 1539 2288 1573 2322
rect 1607 2288 1641 2322
rect 1675 2288 1709 2322
rect 1743 2288 1777 2322
rect 1811 2288 1845 2322
rect 1879 2288 1913 2322
rect 1947 2288 1981 2322
rect 2015 2288 2049 2322
rect 2083 2288 2117 2322
rect 2151 2288 2185 2322
rect 2219 2288 2253 2322
rect 2287 2288 2321 2322
rect 2355 2288 2389 2322
rect 2423 2288 2457 2322
<< mvnsubdiffcont >>
rect 85 7317 119 7351
rect 187 7317 221 7351
rect 255 7317 289 7351
rect 323 7317 357 7351
rect 391 7317 425 7351
rect 459 7317 493 7351
rect 527 7317 561 7351
rect 595 7317 629 7351
rect 663 7317 697 7351
rect 731 7317 765 7351
rect 799 7317 833 7351
rect 867 7317 901 7351
rect 935 7317 969 7351
rect 1003 7317 1037 7351
rect 1071 7317 1105 7351
rect 1139 7317 1173 7351
rect 1207 7317 1241 7351
rect 1275 7317 1309 7351
rect 1343 7317 1377 7351
rect 1411 7317 1445 7351
rect 1479 7317 1513 7351
rect 1547 7317 1581 7351
rect 1615 7317 1649 7351
rect 1683 7317 1717 7351
rect 1751 7317 1785 7351
rect 1819 7317 1853 7351
rect 1887 7317 1921 7351
rect 1955 7317 1989 7351
rect 2023 7317 2057 7351
rect 2091 7317 2125 7351
rect 2159 7317 2193 7351
rect 2227 7317 2261 7351
rect 2295 7317 2329 7351
rect 2363 7317 2397 7351
rect 2431 7317 2465 7351
rect 2499 7317 2533 7351
rect 2567 7317 2601 7351
rect 9 7222 43 7256
rect 9 7154 43 7188
rect 2645 7248 2679 7282
rect 2645 7180 2679 7214
rect 9 7086 43 7120
rect 9 7018 43 7052
rect 9 6950 43 6984
rect 9 6882 43 6916
rect 9 6814 43 6848
rect 9 6746 43 6780
rect 9 6678 43 6712
rect 9 6610 43 6644
rect 9 6542 43 6576
rect 9 6474 43 6508
rect 9 6406 43 6440
rect 9 6338 43 6372
rect 9 6270 43 6304
rect 9 6202 43 6236
rect 9 6134 43 6168
rect 9 6066 43 6100
rect 9 5998 43 6032
rect 9 5930 43 5964
rect 9 5862 43 5896
rect 9 5794 43 5828
rect 9 5726 43 5760
rect 9 5658 43 5692
rect 9 5590 43 5624
rect 9 5522 43 5556
rect 9 5454 43 5488
rect 9 5386 43 5420
rect 9 5318 43 5352
rect 9 5250 43 5284
rect 9 5182 43 5216
rect 9 5114 43 5148
rect 9 5046 43 5080
rect 9 4978 43 5012
rect 9 4910 43 4944
rect 9 4842 43 4876
rect 9 4774 43 4808
rect 9 4706 43 4740
rect 9 4638 43 4672
rect 9 4570 43 4604
rect 9 4502 43 4536
rect 9 4434 43 4468
rect 9 4366 43 4400
rect 9 4298 43 4332
rect 9 4230 43 4264
rect 9 4162 43 4196
rect 9 4094 43 4128
rect 9 4026 43 4060
rect 9 3958 43 3992
rect 9 3890 43 3924
rect 9 3822 43 3856
rect 9 3754 43 3788
rect 9 3686 43 3720
rect 9 3618 43 3652
rect 9 3550 43 3584
rect 9 3482 43 3516
rect 9 3414 43 3448
rect 9 3346 43 3380
rect 9 3278 43 3312
rect 9 3210 43 3244
rect 9 3142 43 3176
rect 9 3074 43 3108
rect 9 3006 43 3040
rect 9 2938 43 2972
rect 9 2870 43 2904
rect 9 2802 43 2836
rect 9 2734 43 2768
rect 9 2666 43 2700
rect 9 2598 43 2632
rect 9 2530 43 2564
rect 9 2462 43 2496
rect 9 2394 43 2428
rect 9 2326 43 2360
rect 9 2258 43 2292
rect 2645 7112 2679 7146
rect 2645 7044 2679 7078
rect 2645 6976 2679 7010
rect 2645 6908 2679 6942
rect 2645 6840 2679 6874
rect 2645 6772 2679 6806
rect 2645 6704 2679 6738
rect 2645 6636 2679 6670
rect 2645 6568 2679 6602
rect 2645 6500 2679 6534
rect 2645 6432 2679 6466
rect 2645 6364 2679 6398
rect 2645 6296 2679 6330
rect 2645 6228 2679 6262
rect 2645 6160 2679 6194
rect 2645 6092 2679 6126
rect 2645 6024 2679 6058
rect 2645 5956 2679 5990
rect 2645 5888 2679 5922
rect 2645 5820 2679 5854
rect 2645 5752 2679 5786
rect 2645 5684 2679 5718
rect 2645 5616 2679 5650
rect 2645 5548 2679 5582
rect 2645 5480 2679 5514
rect 2645 5412 2679 5446
rect 2645 5344 2679 5378
rect 2645 5276 2679 5310
rect 2645 5208 2679 5242
rect 2645 5140 2679 5174
rect 2645 5072 2679 5106
rect 2645 5004 2679 5038
rect 2645 4936 2679 4970
rect 2645 4868 2679 4902
rect 2645 4800 2679 4834
rect 2645 4732 2679 4766
rect 2645 4664 2679 4698
rect 2645 4596 2679 4630
rect 2645 4528 2679 4562
rect 2645 4460 2679 4494
rect 2645 4392 2679 4426
rect 2645 4324 2679 4358
rect 2645 4256 2679 4290
rect 2645 4188 2679 4222
rect 2645 4120 2679 4154
rect 2645 4052 2679 4086
rect 2645 3984 2679 4018
rect 2645 3916 2679 3950
rect 2645 3848 2679 3882
rect 2645 3780 2679 3814
rect 2645 3712 2679 3746
rect 2645 3644 2679 3678
rect 2645 3576 2679 3610
rect 2645 3508 2679 3542
rect 2645 3440 2679 3474
rect 2645 3372 2679 3406
rect 2645 3304 2679 3338
rect 2645 3236 2679 3270
rect 2645 3168 2679 3202
rect 2645 3100 2679 3134
rect 2645 3032 2679 3066
rect 2645 2964 2679 2998
rect 2645 2896 2679 2930
rect 2645 2828 2679 2862
rect 2645 2760 2679 2794
rect 2645 2692 2679 2726
rect 2645 2624 2679 2658
rect 2645 2556 2679 2590
rect 2645 2488 2679 2522
rect 2645 2420 2679 2454
rect 2645 2352 2679 2386
rect 9 2190 43 2224
rect 9 2122 43 2156
rect 2645 2284 2679 2318
rect 2645 2216 2679 2250
rect 2645 2148 2679 2182
rect 128 2099 162 2133
rect 196 2099 230 2133
rect 264 2099 298 2133
rect 332 2099 366 2133
rect 400 2099 434 2133
rect 468 2099 502 2133
rect 536 2099 570 2133
rect 604 2099 638 2133
rect 672 2099 706 2133
rect 740 2099 774 2133
rect 808 2099 842 2133
rect 876 2099 910 2133
rect 944 2099 978 2133
rect 1012 2099 1046 2133
rect 1080 2099 1114 2133
rect 1148 2099 1182 2133
rect 1216 2099 1250 2133
rect 1284 2099 1318 2133
rect 1352 2099 1386 2133
rect 1420 2099 1454 2133
rect 1488 2099 1522 2133
rect 1556 2099 1590 2133
rect 1624 2099 1658 2133
rect 1692 2099 1726 2133
rect 1760 2099 1794 2133
rect 1828 2099 1862 2133
rect 1896 2099 1930 2133
rect 1964 2099 1998 2133
rect 2032 2099 2066 2133
rect 2100 2099 2134 2133
rect 2168 2099 2202 2133
rect 2236 2099 2270 2133
rect 2304 2099 2338 2133
rect 2372 2099 2406 2133
rect 2440 2099 2474 2133
rect 2508 2099 2542 2133
rect 2576 2099 2610 2133
rect 9 2054 43 2088
rect 2645 2080 2679 2114
rect 9 1986 43 2020
rect 9 1918 43 1952
rect 2645 2012 2679 2046
rect 2645 1944 2679 1978
rect 9 1850 43 1884
rect 9 1782 43 1816
rect 9 1714 43 1748
rect 9 1646 43 1680
rect 9 1578 43 1612
rect 9 1510 43 1544
rect 9 1442 43 1476
rect 9 1374 43 1408
rect 9 1306 43 1340
rect 9 1238 43 1272
rect 9 1170 43 1204
rect 9 1102 43 1136
rect 9 1034 43 1068
rect 9 966 43 1000
rect 9 898 43 932
rect 9 830 43 864
rect 9 762 43 796
rect 9 694 43 728
rect 9 626 43 660
rect 9 558 43 592
rect 2645 1876 2679 1910
rect 2645 1808 2679 1842
rect 2645 1740 2679 1774
rect 2645 1672 2679 1706
rect 2645 1604 2679 1638
rect 2645 1536 2679 1570
rect 2645 1468 2679 1502
rect 2645 1400 2679 1434
rect 2645 1332 2679 1366
rect 2645 1264 2679 1298
rect 2645 1196 2679 1230
rect 2645 1128 2679 1162
rect 2645 1060 2679 1094
rect 2645 992 2679 1026
rect 2645 924 2679 958
rect 2645 856 2679 890
rect 2645 788 2679 822
rect 2645 720 2679 754
rect 2645 652 2679 686
rect 2645 584 2679 618
rect 9 490 43 524
rect 9 295 43 329
rect 9 227 43 261
rect 9 159 43 193
rect 2645 516 2679 550
rect 2645 448 2679 482
rect 2645 380 2679 414
rect 2645 312 2679 346
rect 2645 244 2679 278
rect 2645 176 2679 210
rect 9 91 43 125
rect 2645 108 2679 142
<< poly >>
rect 300 8722 500 8738
rect 300 8688 349 8722
rect 383 8688 417 8722
rect 451 8688 500 8722
rect 300 8666 500 8688
rect 556 8722 756 8738
rect 556 8688 605 8722
rect 639 8688 673 8722
rect 707 8688 756 8722
rect 556 8666 756 8688
rect 812 8722 1012 8738
rect 812 8688 861 8722
rect 895 8688 929 8722
rect 963 8688 1012 8722
rect 812 8666 1012 8688
rect 1068 8722 1268 8738
rect 1068 8688 1117 8722
rect 1151 8688 1185 8722
rect 1219 8688 1268 8722
rect 1068 8666 1268 8688
rect 1324 8722 1524 8738
rect 1324 8688 1373 8722
rect 1407 8688 1441 8722
rect 1475 8688 1524 8722
rect 1324 8666 1524 8688
rect 1580 8722 1780 8738
rect 1580 8688 1629 8722
rect 1663 8688 1697 8722
rect 1731 8688 1780 8722
rect 1580 8666 1780 8688
rect 1836 8722 2036 8738
rect 1836 8688 1885 8722
rect 1919 8688 1953 8722
rect 1987 8688 2036 8722
rect 1836 8666 2036 8688
rect 2092 8722 2292 8738
rect 2092 8688 2141 8722
rect 2175 8688 2209 8722
rect 2243 8688 2292 8722
rect 2092 8666 2292 8688
rect 326 7055 460 7071
rect 326 7021 342 7055
rect 376 7021 410 7055
rect 444 7021 460 7055
rect 326 7005 460 7021
rect 516 6999 1316 7071
rect 1372 6999 2172 7071
rect 2228 7055 2362 7071
rect 2228 7021 2244 7055
rect 2278 7021 2312 7055
rect 2346 7021 2362 7055
rect 2228 7005 2362 7021
rect 360 5879 460 5921
rect 2228 5879 2328 5921
rect 326 5863 460 5879
rect 326 5829 342 5863
rect 376 5829 410 5863
rect 444 5829 460 5863
rect 326 5813 460 5829
rect 516 5807 1316 5879
rect 1372 5807 2172 5879
rect 2228 5863 2362 5879
rect 2228 5829 2244 5863
rect 2278 5829 2312 5863
rect 2346 5829 2362 5863
rect 2228 5813 2362 5829
rect 360 4687 460 4729
rect 2228 4687 2328 4729
rect 326 4671 460 4687
rect 326 4637 342 4671
rect 376 4637 410 4671
rect 444 4637 460 4671
rect 326 4621 460 4637
rect 516 4615 1316 4687
rect 1372 4615 2172 4687
rect 2228 4671 2362 4687
rect 2228 4637 2244 4671
rect 2278 4637 2312 4671
rect 2346 4637 2362 4671
rect 2228 4621 2362 4637
rect 360 3495 460 3537
rect 2228 3495 2328 3537
rect 326 3479 460 3495
rect 326 3445 342 3479
rect 376 3445 410 3479
rect 444 3445 460 3479
rect 326 3429 460 3445
rect 516 3423 1316 3495
rect 1372 3423 2172 3495
rect 2228 3479 2362 3495
rect 2228 3445 2244 3479
rect 2278 3445 2312 3479
rect 2346 3445 2362 3479
rect 2228 3429 2362 3445
rect 904 2048 1004 2064
rect 904 2014 937 2048
rect 971 2014 1004 2048
rect 904 1980 1004 2014
rect 904 1950 937 1980
rect 921 1946 937 1950
rect 971 1950 1004 1980
rect 1060 2048 1160 2064
rect 1060 2014 1093 2048
rect 1127 2014 1160 2048
rect 1060 1980 1160 2014
rect 1060 1950 1093 1980
rect 971 1946 987 1950
rect 921 1930 987 1946
rect 1077 1946 1093 1950
rect 1127 1950 1160 1980
rect 1216 2048 1316 2064
rect 1216 2014 1249 2048
rect 1283 2014 1316 2048
rect 1216 1980 1316 2014
rect 1216 1950 1249 1980
rect 1127 1946 1143 1950
rect 1077 1930 1143 1946
rect 1233 1946 1249 1950
rect 1283 1950 1316 1980
rect 1372 2048 1472 2064
rect 1372 2014 1405 2048
rect 1439 2014 1472 2048
rect 1372 1980 1472 2014
rect 1372 1950 1405 1980
rect 1283 1946 1299 1950
rect 1233 1930 1299 1946
rect 1389 1946 1405 1950
rect 1439 1950 1472 1980
rect 1528 2048 1628 2064
rect 1528 2014 1561 2048
rect 1595 2014 1628 2048
rect 1528 1980 1628 2014
rect 1528 1950 1561 1980
rect 1439 1946 1455 1950
rect 1389 1930 1455 1946
rect 1545 1946 1561 1950
rect 1595 1950 1628 1980
rect 1684 2048 1784 2064
rect 1684 2014 1717 2048
rect 1751 2014 1784 2048
rect 1684 1980 1784 2014
rect 1684 1950 1717 1980
rect 1595 1946 1611 1950
rect 1545 1930 1611 1946
rect 1701 1946 1717 1950
rect 1751 1950 1784 1980
rect 1751 1946 1767 1950
rect 1701 1930 1767 1946
rect 163 530 263 543
rect 319 530 419 543
rect 475 530 575 543
rect 2113 530 2213 543
rect 2269 530 2369 543
rect 2425 530 2525 543
rect 163 80 197 146
rect 1283 80 1316 146
rect 1372 80 1405 146
rect 2491 80 2525 146
<< polycont >>
rect 349 8688 383 8722
rect 417 8688 451 8722
rect 605 8688 639 8722
rect 673 8688 707 8722
rect 861 8688 895 8722
rect 929 8688 963 8722
rect 1117 8688 1151 8722
rect 1185 8688 1219 8722
rect 1373 8688 1407 8722
rect 1441 8688 1475 8722
rect 1629 8688 1663 8722
rect 1697 8688 1731 8722
rect 1885 8688 1919 8722
rect 1953 8688 1987 8722
rect 2141 8688 2175 8722
rect 2209 8688 2243 8722
rect 342 7021 376 7055
rect 410 7021 444 7055
rect 2244 7021 2278 7055
rect 2312 7021 2346 7055
rect 342 5829 376 5863
rect 410 5829 444 5863
rect 2244 5829 2278 5863
rect 2312 5829 2346 5863
rect 342 4637 376 4671
rect 410 4637 444 4671
rect 2244 4637 2278 4671
rect 2312 4637 2346 4671
rect 342 3445 376 3479
rect 410 3445 444 3479
rect 2244 3445 2278 3479
rect 2312 3445 2346 3479
rect 937 2014 971 2048
rect 937 1946 971 1980
rect 1093 2014 1127 2048
rect 1093 1946 1127 1980
rect 1249 2014 1283 2048
rect 1249 1946 1283 1980
rect 1405 2014 1439 2048
rect 1405 1946 1439 1980
rect 1561 2014 1595 2048
rect 1561 1946 1595 1980
rect 1717 2014 1751 2048
rect 1717 1946 1751 1980
<< locali >>
rect 1357 8722 1491 8772
rect 333 8688 349 8722
rect 407 8688 417 8722
rect 485 8688 529 8722
rect 563 8688 605 8722
rect 641 8688 673 8722
rect 719 8688 763 8722
rect 797 8688 841 8722
rect 895 8688 919 8722
rect 963 8688 997 8722
rect 1031 8688 1075 8722
rect 1109 8688 1117 8722
rect 1151 8688 1153 8722
rect 1219 8688 1230 8722
rect 1357 8688 1373 8722
rect 1407 8688 1441 8722
rect 1475 8688 1491 8722
rect 1617 8688 1629 8722
rect 1696 8688 1697 8722
rect 1731 8688 1741 8722
rect 1775 8688 1820 8722
rect 1854 8688 1885 8722
rect 1933 8688 1953 8722
rect 2012 8688 2057 8722
rect 2091 8688 2135 8722
rect 2175 8688 2209 8722
rect 2247 8688 2259 8722
rect 55 7540 2680 7541
rect 55 7506 89 7540
rect 123 7506 157 7540
rect 191 7506 225 7540
rect 259 7506 293 7540
rect 327 7506 361 7540
rect 395 7506 429 7540
rect 463 7506 497 7540
rect 531 7506 565 7540
rect 599 7506 633 7540
rect 667 7506 701 7540
rect 735 7506 769 7540
rect 803 7506 837 7540
rect 871 7506 905 7540
rect 939 7506 973 7540
rect 1007 7506 1041 7540
rect 1075 7506 1109 7540
rect 1143 7506 1177 7540
rect 1211 7506 1245 7540
rect 1279 7506 1313 7540
rect 1347 7506 1381 7540
rect 1415 7506 1449 7540
rect 1483 7506 1517 7540
rect 1551 7506 1585 7540
rect 1619 7506 1653 7540
rect 1687 7506 1721 7540
rect 1755 7506 1789 7540
rect 1823 7506 1857 7540
rect 1891 7506 1925 7540
rect 1959 7506 1993 7540
rect 2027 7506 2061 7540
rect 2095 7506 2129 7540
rect 2163 7506 2197 7540
rect 2231 7506 2265 7540
rect 2299 7506 2333 7540
rect 2367 7506 2401 7540
rect 2435 7506 2469 7540
rect 2503 7506 2537 7540
rect 2571 7506 2605 7540
rect 2639 7506 2680 7540
rect 55 7505 2680 7506
rect 8 7351 2680 7352
rect 8 7317 85 7351
rect 119 7317 187 7351
rect 221 7317 255 7351
rect 289 7317 323 7351
rect 357 7317 391 7351
rect 425 7317 459 7351
rect 493 7317 527 7351
rect 561 7317 595 7351
rect 629 7317 663 7351
rect 697 7317 731 7351
rect 765 7317 799 7351
rect 833 7317 867 7351
rect 901 7317 935 7351
rect 969 7317 1003 7351
rect 1037 7317 1071 7351
rect 1105 7317 1139 7351
rect 1173 7317 1207 7351
rect 1241 7317 1275 7351
rect 1309 7317 1343 7351
rect 1377 7317 1411 7351
rect 1445 7317 1479 7351
rect 1513 7317 1547 7351
rect 1581 7317 1615 7351
rect 1649 7317 1683 7351
rect 1717 7317 1751 7351
rect 1785 7317 1819 7351
rect 1853 7317 1887 7351
rect 1921 7317 1955 7351
rect 1989 7317 2023 7351
rect 2057 7317 2091 7351
rect 2125 7317 2159 7351
rect 2193 7317 2227 7351
rect 2261 7317 2295 7351
rect 2329 7317 2363 7351
rect 2397 7317 2431 7351
rect 2465 7317 2499 7351
rect 2533 7317 2567 7351
rect 2601 7317 2680 7351
rect 8 7316 2680 7317
rect 8 7256 44 7316
rect 8 7222 9 7256
rect 43 7222 44 7256
rect 8 7188 44 7222
rect 8 7154 9 7188
rect 43 7154 44 7188
rect 8 7120 44 7154
rect 2644 7282 2680 7316
rect 2644 7248 2645 7282
rect 2679 7248 2680 7282
rect 2644 7214 2680 7248
rect 2644 7180 2645 7214
rect 2679 7180 2680 7214
rect 2644 7146 2680 7180
rect 8 7086 9 7120
rect 43 7086 44 7120
rect 8 7052 44 7086
rect 8 7018 9 7052
rect 43 7018 44 7052
rect 8 6984 44 7018
rect 8 6950 9 6984
rect 43 6950 44 6984
rect 8 6916 44 6950
rect 8 6882 9 6916
rect 43 6882 44 6916
rect 8 6848 44 6882
rect 8 6814 9 6848
rect 43 6814 44 6848
rect 8 6780 44 6814
rect 8 6746 9 6780
rect 43 6746 44 6780
rect 8 6712 44 6746
rect 8 6678 9 6712
rect 43 6678 44 6712
rect 8 6644 44 6678
rect 8 6610 9 6644
rect 43 6610 44 6644
rect 8 6576 44 6610
rect 8 6542 9 6576
rect 43 6542 44 6576
rect 8 6508 44 6542
rect 8 6474 9 6508
rect 43 6474 44 6508
rect 8 6440 44 6474
rect 8 6406 9 6440
rect 43 6406 44 6440
rect 8 6372 44 6406
rect 8 6338 9 6372
rect 43 6338 44 6372
rect 8 6304 44 6338
rect 8 6270 9 6304
rect 43 6270 44 6304
rect 8 6236 44 6270
rect 8 6202 9 6236
rect 43 6202 44 6236
rect 8 6168 44 6202
rect 8 6134 9 6168
rect 43 6134 44 6168
rect 8 6100 44 6134
rect 8 6066 9 6100
rect 43 6066 44 6100
rect 8 6032 44 6066
rect 8 5998 9 6032
rect 43 5998 44 6032
rect 8 5964 44 5998
rect 8 5930 9 5964
rect 43 5930 44 5964
rect 8 5896 44 5930
rect 8 5862 9 5896
rect 43 5862 44 5896
rect 8 5828 44 5862
rect 8 5794 9 5828
rect 43 5794 44 5828
rect 8 5760 44 5794
rect 8 5726 9 5760
rect 43 5726 44 5760
rect 8 5692 44 5726
rect 8 5658 9 5692
rect 43 5658 44 5692
rect 8 5624 44 5658
rect 8 5590 9 5624
rect 43 5590 44 5624
rect 8 5556 44 5590
rect 8 5522 9 5556
rect 43 5522 44 5556
rect 8 5488 44 5522
rect 8 5454 9 5488
rect 43 5454 44 5488
rect 8 5420 44 5454
rect 8 5386 9 5420
rect 43 5386 44 5420
rect 8 5352 44 5386
rect 8 5318 9 5352
rect 43 5318 44 5352
rect 8 5284 44 5318
rect 8 5250 9 5284
rect 43 5250 44 5284
rect 8 5216 44 5250
rect 8 5182 9 5216
rect 43 5182 44 5216
rect 8 5148 44 5182
rect 8 5114 9 5148
rect 43 5114 44 5148
rect 8 5080 44 5114
rect 8 5046 9 5080
rect 43 5046 44 5080
rect 8 5012 44 5046
rect 8 4978 9 5012
rect 43 4978 44 5012
rect 8 4944 44 4978
rect 8 4910 9 4944
rect 43 4910 44 4944
rect 8 4876 44 4910
rect 8 4842 9 4876
rect 43 4842 44 4876
rect 8 4808 44 4842
rect 8 4774 9 4808
rect 43 4774 44 4808
rect 8 4740 44 4774
rect 8 4706 9 4740
rect 43 4706 44 4740
rect 8 4672 44 4706
rect 8 4638 9 4672
rect 43 4638 44 4672
rect 8 4604 44 4638
rect 8 4570 9 4604
rect 43 4570 44 4604
rect 8 4536 44 4570
rect 8 4502 9 4536
rect 43 4502 44 4536
rect 8 4468 44 4502
rect 8 4434 9 4468
rect 43 4434 44 4468
rect 8 4400 44 4434
rect 8 4366 9 4400
rect 43 4366 44 4400
rect 8 4332 44 4366
rect 8 4298 9 4332
rect 43 4298 44 4332
rect 8 4264 44 4298
rect 8 4230 9 4264
rect 43 4230 44 4264
rect 8 4196 44 4230
rect 8 4162 9 4196
rect 43 4162 44 4196
rect 8 4128 44 4162
rect 8 4094 9 4128
rect 43 4094 44 4128
rect 8 4060 44 4094
rect 8 4026 9 4060
rect 43 4026 44 4060
rect 8 3992 44 4026
rect 8 3958 9 3992
rect 43 3958 44 3992
rect 8 3924 44 3958
rect 8 3890 9 3924
rect 43 3890 44 3924
rect 8 3856 44 3890
rect 8 3822 9 3856
rect 43 3822 44 3856
rect 8 3788 44 3822
rect 8 3754 9 3788
rect 43 3754 44 3788
rect 8 3720 44 3754
rect 8 3686 9 3720
rect 43 3686 44 3720
rect 8 3652 44 3686
rect 8 3618 9 3652
rect 43 3618 44 3652
rect 8 3584 44 3618
rect 8 3550 9 3584
rect 43 3550 44 3584
rect 8 3516 44 3550
rect 8 3482 9 3516
rect 43 3482 44 3516
rect 8 3448 44 3482
rect 8 3414 9 3448
rect 43 3414 44 3448
rect 8 3380 44 3414
rect 8 3346 9 3380
rect 43 3346 44 3380
rect 8 3312 44 3346
rect 8 3278 9 3312
rect 43 3278 44 3312
rect 8 3244 44 3278
rect 8 3210 9 3244
rect 43 3210 44 3244
rect 8 3176 44 3210
rect 8 3142 9 3176
rect 43 3142 44 3176
rect 8 3108 44 3142
rect 8 3074 9 3108
rect 43 3074 44 3108
rect 8 3040 44 3074
rect 8 3006 9 3040
rect 43 3006 44 3040
rect 8 2972 44 3006
rect 8 2938 9 2972
rect 43 2938 44 2972
rect 8 2904 44 2938
rect 8 2870 9 2904
rect 43 2870 44 2904
rect 8 2836 44 2870
rect 8 2802 9 2836
rect 43 2802 44 2836
rect 8 2768 44 2802
rect 8 2734 9 2768
rect 43 2734 44 2768
rect 8 2700 44 2734
rect 8 2666 9 2700
rect 43 2666 44 2700
rect 8 2632 44 2666
rect 8 2598 9 2632
rect 43 2598 44 2632
rect 8 2564 44 2598
rect 8 2530 9 2564
rect 43 2530 44 2564
rect 8 2496 44 2530
rect 8 2462 9 2496
rect 43 2462 44 2496
rect 8 2428 44 2462
rect 8 2394 9 2428
rect 43 2394 44 2428
rect 8 2360 44 2394
rect 8 2326 9 2360
rect 43 2326 44 2360
rect 8 2292 44 2326
rect 8 2258 9 2292
rect 43 2258 44 2292
rect 197 7140 2491 7141
rect 197 7106 231 7140
rect 265 7106 299 7140
rect 333 7106 367 7140
rect 401 7106 435 7140
rect 469 7106 503 7140
rect 537 7106 571 7140
rect 605 7106 639 7140
rect 673 7106 707 7140
rect 741 7106 775 7140
rect 809 7106 843 7140
rect 877 7106 911 7140
rect 945 7106 979 7140
rect 1013 7106 1047 7140
rect 1081 7106 1115 7140
rect 1149 7106 1183 7140
rect 1217 7106 1251 7140
rect 1285 7106 1319 7140
rect 1353 7106 1387 7140
rect 1421 7106 1455 7140
rect 1489 7106 1523 7140
rect 1557 7106 1591 7140
rect 1625 7106 1659 7140
rect 1693 7106 1727 7140
rect 1761 7106 1795 7140
rect 1829 7106 1863 7140
rect 1897 7106 1931 7140
rect 1965 7106 1999 7140
rect 2033 7106 2067 7140
rect 2101 7106 2135 7140
rect 2169 7106 2203 7140
rect 2237 7106 2271 7140
rect 2305 7106 2339 7140
rect 2373 7107 2491 7140
rect 2373 7106 2456 7107
rect 197 7105 2456 7106
rect 197 7047 233 7105
rect 2455 7073 2456 7105
rect 2490 7073 2491 7107
rect 197 7013 198 7047
rect 232 7013 233 7047
rect 294 7055 444 7071
rect 294 7035 342 7055
rect 197 6979 233 7013
rect 197 6945 198 6979
rect 232 6945 233 6979
rect 197 6911 233 6945
rect 315 7021 342 7035
rect 376 7021 410 7055
rect 315 7005 444 7021
rect 2244 7055 2394 7071
rect 2278 7021 2312 7055
rect 2346 7035 2394 7055
rect 2455 7039 2491 7073
rect 2346 7021 2373 7035
rect 2244 7005 2373 7021
rect 315 6919 349 7005
rect 2339 6919 2373 7005
rect 2455 7005 2456 7039
rect 2490 7005 2491 7039
rect 2455 6971 2491 7005
rect 2455 6937 2456 6971
rect 2490 6937 2491 6971
rect 197 6877 198 6911
rect 232 6877 233 6911
rect 197 6843 233 6877
rect 197 6809 198 6843
rect 232 6809 233 6843
rect 197 6775 233 6809
rect 197 6741 198 6775
rect 232 6741 233 6775
rect 197 6707 233 6741
rect 197 6673 198 6707
rect 232 6673 233 6707
rect 197 6639 233 6673
rect 197 6605 198 6639
rect 232 6605 233 6639
rect 197 6571 233 6605
rect 197 6537 198 6571
rect 232 6537 233 6571
rect 197 6503 233 6537
rect 197 6469 198 6503
rect 232 6469 233 6503
rect 197 6435 233 6469
rect 197 6401 198 6435
rect 232 6401 233 6435
rect 197 6367 233 6401
rect 197 6333 198 6367
rect 232 6333 233 6367
rect 197 6299 233 6333
rect 197 6265 198 6299
rect 232 6265 233 6299
rect 197 6231 233 6265
rect 197 6197 198 6231
rect 232 6197 233 6231
rect 197 6163 233 6197
rect 197 6129 198 6163
rect 232 6129 233 6163
rect 197 6095 233 6129
rect 197 6061 198 6095
rect 232 6061 233 6095
rect 197 6027 233 6061
rect 197 5993 198 6027
rect 232 5993 233 6027
rect 197 5959 233 5993
rect 2455 6903 2491 6937
rect 2455 6869 2456 6903
rect 2490 6869 2491 6903
rect 2455 6835 2491 6869
rect 2455 6801 2456 6835
rect 2490 6801 2491 6835
rect 2455 6767 2491 6801
rect 2455 6733 2456 6767
rect 2490 6733 2491 6767
rect 2455 6699 2491 6733
rect 2455 6665 2456 6699
rect 2490 6665 2491 6699
rect 2455 6631 2491 6665
rect 2455 6597 2456 6631
rect 2490 6597 2491 6631
rect 2455 6563 2491 6597
rect 2455 6529 2456 6563
rect 2490 6529 2491 6563
rect 2455 6495 2491 6529
rect 2455 6461 2456 6495
rect 2490 6461 2491 6495
rect 2455 6427 2491 6461
rect 2455 6393 2456 6427
rect 2490 6393 2491 6427
rect 2455 6359 2491 6393
rect 2455 6325 2456 6359
rect 2490 6325 2491 6359
rect 2455 6291 2491 6325
rect 2455 6257 2456 6291
rect 2490 6257 2491 6291
rect 2455 6223 2491 6257
rect 2455 6189 2456 6223
rect 2490 6189 2491 6223
rect 2455 6155 2491 6189
rect 2455 6121 2456 6155
rect 2490 6121 2491 6155
rect 2455 6087 2491 6121
rect 2455 6053 2456 6087
rect 2490 6053 2491 6087
rect 2455 6019 2491 6053
rect 2455 5985 2456 6019
rect 2490 5985 2491 6019
rect 197 5925 198 5959
rect 232 5925 233 5959
rect 197 5891 233 5925
rect 197 5857 198 5891
rect 232 5857 233 5891
rect 197 5823 233 5857
rect 197 5789 198 5823
rect 232 5789 233 5823
rect 197 5755 233 5789
rect 197 5721 198 5755
rect 232 5721 233 5755
rect 315 5879 349 5969
rect 2339 5879 2373 5969
rect 315 5863 444 5879
rect 315 5829 342 5863
rect 376 5829 410 5863
rect 315 5813 444 5829
rect 2244 5863 2373 5879
rect 2278 5829 2312 5863
rect 2346 5829 2373 5863
rect 2244 5813 2373 5829
rect 315 5727 349 5813
rect 2339 5727 2373 5813
rect 2455 5951 2491 5985
rect 2455 5917 2456 5951
rect 2490 5917 2491 5951
rect 2455 5883 2491 5917
rect 2455 5849 2456 5883
rect 2490 5849 2491 5883
rect 2455 5815 2491 5849
rect 2455 5781 2456 5815
rect 2490 5781 2491 5815
rect 2455 5747 2491 5781
rect 197 5687 233 5721
rect 197 5653 198 5687
rect 232 5653 233 5687
rect 197 5619 233 5653
rect 197 5585 198 5619
rect 232 5585 233 5619
rect 197 5551 233 5585
rect 197 5517 198 5551
rect 232 5517 233 5551
rect 197 5483 233 5517
rect 197 5449 198 5483
rect 232 5449 233 5483
rect 197 5415 233 5449
rect 197 5381 198 5415
rect 232 5381 233 5415
rect 197 5347 233 5381
rect 197 5313 198 5347
rect 232 5313 233 5347
rect 197 5279 233 5313
rect 197 5245 198 5279
rect 232 5245 233 5279
rect 197 5211 233 5245
rect 197 5177 198 5211
rect 232 5177 233 5211
rect 197 5143 233 5177
rect 197 5109 198 5143
rect 232 5109 233 5143
rect 197 5075 233 5109
rect 197 5041 198 5075
rect 232 5041 233 5075
rect 197 5007 233 5041
rect 197 4973 198 5007
rect 232 4973 233 5007
rect 197 4939 233 4973
rect 197 4905 198 4939
rect 232 4905 233 4939
rect 197 4871 233 4905
rect 197 4837 198 4871
rect 232 4837 233 4871
rect 197 4803 233 4837
rect 197 4769 198 4803
rect 232 4769 233 4803
rect 2455 5713 2456 5747
rect 2490 5713 2491 5747
rect 2455 5679 2491 5713
rect 2455 5645 2456 5679
rect 2490 5645 2491 5679
rect 2455 5611 2491 5645
rect 2455 5577 2456 5611
rect 2490 5577 2491 5611
rect 2455 5543 2491 5577
rect 2455 5509 2456 5543
rect 2490 5509 2491 5543
rect 2455 5475 2491 5509
rect 2455 5441 2456 5475
rect 2490 5441 2491 5475
rect 2455 5407 2491 5441
rect 2455 5373 2456 5407
rect 2490 5373 2491 5407
rect 2455 5339 2491 5373
rect 2455 5305 2456 5339
rect 2490 5305 2491 5339
rect 2455 5271 2491 5305
rect 2455 5237 2456 5271
rect 2490 5237 2491 5271
rect 2455 5203 2491 5237
rect 2455 5169 2456 5203
rect 2490 5169 2491 5203
rect 2455 5135 2491 5169
rect 2455 5101 2456 5135
rect 2490 5101 2491 5135
rect 2455 5067 2491 5101
rect 2455 5033 2456 5067
rect 2490 5033 2491 5067
rect 2455 4999 2491 5033
rect 2455 4965 2456 4999
rect 2490 4965 2491 4999
rect 2455 4931 2491 4965
rect 2455 4897 2456 4931
rect 2490 4897 2491 4931
rect 2455 4863 2491 4897
rect 2455 4829 2456 4863
rect 2490 4829 2491 4863
rect 2455 4795 2491 4829
rect 197 4735 233 4769
rect 197 4701 198 4735
rect 232 4701 233 4735
rect 197 4667 233 4701
rect 197 4633 198 4667
rect 232 4633 233 4667
rect 197 4599 233 4633
rect 197 4565 198 4599
rect 232 4565 233 4599
rect 197 4531 233 4565
rect 315 4687 349 4777
rect 2339 4687 2373 4777
rect 315 4671 444 4687
rect 315 4637 342 4671
rect 376 4637 410 4671
rect 315 4621 444 4637
rect 2244 4671 2373 4687
rect 2278 4637 2312 4671
rect 2346 4637 2373 4671
rect 2244 4621 2373 4637
rect 315 4535 349 4621
rect 2339 4535 2373 4621
rect 2455 4761 2456 4795
rect 2490 4761 2491 4795
rect 2455 4727 2491 4761
rect 2455 4693 2456 4727
rect 2490 4693 2491 4727
rect 2455 4659 2491 4693
rect 2455 4625 2456 4659
rect 2490 4625 2491 4659
rect 2455 4591 2491 4625
rect 2455 4557 2456 4591
rect 2490 4557 2491 4591
rect 197 4497 198 4531
rect 232 4497 233 4531
rect 197 4463 233 4497
rect 197 4429 198 4463
rect 232 4429 233 4463
rect 197 4395 233 4429
rect 197 4361 198 4395
rect 232 4361 233 4395
rect 197 4327 233 4361
rect 197 4293 198 4327
rect 232 4293 233 4327
rect 197 4259 233 4293
rect 197 4225 198 4259
rect 232 4225 233 4259
rect 197 4191 233 4225
rect 197 4157 198 4191
rect 232 4157 233 4191
rect 197 4123 233 4157
rect 197 4089 198 4123
rect 232 4089 233 4123
rect 197 4055 233 4089
rect 197 4021 198 4055
rect 232 4021 233 4055
rect 197 3987 233 4021
rect 197 3953 198 3987
rect 232 3953 233 3987
rect 197 3919 233 3953
rect 197 3885 198 3919
rect 232 3885 233 3919
rect 197 3851 233 3885
rect 197 3817 198 3851
rect 232 3817 233 3851
rect 197 3783 233 3817
rect 197 3749 198 3783
rect 232 3749 233 3783
rect 197 3715 233 3749
rect 197 3681 198 3715
rect 232 3681 233 3715
rect 197 3647 233 3681
rect 197 3613 198 3647
rect 232 3613 233 3647
rect 197 3579 233 3613
rect 2455 4523 2491 4557
rect 2455 4489 2456 4523
rect 2490 4489 2491 4523
rect 2455 4455 2491 4489
rect 2455 4421 2456 4455
rect 2490 4421 2491 4455
rect 2455 4387 2491 4421
rect 2455 4353 2456 4387
rect 2490 4353 2491 4387
rect 2455 4319 2491 4353
rect 2455 4285 2456 4319
rect 2490 4285 2491 4319
rect 2455 4251 2491 4285
rect 2455 4217 2456 4251
rect 2490 4217 2491 4251
rect 2455 4183 2491 4217
rect 2455 4149 2456 4183
rect 2490 4149 2491 4183
rect 2455 4115 2491 4149
rect 2455 4081 2456 4115
rect 2490 4081 2491 4115
rect 2455 4047 2491 4081
rect 2455 4013 2456 4047
rect 2490 4013 2491 4047
rect 2455 3979 2491 4013
rect 2455 3945 2456 3979
rect 2490 3945 2491 3979
rect 2455 3911 2491 3945
rect 2455 3877 2456 3911
rect 2490 3877 2491 3911
rect 2455 3843 2491 3877
rect 2455 3809 2456 3843
rect 2490 3809 2491 3843
rect 2455 3775 2491 3809
rect 2455 3741 2456 3775
rect 2490 3741 2491 3775
rect 2455 3707 2491 3741
rect 2455 3673 2456 3707
rect 2490 3673 2491 3707
rect 2455 3639 2491 3673
rect 2455 3605 2456 3639
rect 2490 3605 2491 3639
rect 197 3545 198 3579
rect 232 3545 233 3579
rect 197 3511 233 3545
rect 197 3477 198 3511
rect 232 3477 233 3511
rect 197 3443 233 3477
rect 197 3409 198 3443
rect 232 3409 233 3443
rect 197 3375 233 3409
rect 197 3341 198 3375
rect 232 3341 233 3375
rect 315 3495 349 3585
rect 2339 3495 2373 3585
rect 315 3479 444 3495
rect 315 3445 342 3479
rect 376 3445 410 3479
rect 315 3429 444 3445
rect 2244 3479 2373 3495
rect 2278 3445 2312 3479
rect 2346 3445 2373 3479
rect 2244 3429 2373 3445
rect 315 3343 349 3429
rect 2339 3343 2373 3429
rect 2455 3571 2491 3605
rect 2455 3537 2456 3571
rect 2490 3537 2491 3571
rect 2455 3503 2491 3537
rect 2455 3469 2456 3503
rect 2490 3469 2491 3503
rect 2455 3435 2491 3469
rect 2455 3401 2456 3435
rect 2490 3401 2491 3435
rect 2455 3367 2491 3401
rect 197 3307 233 3341
rect 197 3273 198 3307
rect 232 3273 233 3307
rect 197 3239 233 3273
rect 197 3205 198 3239
rect 232 3205 233 3239
rect 197 3171 233 3205
rect 197 3137 198 3171
rect 232 3137 233 3171
rect 197 3103 233 3137
rect 197 3069 198 3103
rect 232 3069 233 3103
rect 197 3035 233 3069
rect 197 3001 198 3035
rect 232 3001 233 3035
rect 197 2967 233 3001
rect 197 2933 198 2967
rect 232 2933 233 2967
rect 197 2899 233 2933
rect 197 2865 198 2899
rect 232 2865 233 2899
rect 197 2831 233 2865
rect 197 2797 198 2831
rect 232 2797 233 2831
rect 197 2763 233 2797
rect 197 2729 198 2763
rect 232 2729 233 2763
rect 197 2695 233 2729
rect 197 2661 198 2695
rect 232 2661 233 2695
rect 197 2627 233 2661
rect 197 2593 198 2627
rect 232 2593 233 2627
rect 197 2559 233 2593
rect 197 2525 198 2559
rect 232 2525 233 2559
rect 197 2491 233 2525
rect 197 2457 198 2491
rect 232 2457 233 2491
rect 197 2423 233 2457
rect 197 2389 198 2423
rect 232 2389 233 2423
rect 197 2355 233 2389
rect 197 2321 198 2355
rect 232 2323 233 2355
rect 2455 3333 2456 3367
rect 2490 3333 2491 3367
rect 2455 3299 2491 3333
rect 2455 3265 2456 3299
rect 2490 3265 2491 3299
rect 2455 3231 2491 3265
rect 2455 3197 2456 3231
rect 2490 3197 2491 3231
rect 2455 3163 2491 3197
rect 2455 3129 2456 3163
rect 2490 3129 2491 3163
rect 2455 3095 2491 3129
rect 2455 3061 2456 3095
rect 2490 3061 2491 3095
rect 2455 3027 2491 3061
rect 2455 2993 2456 3027
rect 2490 2993 2491 3027
rect 2455 2959 2491 2993
rect 2455 2925 2456 2959
rect 2490 2925 2491 2959
rect 2455 2891 2491 2925
rect 2455 2857 2456 2891
rect 2490 2857 2491 2891
rect 2455 2823 2491 2857
rect 2455 2789 2456 2823
rect 2490 2789 2491 2823
rect 2455 2755 2491 2789
rect 2455 2721 2456 2755
rect 2490 2721 2491 2755
rect 2455 2687 2491 2721
rect 2455 2653 2456 2687
rect 2490 2653 2491 2687
rect 2455 2619 2491 2653
rect 2455 2585 2456 2619
rect 2490 2585 2491 2619
rect 2455 2551 2491 2585
rect 2455 2517 2456 2551
rect 2490 2517 2491 2551
rect 2455 2483 2491 2517
rect 2455 2449 2456 2483
rect 2490 2449 2491 2483
rect 2455 2323 2491 2449
rect 232 2322 2491 2323
rect 232 2321 315 2322
rect 197 2288 315 2321
rect 349 2288 383 2322
rect 417 2288 451 2322
rect 485 2288 519 2322
rect 553 2288 587 2322
rect 621 2288 655 2322
rect 689 2288 723 2322
rect 757 2288 791 2322
rect 825 2288 859 2322
rect 893 2288 927 2322
rect 961 2288 995 2322
rect 1029 2288 1063 2322
rect 1097 2288 1131 2322
rect 1165 2288 1199 2322
rect 1233 2288 1267 2322
rect 1301 2288 1335 2322
rect 1369 2288 1403 2322
rect 1437 2288 1471 2322
rect 1505 2288 1539 2322
rect 1573 2288 1607 2322
rect 1641 2288 1675 2322
rect 1709 2288 1743 2322
rect 1777 2288 1811 2322
rect 1845 2288 1879 2322
rect 1913 2288 1947 2322
rect 1981 2288 2015 2322
rect 2049 2288 2083 2322
rect 2117 2288 2151 2322
rect 2185 2288 2219 2322
rect 2253 2288 2271 2322
rect 2321 2288 2343 2322
rect 2389 2288 2423 2322
rect 2457 2288 2491 2322
rect 197 2287 2491 2288
rect 2644 7112 2645 7146
rect 2679 7112 2680 7146
rect 2644 7078 2680 7112
rect 2644 7044 2645 7078
rect 2679 7044 2680 7078
rect 2644 7010 2680 7044
rect 2644 6976 2645 7010
rect 2679 6976 2680 7010
rect 2644 6942 2680 6976
rect 2644 6908 2645 6942
rect 2679 6908 2680 6942
rect 2644 6874 2680 6908
rect 2644 6840 2645 6874
rect 2679 6840 2680 6874
rect 2644 6806 2680 6840
rect 2644 6772 2645 6806
rect 2679 6772 2680 6806
rect 2644 6738 2680 6772
rect 2644 6704 2645 6738
rect 2679 6704 2680 6738
rect 2644 6670 2680 6704
rect 2644 6636 2645 6670
rect 2679 6636 2680 6670
rect 2644 6602 2680 6636
rect 2644 6568 2645 6602
rect 2679 6568 2680 6602
rect 2644 6534 2680 6568
rect 2644 6500 2645 6534
rect 2679 6500 2680 6534
rect 2644 6466 2680 6500
rect 2644 6432 2645 6466
rect 2679 6432 2680 6466
rect 2644 6398 2680 6432
rect 2644 6364 2645 6398
rect 2679 6364 2680 6398
rect 2644 6330 2680 6364
rect 2644 6296 2645 6330
rect 2679 6296 2680 6330
rect 2644 6262 2680 6296
rect 2644 6228 2645 6262
rect 2679 6228 2680 6262
rect 2644 6194 2680 6228
rect 2644 6160 2645 6194
rect 2679 6160 2680 6194
rect 2644 6126 2680 6160
rect 2644 6092 2645 6126
rect 2679 6092 2680 6126
rect 2644 6058 2680 6092
rect 2644 6024 2645 6058
rect 2679 6024 2680 6058
rect 2644 5990 2680 6024
rect 2644 5956 2645 5990
rect 2679 5956 2680 5990
rect 2644 5922 2680 5956
rect 2644 5888 2645 5922
rect 2679 5888 2680 5922
rect 2644 5854 2680 5888
rect 2644 5820 2645 5854
rect 2679 5820 2680 5854
rect 2644 5786 2680 5820
rect 2644 5752 2645 5786
rect 2679 5752 2680 5786
rect 2644 5718 2680 5752
rect 2644 5684 2645 5718
rect 2679 5684 2680 5718
rect 2644 5650 2680 5684
rect 2644 5616 2645 5650
rect 2679 5616 2680 5650
rect 2644 5582 2680 5616
rect 2644 5548 2645 5582
rect 2679 5548 2680 5582
rect 2644 5514 2680 5548
rect 2644 5480 2645 5514
rect 2679 5480 2680 5514
rect 2644 5446 2680 5480
rect 2644 5412 2645 5446
rect 2679 5412 2680 5446
rect 2644 5378 2680 5412
rect 2644 5344 2645 5378
rect 2679 5344 2680 5378
rect 2644 5310 2680 5344
rect 2644 5276 2645 5310
rect 2679 5276 2680 5310
rect 2644 5242 2680 5276
rect 2644 5208 2645 5242
rect 2679 5208 2680 5242
rect 2644 5174 2680 5208
rect 2644 5140 2645 5174
rect 2679 5140 2680 5174
rect 2644 5106 2680 5140
rect 2644 5072 2645 5106
rect 2679 5072 2680 5106
rect 2644 5038 2680 5072
rect 2644 5004 2645 5038
rect 2679 5004 2680 5038
rect 2644 4970 2680 5004
rect 2644 4936 2645 4970
rect 2679 4936 2680 4970
rect 2644 4902 2680 4936
rect 2644 4868 2645 4902
rect 2679 4868 2680 4902
rect 2644 4834 2680 4868
rect 2644 4800 2645 4834
rect 2679 4800 2680 4834
rect 2644 4766 2680 4800
rect 2644 4732 2645 4766
rect 2679 4732 2680 4766
rect 2644 4698 2680 4732
rect 2644 4664 2645 4698
rect 2679 4664 2680 4698
rect 2644 4630 2680 4664
rect 2644 4596 2645 4630
rect 2679 4596 2680 4630
rect 2644 4562 2680 4596
rect 2644 4528 2645 4562
rect 2679 4528 2680 4562
rect 2644 4494 2680 4528
rect 2644 4460 2645 4494
rect 2679 4460 2680 4494
rect 2644 4426 2680 4460
rect 2644 4392 2645 4426
rect 2679 4392 2680 4426
rect 2644 4358 2680 4392
rect 2644 4324 2645 4358
rect 2679 4324 2680 4358
rect 2644 4290 2680 4324
rect 2644 4256 2645 4290
rect 2679 4256 2680 4290
rect 2644 4222 2680 4256
rect 2644 4188 2645 4222
rect 2679 4188 2680 4222
rect 2644 4154 2680 4188
rect 2644 4120 2645 4154
rect 2679 4120 2680 4154
rect 2644 4086 2680 4120
rect 2644 4052 2645 4086
rect 2679 4052 2680 4086
rect 2644 4018 2680 4052
rect 2644 3984 2645 4018
rect 2679 3984 2680 4018
rect 2644 3950 2680 3984
rect 2644 3916 2645 3950
rect 2679 3916 2680 3950
rect 2644 3882 2680 3916
rect 2644 3848 2645 3882
rect 2679 3848 2680 3882
rect 2644 3814 2680 3848
rect 2644 3780 2645 3814
rect 2679 3780 2680 3814
rect 2644 3746 2680 3780
rect 2644 3712 2645 3746
rect 2679 3712 2680 3746
rect 2644 3678 2680 3712
rect 2644 3644 2645 3678
rect 2679 3644 2680 3678
rect 2644 3610 2680 3644
rect 2644 3576 2645 3610
rect 2679 3576 2680 3610
rect 2644 3542 2680 3576
rect 2644 3508 2645 3542
rect 2679 3508 2680 3542
rect 2644 3474 2680 3508
rect 2644 3440 2645 3474
rect 2679 3440 2680 3474
rect 2644 3406 2680 3440
rect 2644 3372 2645 3406
rect 2679 3372 2680 3406
rect 2644 3338 2680 3372
rect 2644 3304 2645 3338
rect 2679 3304 2680 3338
rect 2644 3270 2680 3304
rect 2644 3236 2645 3270
rect 2679 3236 2680 3270
rect 2644 3202 2680 3236
rect 2644 3168 2645 3202
rect 2679 3168 2680 3202
rect 2644 3134 2680 3168
rect 2644 3100 2645 3134
rect 2679 3100 2680 3134
rect 2644 3066 2680 3100
rect 2644 3032 2645 3066
rect 2679 3032 2680 3066
rect 2644 2998 2680 3032
rect 2644 2964 2645 2998
rect 2679 2964 2680 2998
rect 2644 2930 2680 2964
rect 2644 2896 2645 2930
rect 2679 2896 2680 2930
rect 2644 2862 2680 2896
rect 2644 2828 2645 2862
rect 2679 2828 2680 2862
rect 2644 2794 2680 2828
rect 2644 2760 2645 2794
rect 2679 2760 2680 2794
rect 2644 2726 2680 2760
rect 2644 2692 2645 2726
rect 2679 2692 2680 2726
rect 2644 2658 2680 2692
rect 2644 2624 2645 2658
rect 2679 2624 2680 2658
rect 2644 2590 2680 2624
rect 2644 2556 2645 2590
rect 2679 2556 2680 2590
rect 2644 2522 2680 2556
rect 2644 2488 2645 2522
rect 2679 2488 2680 2522
rect 2644 2454 2680 2488
rect 2644 2420 2645 2454
rect 2679 2420 2680 2454
rect 2644 2386 2680 2420
rect 2644 2352 2645 2386
rect 2679 2352 2680 2386
rect 2644 2318 2680 2352
rect 8 2224 44 2258
rect 8 2190 9 2224
rect 43 2190 44 2224
rect 8 2156 44 2190
rect 8 2122 9 2156
rect 43 2134 44 2156
rect 2644 2284 2645 2318
rect 2679 2284 2680 2318
rect 2644 2250 2680 2284
rect 2644 2216 2645 2250
rect 2679 2216 2680 2250
rect 2644 2182 2680 2216
rect 2644 2148 2645 2182
rect 2679 2148 2680 2182
rect 2644 2134 2680 2148
rect 43 2133 2680 2134
rect 43 2122 96 2133
rect 8 2099 96 2122
rect 162 2099 168 2133
rect 230 2099 240 2133
rect 298 2099 312 2133
rect 366 2099 384 2133
rect 434 2099 456 2133
rect 502 2099 536 2133
rect 570 2099 604 2133
rect 638 2099 672 2133
rect 706 2099 740 2133
rect 774 2099 808 2133
rect 842 2099 876 2133
rect 910 2099 944 2133
rect 978 2099 1012 2133
rect 1046 2099 1080 2133
rect 1114 2099 1148 2133
rect 1182 2099 1216 2133
rect 1250 2099 1284 2133
rect 1318 2099 1352 2133
rect 1386 2099 1420 2133
rect 1454 2099 1488 2133
rect 1522 2099 1556 2133
rect 1590 2099 1624 2133
rect 1658 2099 1692 2133
rect 1726 2099 1760 2133
rect 1794 2099 1828 2133
rect 1862 2099 1896 2133
rect 1930 2099 1964 2133
rect 1998 2099 2032 2133
rect 2066 2099 2100 2133
rect 2134 2099 2168 2133
rect 2202 2099 2236 2133
rect 2270 2099 2304 2133
rect 2338 2099 2372 2133
rect 2406 2099 2440 2133
rect 2474 2099 2508 2133
rect 2542 2099 2576 2133
rect 2610 2114 2680 2133
rect 2610 2099 2645 2114
rect 8 2098 2645 2099
rect 8 2088 44 2098
rect 8 2054 9 2088
rect 43 2054 44 2088
rect 8 2020 44 2054
rect 2644 2080 2645 2098
rect 2679 2080 2680 2114
rect 8 1986 9 2020
rect 43 1986 44 2020
rect 8 1952 44 1986
rect 859 2014 937 2048
rect 971 2014 987 2048
rect 859 1980 987 2014
rect 8 1918 9 1952
rect 43 1918 44 1952
rect 8 1884 44 1918
rect 8 1850 9 1884
rect 43 1850 44 1884
rect 8 1816 44 1850
rect 8 1782 9 1816
rect 43 1782 44 1816
rect 8 1748 44 1782
rect 8 1714 9 1748
rect 43 1714 44 1748
rect 8 1680 44 1714
rect 8 1646 9 1680
rect 43 1646 44 1680
rect 8 1612 44 1646
rect 8 1578 9 1612
rect 43 1578 44 1612
rect 8 1544 44 1578
rect 8 1510 9 1544
rect 43 1510 44 1544
rect 8 1476 44 1510
rect 8 1442 9 1476
rect 43 1442 44 1476
rect 8 1408 44 1442
rect 8 1374 9 1408
rect 43 1374 44 1408
rect 8 1340 44 1374
rect 8 1306 9 1340
rect 43 1306 44 1340
rect 8 1272 44 1306
rect 8 1238 9 1272
rect 43 1238 44 1272
rect 8 1204 44 1238
rect 8 1170 9 1204
rect 43 1170 44 1204
rect 8 1136 44 1170
rect 8 1102 9 1136
rect 43 1102 44 1136
rect 8 1068 44 1102
rect 8 1034 9 1068
rect 43 1034 44 1068
rect 8 1000 44 1034
rect 8 966 9 1000
rect 43 966 44 1000
rect 8 932 44 966
rect 8 898 9 932
rect 43 898 44 932
rect 8 864 44 898
rect 8 830 9 864
rect 43 830 44 864
rect 8 796 44 830
rect 8 762 9 796
rect 43 762 44 796
rect 8 728 44 762
rect 8 694 9 728
rect 43 694 44 728
rect 8 660 44 694
rect 8 626 9 660
rect 43 626 44 660
rect 8 592 44 626
rect 8 558 9 592
rect 43 558 44 592
rect 8 524 44 558
rect 8 490 9 524
rect 43 490 44 524
rect 8 329 44 490
rect 118 444 152 591
rect 8 295 9 329
rect 43 295 44 329
rect 8 261 44 295
rect 8 227 9 261
rect 43 227 44 261
rect 8 193 44 227
rect 8 159 9 193
rect 43 159 44 193
rect 216 174 366 1975
rect 859 1946 937 1980
rect 971 1946 987 1980
rect 1077 2004 1093 2048
rect 1127 2004 1143 2048
rect 1077 1980 1143 2004
rect 1077 1946 1093 1980
rect 1127 1946 1143 1980
rect 1233 2004 1249 2048
rect 1283 2004 1299 2048
rect 1233 1980 1299 2004
rect 1233 1946 1249 1980
rect 1283 1946 1299 1980
rect 1389 2004 1405 2048
rect 1439 2004 1455 2048
rect 1389 1980 1455 2004
rect 1389 1946 1405 1980
rect 1439 1946 1455 1980
rect 1545 2004 1561 2048
rect 1595 2004 1611 2048
rect 1545 1980 1611 2004
rect 1545 1946 1561 1980
rect 1595 1946 1611 1980
rect 1701 2014 1717 2048
rect 1751 2014 1829 2048
rect 1701 1980 1829 2014
rect 1701 1946 1717 1980
rect 1751 1946 1829 1980
rect 2644 2046 2680 2080
rect 2644 2012 2645 2046
rect 2679 2012 2680 2046
rect 2644 1978 2680 2012
rect 859 1884 893 1946
rect 859 1812 893 1850
rect 1795 1884 1829 1946
rect 1015 1767 1049 1805
rect 1015 1695 1049 1733
rect 1327 1767 1361 1805
rect 1171 1637 1205 1675
rect 1327 1695 1361 1733
rect 1639 1767 1673 1805
rect 1795 1812 1829 1850
rect 1327 1623 1361 1661
rect 1483 1637 1517 1675
rect 1639 1695 1673 1733
rect 430 444 464 591
rect 586 174 737 1471
rect 859 382 893 434
rect 957 174 1107 1471
rect 1171 382 1205 434
rect 1269 174 1419 1471
rect 1483 382 1517 434
rect 1581 174 1731 1471
rect 1795 382 1829 434
rect 1951 174 2102 1471
rect 2224 444 2258 591
rect 2322 174 2472 1975
rect 2644 1944 2645 1978
rect 2679 1944 2680 1978
rect 2644 1910 2680 1944
rect 2644 1876 2645 1910
rect 2679 1876 2680 1910
rect 2644 1842 2680 1876
rect 2644 1808 2645 1842
rect 2679 1808 2680 1842
rect 2644 1774 2680 1808
rect 2644 1740 2645 1774
rect 2679 1740 2680 1774
rect 2644 1706 2680 1740
rect 2644 1672 2645 1706
rect 2679 1672 2680 1706
rect 2644 1638 2680 1672
rect 2644 1604 2645 1638
rect 2679 1604 2680 1638
rect 2644 1570 2680 1604
rect 2644 1536 2645 1570
rect 2679 1536 2680 1570
rect 2644 1502 2680 1536
rect 2644 1468 2645 1502
rect 2679 1468 2680 1502
rect 2644 1434 2680 1468
rect 2644 1400 2645 1434
rect 2679 1400 2680 1434
rect 2644 1366 2680 1400
rect 2644 1332 2645 1366
rect 2679 1332 2680 1366
rect 2644 1298 2680 1332
rect 2644 1264 2645 1298
rect 2679 1264 2680 1298
rect 2644 1230 2680 1264
rect 2644 1196 2645 1230
rect 2679 1196 2680 1230
rect 2644 1162 2680 1196
rect 2644 1128 2645 1162
rect 2679 1128 2680 1162
rect 2644 1094 2680 1128
rect 2644 1060 2645 1094
rect 2679 1060 2680 1094
rect 2644 1026 2680 1060
rect 2644 992 2645 1026
rect 2679 992 2680 1026
rect 2644 958 2680 992
rect 2644 924 2645 958
rect 2679 924 2680 958
rect 2644 890 2680 924
rect 2644 856 2645 890
rect 2679 856 2680 890
rect 2644 822 2680 856
rect 2644 788 2645 822
rect 2679 788 2680 822
rect 2644 754 2680 788
rect 2644 720 2645 754
rect 2679 720 2680 754
rect 2644 686 2680 720
rect 2644 652 2645 686
rect 2679 652 2680 686
rect 2644 618 2680 652
rect 2536 444 2570 591
rect 2644 584 2645 618
rect 2679 584 2680 618
rect 2644 550 2680 584
rect 2644 516 2645 550
rect 2679 516 2680 550
rect 2644 482 2680 516
rect 2644 448 2645 482
rect 2679 448 2680 482
rect 2644 414 2680 448
rect 2644 380 2645 414
rect 2679 380 2680 414
rect 2644 346 2680 380
rect 2644 312 2645 346
rect 2679 312 2680 346
rect 2644 278 2680 312
rect 2644 244 2645 278
rect 2679 244 2680 278
rect 2644 210 2680 244
rect 2644 176 2645 210
rect 2679 176 2680 210
rect 8 125 44 159
rect 2644 142 2680 176
rect 8 91 9 125
rect 43 91 44 125
rect 672 96 710 130
rect 2407 96 2445 130
rect 2644 108 2645 142
rect 2679 108 2680 142
rect 8 57 44 91
rect 2644 57 2680 108
<< viali >>
rect 373 8688 383 8722
rect 383 8688 407 8722
rect 451 8688 485 8722
rect 529 8688 563 8722
rect 607 8688 639 8722
rect 639 8688 641 8722
rect 685 8688 707 8722
rect 707 8688 719 8722
rect 763 8688 797 8722
rect 841 8688 861 8722
rect 861 8688 875 8722
rect 919 8688 929 8722
rect 929 8688 953 8722
rect 997 8688 1031 8722
rect 1075 8688 1109 8722
rect 1153 8688 1185 8722
rect 1185 8688 1187 8722
rect 1230 8688 1264 8722
rect 1583 8688 1617 8722
rect 1662 8688 1663 8722
rect 1663 8688 1696 8722
rect 1741 8688 1775 8722
rect 1820 8688 1854 8722
rect 1899 8688 1919 8722
rect 1919 8688 1933 8722
rect 1978 8688 1987 8722
rect 1987 8688 2012 8722
rect 2057 8688 2091 8722
rect 2135 8688 2141 8722
rect 2141 8688 2169 8722
rect 2213 8688 2243 8722
rect 2243 8688 2247 8722
rect 2271 2288 2287 2322
rect 2287 2288 2305 2322
rect 2343 2288 2355 2322
rect 2355 2288 2377 2322
rect 96 2099 128 2133
rect 128 2099 130 2133
rect 168 2099 196 2133
rect 196 2099 202 2133
rect 240 2099 264 2133
rect 264 2099 274 2133
rect 312 2099 332 2133
rect 332 2099 346 2133
rect 384 2099 400 2133
rect 400 2099 418 2133
rect 456 2099 468 2133
rect 468 2099 490 2133
rect 1093 2014 1127 2038
rect 1093 2004 1127 2014
rect 1093 1946 1127 1966
rect 1249 2014 1283 2038
rect 1249 2004 1283 2014
rect 1249 1946 1283 1966
rect 1405 2014 1439 2038
rect 1405 2004 1439 2014
rect 1405 1946 1439 1966
rect 1561 2014 1595 2038
rect 1561 2004 1595 2014
rect 1561 1946 1595 1966
rect 1093 1932 1127 1946
rect 1249 1932 1283 1946
rect 1405 1932 1439 1946
rect 1561 1932 1595 1946
rect 859 1850 893 1884
rect 1795 1850 1829 1884
rect 859 1778 893 1812
rect 1015 1805 1049 1839
rect 1015 1733 1049 1767
rect 1327 1805 1361 1839
rect 1327 1733 1361 1767
rect 1015 1661 1049 1695
rect 1171 1675 1205 1709
rect 1171 1603 1205 1637
rect 1639 1805 1673 1839
rect 1795 1778 1829 1812
rect 1639 1733 1673 1767
rect 1327 1661 1361 1695
rect 1327 1589 1361 1623
rect 1483 1675 1517 1709
rect 1639 1661 1673 1695
rect 1483 1603 1517 1637
rect 638 96 672 130
rect 710 96 744 130
rect 2373 96 2407 130
rect 2445 96 2479 130
<< metal1 >>
rect 291 8722 2259 8728
rect 291 8688 373 8722
rect 407 8688 451 8722
rect 485 8688 529 8722
rect 563 8688 607 8722
rect 641 8688 685 8722
rect 719 8688 763 8722
rect 797 8688 841 8722
rect 875 8688 919 8722
rect 953 8688 997 8722
rect 1031 8688 1075 8722
rect 1109 8688 1153 8722
rect 1187 8688 1230 8722
rect 1264 8688 1583 8722
rect 1617 8688 1662 8722
rect 1696 8688 1741 8722
rect 1775 8688 1820 8722
rect 1854 8688 1899 8722
rect 1933 8688 1978 8722
rect 2012 8688 2057 8722
rect 2091 8688 2135 8722
rect 2169 8688 2213 8722
rect 2247 8688 2259 8722
rect 291 8682 2259 8688
rect 243 8620 2405 8626
rect 243 8568 567 8620
rect 619 8568 2405 8620
rect 243 8556 2405 8568
rect 243 8504 567 8556
rect 619 8504 2405 8556
rect 243 8492 2405 8504
rect 243 8440 567 8492
rect 619 8440 2405 8492
rect 243 8434 2405 8440
rect 243 8399 301 8434
tri 301 8409 326 8434 nw
tri 730 8409 755 8434 ne
tri 813 8409 838 8434 nw
tri 1242 8409 1267 8434 ne
tri 1325 8409 1350 8434 nw
tri 1754 8409 1779 8434 ne
tri 1837 8409 1862 8434 nw
tri 2266 8409 2291 8434 ne
rect 2291 8399 2349 8434
tri 2349 8409 2374 8434 nw
rect 499 7750 557 7802
rect 500 7748 556 7749
rect 1011 7750 1069 7802
rect 1012 7748 1068 7749
rect 500 7711 556 7712
rect 1012 7711 1068 7712
rect 499 7685 557 7710
tri 557 7685 582 7710 sw
tri 986 7685 1011 7710 se
rect 1011 7685 1069 7710
tri 1069 7685 1094 7710 sw
tri 1498 7685 1523 7710 se
rect 1523 7685 1581 7796
rect 2035 7750 2093 7802
rect 2036 7748 2092 7749
rect 2036 7711 2092 7712
tri 1581 7685 1606 7710 sw
tri 2010 7685 2035 7710 se
rect 2035 7685 2093 7710
rect 499 7658 2093 7685
tri 499 7633 524 7658 ne
rect 524 7633 2068 7658
tri 2068 7633 2093 7658 nw
tri 1290 7608 1315 7633 ne
rect 10 7538 1187 7546
rect 10 7422 43 7538
rect 223 7422 308 7538
rect 488 7486 567 7538
rect 619 7486 1187 7538
rect 488 7474 1187 7486
rect 488 7422 567 7474
rect 619 7422 1187 7474
rect 10 7413 1187 7422
rect -3 7305 107 7357
rect 159 7305 171 7357
rect 223 7305 229 7357
tri 229 7305 235 7311 nw
rect -3 7264 55 7305
tri 55 7271 89 7305 nw
tri 186 7120 212 7146 se
rect 212 7120 293 7146
rect 186 7113 293 7120
rect 244 7100 293 7113
rect 186 2378 337 7100
tri 337 7075 362 7100 nw
rect 1113 7061 1165 7067
tri 1087 6983 1113 7009 ne
rect 1113 6997 1165 7009
tri 1165 6983 1191 7009 nw
rect 1113 6939 1165 6945
rect 465 5937 511 5957
tri 511 5937 531 5957 sw
tri 465 5901 501 5937 ne
rect 501 5901 531 5937
tri 531 5901 567 5937 sw
tri 501 5875 527 5901 ne
rect 527 5875 567 5901
tri 567 5875 593 5901 sw
tri 527 5835 567 5875 ne
rect 567 5855 593 5875
tri 593 5855 613 5875 sw
tri 445 4745 511 4811 se
tri 383 4683 445 4745 se
rect 445 4683 449 4745
tri 449 4683 511 4745 nw
tri 561 4683 567 4689 se
rect 567 4683 613 5855
rect 1221 5869 1273 5875
tri 1195 5791 1221 5817 ne
rect 1221 5805 1273 5817
rect 1221 5747 1273 5753
rect 1005 5620 1273 5626
rect 1057 5568 1221 5620
rect 1005 5556 1273 5568
rect 1057 5504 1221 5556
rect 1005 5498 1273 5504
tri 379 4679 383 4683 se
rect 383 4679 445 4683
tri 445 4679 449 4683 nw
tri 557 4679 561 4683 se
rect 561 4679 613 4683
rect 379 3461 425 4679
tri 425 4659 445 4679 nw
tri 537 4659 557 4679 se
rect 557 4669 613 4679
rect 557 4659 597 4669
tri 531 4653 537 4659 se
rect 537 4653 597 4659
tri 597 4653 613 4669 nw
rect 1113 4677 1165 4683
tri 465 4587 531 4653 se
rect 531 4623 567 4653
tri 567 4623 597 4653 nw
tri 1087 4623 1089 4625 ne
rect 1089 4623 1165 4625
tri 531 4587 567 4623 nw
tri 1089 4599 1113 4623 ne
rect 1113 4613 1165 4623
rect 465 4567 511 4587
tri 511 4567 531 4587 nw
tri 1165 4599 1191 4625 nw
rect 1113 4555 1165 4561
rect 1005 3804 1273 3810
rect 1057 3752 1221 3804
rect 1005 3740 1273 3752
rect 1057 3688 1221 3740
rect 1005 3682 1273 3688
rect 465 3553 511 3573
tri 465 3507 511 3553 ne
tri 511 3507 577 3573 sw
tri 511 3481 537 3507 ne
rect 537 3491 577 3507
tri 577 3491 593 3507 sw
rect 537 3481 593 3491
tri 593 3481 603 3491 sw
rect 1221 3485 1273 3491
tri 379 3415 425 3461 ne
tri 425 3415 491 3481 sw
tri 537 3471 547 3481 ne
rect 547 3471 603 3481
tri 603 3471 613 3481 sw
tri 547 3451 567 3471 ne
tri 425 3395 445 3415 ne
rect 445 3395 491 3415
tri 491 3395 511 3415 sw
tri 445 3363 477 3395 ne
rect 477 3363 511 3395
tri 477 3329 511 3363 ne
rect 567 2455 613 3471
tri 1195 3407 1221 3433 ne
rect 1221 3421 1273 3433
rect 1221 3363 1273 3369
tri 613 2455 619 2461 sw
rect 567 2449 619 2455
tri 241 2288 257 2304 se
rect 257 2298 309 2304
tri 175 2222 241 2288 se
rect 241 2246 257 2288
rect 241 2234 309 2246
rect 241 2222 257 2234
rect 70 2182 257 2222
rect 465 2254 511 2389
rect 567 2385 619 2397
rect 1315 2381 1373 7633
tri 1373 7608 1398 7633 nw
tri 2266 7546 2291 7571 se
rect 2291 7546 2349 7633
tri 2349 7546 2374 7571 sw
rect 1429 7538 2403 7546
rect 1429 7422 2200 7538
rect 2380 7422 2403 7538
rect 1429 7413 2403 7422
tri 2453 7305 2459 7311 ne
rect 2459 7305 2465 7357
rect 2517 7305 2529 7357
rect 2581 7305 2691 7357
tri 2598 7270 2633 7305 ne
rect 2633 7265 2691 7305
rect 2395 7120 2476 7146
tri 2476 7120 2502 7146 sw
rect 2395 7113 2502 7120
rect 2395 7100 2444 7113
tri 2326 7075 2351 7100 ne
rect 1523 7061 1575 7067
tri 1497 6983 1523 7009 ne
rect 1523 6997 1575 7009
tri 1575 6983 1601 7009 nw
rect 1523 6939 1575 6945
rect 2351 6209 2502 7100
tri 2165 5945 2177 5957 se
rect 2177 5945 2223 5957
rect 1415 5939 1467 5945
tri 2141 5921 2165 5945 se
rect 2165 5937 2223 5945
rect 2165 5921 2207 5937
tri 2207 5921 2223 5937 nw
tri 2121 5901 2141 5921 se
rect 2141 5901 2177 5921
rect 1415 5875 1467 5887
tri 1467 5875 1493 5901 sw
tri 2095 5875 2121 5901 se
rect 2121 5891 2177 5901
tri 2177 5891 2207 5921 nw
rect 2121 5875 2141 5891
rect 1415 5817 1467 5823
tri 2075 5855 2095 5875 se
rect 2095 5855 2141 5875
tri 2141 5855 2177 5891 nw
rect 1415 5620 1683 5626
rect 1467 5568 1631 5620
rect 1415 5556 1683 5568
rect 1467 5504 1631 5556
rect 1415 5498 1683 5504
rect 2075 4683 2121 5855
tri 2121 5835 2141 5855 nw
tri 2177 4745 2243 4811 sw
tri 2177 4725 2197 4745 ne
rect 2197 4725 2243 4745
tri 2243 4725 2263 4745 sw
tri 2197 4689 2233 4725 ne
rect 2233 4689 2263 4725
tri 2121 4683 2127 4689 sw
tri 2233 4683 2239 4689 ne
rect 2239 4683 2263 4689
rect 1523 4677 1575 4683
rect 2075 4669 2127 4683
tri 2075 4625 2119 4669 ne
rect 2119 4625 2127 4669
tri 2127 4625 2185 4683 sw
tri 2239 4659 2263 4683 ne
tri 2263 4679 2309 4725 sw
tri 1497 4599 1523 4625 ne
rect 1523 4613 1575 4625
tri 1575 4599 1601 4625 nw
tri 2119 4623 2121 4625 ne
rect 2121 4623 2185 4625
tri 2185 4623 2187 4625 sw
tri 2121 4599 2145 4623 ne
rect 2145 4599 2187 4623
tri 2187 4599 2211 4623 sw
tri 2145 4587 2157 4599 ne
rect 2157 4587 2211 4599
tri 2211 4587 2223 4599 sw
tri 2157 4567 2177 4587 ne
rect 2177 4567 2223 4587
rect 1523 4555 1575 4561
rect 1415 3804 1683 3810
rect 1467 3752 1631 3804
rect 1415 3740 1683 3752
rect 1467 3688 1631 3740
rect 1415 3682 1683 3688
tri 2165 3561 2177 3573 se
rect 2177 3561 2223 3573
rect 1415 3555 1467 3561
tri 2141 3537 2165 3561 se
rect 2165 3553 2223 3561
rect 2165 3537 2207 3553
tri 2207 3537 2223 3553 nw
tri 2121 3517 2141 3537 se
rect 2141 3517 2177 3537
rect 1415 3491 1467 3503
tri 1467 3491 1493 3517 sw
tri 2095 3491 2121 3517 se
rect 2121 3507 2177 3517
tri 2177 3507 2207 3537 nw
rect 2121 3491 2141 3507
rect 1415 3433 1467 3439
tri 2075 3471 2095 3491 se
rect 2095 3471 2141 3491
tri 2141 3471 2177 3507 nw
tri 2253 3471 2263 3481 se
rect 2263 3471 2309 4679
tri 2069 2455 2075 2461 se
rect 2075 2455 2121 3471
tri 2121 3451 2141 3471 nw
tri 2243 3461 2253 3471 se
rect 2253 3461 2309 3471
tri 2233 3451 2243 3461 se
tri 2177 3395 2233 3451 se
rect 2233 3395 2243 3451
tri 2243 3395 2309 3461 nw
tri 2177 3329 2243 3395 nw
rect 2069 2449 2121 2455
rect 2069 2385 2121 2397
rect 567 2327 619 2333
tri 1274 2328 1280 2334 se
rect 1280 2328 1286 2334
rect 1229 2282 1286 2328
rect 1338 2282 1350 2334
rect 1402 2328 1408 2334
tri 1408 2328 1414 2334 sw
rect 1402 2282 1459 2328
tri 511 2254 536 2279 sw
tri 2044 2254 2069 2279 se
rect 2069 2254 2121 2333
rect 465 2251 2121 2254
tri 465 2225 491 2251 ne
rect 491 2225 2095 2251
tri 2095 2225 2121 2251 nw
tri 2150 2196 2177 2223 se
rect 2177 2203 2223 2389
tri 2326 2328 2351 2353 se
rect 2351 2328 2502 6039
rect 2259 2322 2444 2328
rect 2259 2288 2271 2322
rect 2305 2288 2343 2322
rect 2377 2315 2444 2322
rect 2377 2308 2502 2315
rect 2377 2288 2476 2308
rect 2259 2282 2476 2288
tri 2476 2282 2502 2308 nw
rect 2177 2196 2216 2203
tri 2216 2196 2223 2203 nw
tri 2663 2196 2691 2224 se
tri 591 2194 593 2196 se
rect 593 2194 2214 2196
tri 2214 2194 2216 2196 nw
tri 2661 2194 2663 2196 se
rect 2663 2194 2691 2196
rect 70 2176 309 2182
tri 573 2176 591 2194 se
rect 591 2176 2187 2194
tri 567 2170 573 2176 se
rect 573 2170 2187 2176
rect 567 2167 2187 2170
tri 2187 2167 2214 2194 nw
tri 2634 2167 2661 2194 se
rect 2661 2167 2691 2194
rect 567 2142 620 2167
tri 620 2142 645 2167 nw
tri 1062 2142 1087 2167 ne
rect -3 2133 502 2139
rect -3 2099 96 2133
rect 130 2099 168 2133
rect 202 2099 240 2133
rect 274 2099 312 2133
rect 346 2099 384 2133
rect 418 2099 456 2133
rect 490 2099 502 2133
rect -3 1884 502 2099
rect 567 2059 619 2142
tri 619 2141 620 2142 nw
rect 567 1995 619 2007
rect 1087 2038 1133 2167
tri 1133 2142 1158 2167 nw
tri 1218 2142 1243 2167 ne
rect 1243 2142 1289 2167
tri 1289 2142 1314 2167 nw
tri 1374 2142 1399 2167 ne
rect 1244 2140 1288 2141
rect 1087 2004 1093 2038
rect 1127 2004 1133 2038
rect 1087 1966 1133 2004
tri 619 1945 625 1951 sw
rect 619 1943 625 1945
rect 567 1937 625 1943
tri 625 1937 633 1945 sw
tri 567 1932 572 1937 ne
rect 572 1932 633 1937
tri 633 1932 638 1937 sw
rect 1087 1932 1093 1966
rect 1127 1932 1133 1966
tri 572 1905 599 1932 ne
rect 599 1920 638 1932
tri 638 1920 650 1932 sw
rect 1087 1920 1133 1932
rect 1244 2103 1288 2104
rect 1243 2038 1289 2102
rect 1243 2004 1249 2038
rect 1283 2004 1289 2038
rect 1243 1966 1289 2004
rect 1243 1932 1249 1966
rect 1283 1932 1289 1966
rect 1243 1920 1289 1932
rect 1399 2038 1445 2167
tri 1445 2142 1470 2167 nw
tri 1530 2142 1555 2167 ne
rect 1555 2142 1601 2167
tri 1601 2142 1626 2167 nw
tri 2609 2142 2634 2167 se
rect 2634 2142 2691 2167
tri 2608 2141 2609 2142 se
rect 2609 2141 2691 2142
rect 1556 2140 1600 2141
tri 2607 2140 2608 2141 se
rect 2608 2140 2691 2141
tri 2606 2139 2607 2140 se
rect 2607 2139 2691 2140
rect 1399 2004 1405 2038
rect 1439 2004 1445 2038
rect 1399 1966 1445 2004
rect 1399 1932 1405 1966
rect 1439 1932 1445 1966
rect 1399 1920 1445 1932
rect 1556 2103 1600 2104
rect 1555 2038 1601 2102
tri 2161 2068 2186 2093 ne
rect 1555 2004 1561 2038
rect 1595 2004 1601 2038
rect 1555 1966 1601 2004
rect 1555 1932 1561 1966
rect 1595 1932 1601 1966
rect 2069 2059 2121 2065
rect 2069 1995 2121 2007
tri 2055 1937 2069 1951 se
rect 2069 1937 2121 1943
rect 1555 1920 1601 1932
tri 2038 1920 2055 1937 se
rect 2055 1920 2089 1937
rect 599 1905 650 1920
tri 502 1884 523 1905 sw
tri 599 1884 620 1905 ne
rect 620 1896 650 1905
tri 650 1896 674 1920 sw
rect 1244 1918 1288 1919
rect 620 1884 674 1896
tri 674 1884 686 1896 sw
rect 853 1884 899 1896
tri 899 1884 911 1896 sw
rect -3 1879 523 1884
tri 523 1879 528 1884 sw
tri 620 1879 625 1884 ne
rect 625 1879 686 1884
tri 686 1879 691 1884 sw
rect -3 1850 528 1879
tri 528 1850 557 1879 sw
tri 625 1850 654 1879 ne
rect 654 1850 691 1879
tri 691 1850 720 1879 sw
rect 853 1850 859 1884
rect 893 1876 911 1884
tri 911 1876 919 1884 sw
rect 1243 1882 1289 1918
rect 1244 1881 1288 1882
rect 893 1851 919 1876
tri 919 1851 944 1876 sw
tri 1218 1851 1243 1876 se
rect 1243 1851 1289 1880
tri 2037 1919 2038 1920 se
rect 2038 1919 2089 1920
rect 1556 1918 1600 1919
tri 2036 1918 2037 1919 se
rect 2037 1918 2089 1919
rect 1555 1882 1601 1918
tri 2023 1905 2036 1918 se
rect 2036 1905 2089 1918
tri 2089 1905 2121 1937 nw
tri 2014 1896 2023 1905 se
rect 2023 1896 2069 1905
tri 1777 1884 1789 1896 se
rect 1789 1884 1835 1896
tri 2003 1885 2014 1896 se
rect 2014 1885 2069 1896
tri 2069 1885 2089 1905 nw
tri 2166 1885 2186 1905 se
rect 2186 1885 2691 2139
tri 1775 1882 1777 1884 se
rect 1777 1882 1795 1884
rect 1556 1881 1600 1882
tri 1774 1881 1775 1882 se
rect 1775 1881 1795 1882
tri 1773 1880 1774 1881 se
rect 1774 1880 1795 1881
tri 1289 1851 1314 1876 sw
tri 1530 1851 1555 1876 se
rect 1555 1851 1601 1880
tri 1769 1876 1773 1880 se
rect 1773 1876 1795 1880
tri 1601 1851 1626 1876 sw
tri 1744 1851 1769 1876 se
rect 1769 1851 1795 1876
rect 893 1850 1795 1851
rect 1829 1850 1835 1884
rect -3 1839 557 1850
tri 557 1839 568 1850 sw
tri 654 1839 665 1850 ne
rect 665 1839 720 1850
tri 720 1839 731 1850 sw
rect 853 1839 1835 1850
rect -3 1827 568 1839
tri 568 1827 580 1839 sw
tri 665 1827 677 1839 ne
rect 677 1827 731 1839
tri 731 1827 743 1839 sw
rect -3 1813 580 1827
tri 580 1813 594 1827 sw
tri 677 1813 691 1827 ne
rect 691 1813 743 1827
tri 743 1813 757 1827 sw
rect -3 1812 594 1813
tri 594 1812 595 1813 sw
tri 691 1812 692 1813 ne
rect 692 1812 757 1813
tri 757 1812 758 1813 sw
rect 853 1812 1015 1839
rect -3 1778 595 1812
tri 595 1778 629 1812 sw
tri 692 1778 726 1812 ne
rect 726 1778 758 1812
tri 758 1778 792 1812 sw
rect 853 1778 859 1812
rect 893 1805 1015 1812
rect 1049 1805 1327 1839
rect 1361 1805 1639 1839
rect 1673 1812 1835 1839
tri 1937 1819 2003 1885 se
tri 2003 1819 2069 1885 nw
tri 2100 1819 2166 1885 se
rect 2166 1819 2691 1885
rect 1673 1805 1795 1812
rect 893 1778 1795 1805
rect 1829 1778 1835 1812
rect -3 1767 629 1778
tri 629 1767 640 1778 sw
tri 726 1767 737 1778 ne
rect 737 1767 792 1778
tri 792 1767 803 1778 sw
rect 853 1767 1835 1778
rect -3 1747 640 1767
tri 640 1747 660 1767 sw
tri 737 1747 757 1767 ne
rect 757 1766 803 1767
tri 803 1766 804 1767 sw
rect 853 1766 1015 1767
rect 757 1747 804 1766
tri 804 1747 823 1766 sw
tri 853 1747 872 1766 ne
rect 872 1747 1015 1766
rect -3 1733 660 1747
tri 660 1733 674 1747 sw
tri 757 1733 771 1747 ne
rect 771 1733 823 1747
tri 823 1733 837 1747 sw
tri 872 1733 886 1747 ne
rect 886 1733 1015 1747
rect 1049 1749 1327 1767
rect 1049 1733 1064 1749
tri 1064 1733 1080 1749 nw
tri 1225 1733 1241 1749 ne
rect 1241 1733 1327 1749
rect 1361 1749 1639 1767
rect 1361 1733 1447 1749
tri 1447 1733 1463 1749 nw
tri 1608 1733 1624 1749 ne
rect 1624 1733 1639 1749
rect 1673 1766 1835 1767
tri 1884 1766 1937 1819 se
rect 1673 1753 1822 1766
tri 1822 1753 1835 1766 nw
tri 1871 1753 1884 1766 se
rect 1884 1753 1937 1766
tri 1937 1753 2003 1819 nw
tri 2034 1753 2100 1819 se
rect 2100 1753 2691 1819
rect 1673 1749 1818 1753
tri 1818 1749 1822 1753 nw
tri 1867 1749 1871 1753 se
rect 1673 1733 1786 1749
rect -3 1709 674 1733
tri 674 1709 698 1733 sw
tri 771 1709 795 1733 ne
rect 795 1717 837 1733
tri 837 1717 853 1733 sw
tri 886 1717 902 1733 ne
rect 902 1717 1055 1733
tri 1055 1724 1064 1733 nw
tri 1241 1724 1250 1733 ne
rect 795 1709 853 1717
tri 853 1709 861 1717 sw
tri 902 1709 910 1717 ne
rect 910 1709 1055 1717
rect -3 1695 698 1709
tri 698 1695 712 1709 sw
tri 795 1695 809 1709 ne
rect 809 1695 861 1709
tri 861 1695 875 1709 sw
tri 910 1695 924 1709 ne
rect 924 1695 1055 1709
rect -3 1681 712 1695
tri 712 1681 726 1695 sw
tri 809 1681 823 1695 ne
rect 823 1681 875 1695
tri 875 1681 889 1695 sw
tri 924 1681 938 1695 ne
rect 938 1681 1015 1695
rect -3 1661 726 1681
tri 726 1661 746 1681 sw
tri 823 1661 843 1681 ne
rect 843 1666 889 1681
tri 889 1666 904 1681 sw
tri 938 1666 953 1681 ne
rect 953 1666 1015 1681
rect 843 1661 904 1666
tri 904 1661 909 1666 sw
tri 953 1661 958 1666 ne
rect 958 1661 1015 1666
rect 1049 1661 1055 1695
rect -3 1637 56 1661
tri 56 1637 80 1661 nw
tri 243 1637 267 1661 ne
rect 267 1637 315 1661
tri 315 1637 339 1661 nw
tri 427 1637 451 1661 ne
rect 451 1637 746 1661
tri 746 1637 770 1661 sw
tri 843 1651 853 1661 ne
rect 853 1651 909 1661
tri 853 1649 855 1651 ne
rect 855 1649 909 1651
tri 909 1649 921 1661 sw
tri 958 1649 970 1661 ne
rect 970 1649 1055 1661
rect 1165 1709 1211 1721
rect 1165 1675 1171 1709
rect 1205 1675 1211 1709
tri 855 1637 867 1649 ne
rect 867 1640 921 1649
tri 921 1640 930 1649 sw
rect 867 1637 930 1640
tri 930 1637 933 1640 sw
tri 1162 1637 1165 1640 se
rect 1165 1637 1211 1675
rect -3 522 55 1637
tri 55 1636 56 1637 nw
tri 267 1636 268 1637 ne
rect 268 1636 314 1637
tri 314 1636 315 1637 nw
tri 451 1636 452 1637 ne
rect 452 1636 770 1637
tri 452 1603 485 1636 ne
rect 485 1615 770 1636
tri 770 1615 792 1637 sw
tri 867 1615 889 1637 ne
rect 889 1615 933 1637
tri 933 1615 955 1637 sw
tri 1140 1615 1162 1637 se
rect 1162 1615 1171 1637
rect 485 1603 792 1615
tri 792 1603 804 1615 sw
tri 889 1603 901 1615 ne
rect 901 1603 1171 1615
rect 1205 1603 1211 1637
tri 485 1589 499 1603 ne
rect 499 1600 804 1603
tri 804 1600 807 1603 sw
tri 901 1600 904 1603 ne
rect 904 1600 1211 1603
rect 499 1591 807 1600
tri 807 1591 816 1600 sw
tri 904 1591 913 1600 ne
rect 913 1591 1211 1600
rect 499 1589 816 1591
tri 816 1589 818 1591 sw
tri 913 1589 915 1591 ne
rect 915 1589 1209 1591
tri 1209 1589 1211 1591 nw
rect 1250 1695 1438 1733
tri 1438 1724 1447 1733 nw
tri 1624 1724 1633 1733 ne
rect 1250 1661 1327 1695
rect 1361 1661 1438 1695
rect 1250 1623 1438 1661
rect 1250 1589 1327 1623
rect 1361 1589 1438 1623
tri 499 1508 580 1589 ne
rect 580 1577 818 1589
tri 818 1577 830 1589 sw
tri 915 1577 927 1589 ne
rect 927 1577 1197 1589
tri 1197 1577 1209 1589 nw
rect 580 1569 830 1577
tri 830 1569 838 1577 sw
tri 927 1569 935 1577 ne
rect 935 1569 1189 1577
tri 1189 1569 1197 1577 nw
rect 580 1503 838 1569
tri 838 1503 904 1569 sw
rect 1250 1531 1438 1589
rect 1477 1709 1523 1721
rect 1477 1675 1483 1709
rect 1517 1675 1523 1709
rect 1477 1637 1523 1675
rect 1633 1717 1786 1733
tri 1786 1717 1818 1749 nw
tri 1835 1717 1867 1749 se
rect 1867 1717 1871 1749
rect 1633 1695 1756 1717
rect 1633 1661 1639 1695
rect 1673 1687 1756 1695
tri 1756 1687 1786 1717 nw
tri 1805 1687 1835 1717 se
rect 1835 1687 1871 1717
tri 1871 1687 1937 1753 nw
tri 1968 1687 2034 1753 se
rect 2034 1687 2691 1753
rect 1673 1661 1718 1687
rect 1633 1649 1718 1661
tri 1718 1649 1756 1687 nw
tri 1767 1649 1805 1687 se
rect 1805 1683 1867 1687
tri 1867 1683 1871 1687 nw
tri 1964 1683 1968 1687 se
rect 1968 1683 2691 1687
rect 1805 1651 1835 1683
tri 1835 1651 1867 1683 nw
tri 1932 1651 1964 1683 se
rect 1964 1661 2691 1683
rect 1964 1651 2186 1661
rect 1805 1649 1833 1651
tri 1833 1649 1835 1651 nw
tri 1930 1649 1932 1651 se
rect 1932 1649 2186 1651
tri 1758 1640 1767 1649 se
rect 1767 1640 1805 1649
rect 1477 1603 1483 1637
rect 1517 1621 1523 1637
tri 1523 1621 1542 1640 sw
tri 1739 1621 1758 1640 se
rect 1758 1621 1805 1640
tri 1805 1621 1833 1649 nw
tri 1902 1621 1930 1649 se
rect 1930 1621 2186 1649
rect 1517 1615 1542 1621
tri 1542 1615 1548 1621 sw
tri 1733 1615 1739 1621 se
rect 1739 1615 1799 1621
tri 1799 1615 1805 1621 nw
tri 1896 1615 1902 1621 se
rect 1902 1615 2186 1621
rect 1517 1603 1775 1615
rect 1477 1591 1775 1603
tri 1775 1591 1799 1615 nw
tri 1872 1591 1896 1615 se
rect 1896 1591 2186 1615
tri 1477 1577 1491 1591 ne
rect 1491 1577 1753 1591
tri 1491 1569 1499 1577 ne
rect 1499 1569 1753 1577
tri 1753 1569 1775 1591 nw
tri 1867 1586 1872 1591 se
rect 1872 1586 2186 1591
tri 2186 1586 2261 1661 nw
tri 2349 1636 2374 1661 ne
rect 2374 1636 2420 1661
tri 2420 1636 2445 1661 nw
tri 2608 1636 2633 1661 ne
tri 1850 1569 1867 1586 se
rect 1867 1569 2108 1586
tri 1812 1531 1850 1569 se
rect 1850 1531 2108 1569
tri 1784 1503 1812 1531 se
rect 1812 1503 2108 1531
tri 2108 1508 2186 1586 nw
rect 580 1286 2108 1503
rect 580 477 743 1286
tri 743 1236 793 1286 nw
tri 984 1261 1009 1286 ne
rect 1009 1261 1055 1286
tri 1055 1261 1080 1286 nw
tri 1296 1261 1321 1286 ne
rect 1321 1261 1367 1286
tri 1367 1261 1392 1286 nw
tri 1608 1261 1633 1286 ne
rect 1633 1261 1679 1286
tri 1679 1261 1704 1286 nw
tri 1895 1261 1920 1286 ne
rect 1920 1261 2108 1286
tri 1920 1236 1945 1261 ne
rect 1945 477 2108 1261
tri 2522 477 2530 485 se
rect 2530 477 2576 485
tri 2500 455 2522 477 se
rect 2522 455 2576 477
tri 80 423 112 455 se
rect 112 423 158 455
tri 158 423 190 455 sw
tri 392 423 424 455 se
rect 424 423 470 455
tri 470 423 502 455 sw
tri 821 423 853 455 se
rect 853 423 899 455
tri 899 423 931 455 sw
tri 1133 423 1165 455 se
rect 1165 423 1211 455
tri 1445 423 1477 455 se
rect 1477 423 1523 455
tri 1523 423 1555 455 sw
tri 1757 423 1789 455 se
rect 1789 423 1835 455
tri 1835 423 1867 455 sw
tri 2186 423 2218 455 se
rect 2218 423 2264 455
tri 2264 423 2296 455 sw
tri 2468 423 2500 455 se
rect 2500 423 2576 455
rect -3 309 1211 423
rect -3 281 383 309
tri 383 281 411 309 nw
tri 1261 281 1286 306 se
rect 1286 281 2576 423
rect -3 153 255 281
tri 255 153 383 281 nw
rect 423 275 2576 281
rect 603 167 2576 275
rect 2633 171 2691 1661
rect 423 153 603 159
tri 603 153 617 167 nw
rect -3 136 238 153
tri 238 136 255 153 nw
rect -3 130 232 136
tri 232 130 238 136 nw
tri 620 130 626 136 se
rect 626 130 756 136
rect -3 96 198 130
tri 198 96 232 130 nw
tri 586 96 620 130 se
rect 620 96 638 130
rect 672 96 710 130
rect 744 96 756 130
rect -3 90 192 96
tri 192 90 198 96 nw
tri 580 90 586 96 se
rect 586 90 756 96
rect 2361 130 2694 136
rect 2361 96 2373 130
rect 2407 96 2445 130
rect 2479 96 2694 130
rect 2361 90 2694 96
tri 567 77 580 90 se
rect 580 86 756 90
rect 580 77 747 86
tri 747 77 756 86 nw
rect 567 71 683 77
rect 619 19 631 71
rect 567 13 683 19
tri 683 13 747 77 nw
<< rmetal1 >>
rect 499 7749 557 7750
rect 499 7748 500 7749
rect 556 7748 557 7749
rect 1011 7749 1069 7750
rect 1011 7748 1012 7749
rect 1068 7748 1069 7749
rect 499 7711 500 7712
rect 556 7711 557 7712
rect 499 7710 557 7711
rect 1011 7711 1012 7712
rect 1068 7711 1069 7712
rect 1011 7710 1069 7711
rect 2035 7749 2093 7750
rect 2035 7748 2036 7749
rect 2092 7748 2093 7749
rect 2035 7711 2036 7712
rect 2092 7711 2093 7712
rect 2035 7710 2093 7711
rect 1243 2141 1289 2142
rect 1243 2140 1244 2141
rect 1288 2140 1289 2141
rect 1243 2103 1244 2104
rect 1288 2103 1289 2104
rect 1243 2102 1289 2103
rect 1555 2141 1601 2142
rect 1555 2140 1556 2141
rect 1600 2140 1601 2141
rect 1555 2103 1556 2104
rect 1600 2103 1601 2104
rect 1555 2102 1601 2103
rect 1243 1919 1289 1920
rect 1243 1918 1244 1919
rect 1288 1918 1289 1919
rect 1243 1881 1244 1882
rect 1288 1881 1289 1882
rect 1243 1880 1289 1881
rect 1555 1919 1601 1920
rect 1555 1918 1556 1919
rect 1600 1918 1601 1919
rect 1555 1881 1556 1882
rect 1600 1881 1601 1882
rect 1555 1880 1601 1881
<< via1 >>
rect 567 8568 619 8620
rect 567 8504 619 8556
rect 567 8440 619 8492
rect 43 7422 223 7538
rect 308 7422 488 7538
rect 567 7486 619 7538
rect 567 7422 619 7474
rect 107 7305 159 7357
rect 171 7305 223 7357
rect 1113 7009 1165 7061
rect 1113 6945 1165 6997
rect 1221 5817 1273 5869
rect 1221 5753 1273 5805
rect 1005 5568 1057 5620
rect 1221 5568 1273 5620
rect 1005 5504 1057 5556
rect 1221 5504 1273 5556
rect 1113 4625 1165 4677
rect 1113 4561 1165 4613
rect 1005 3752 1057 3804
rect 1221 3752 1273 3804
rect 1005 3688 1057 3740
rect 1221 3688 1273 3740
rect 1221 3433 1273 3485
rect 1221 3369 1273 3421
rect 567 2397 619 2449
rect 257 2246 309 2298
rect 257 2182 309 2234
rect 567 2333 619 2385
rect 2200 7422 2380 7538
rect 2465 7305 2517 7357
rect 2529 7305 2581 7357
rect 1523 7009 1575 7061
rect 1523 6945 1575 6997
rect 1415 5887 1467 5939
rect 1415 5823 1467 5875
rect 1415 5568 1467 5620
rect 1631 5568 1683 5620
rect 1415 5504 1467 5556
rect 1631 5504 1683 5556
rect 1523 4625 1575 4677
rect 1523 4561 1575 4613
rect 1415 3752 1467 3804
rect 1631 3752 1683 3804
rect 1415 3688 1467 3740
rect 1631 3688 1683 3740
rect 1415 3503 1467 3555
rect 1415 3439 1467 3491
rect 2069 2397 2121 2449
rect 1286 2282 1338 2334
rect 1350 2282 1402 2334
rect 2069 2333 2121 2385
rect 567 2007 619 2059
rect 567 1943 619 1995
rect 2069 2007 2121 2059
rect 2069 1943 2121 1995
rect 423 159 603 275
rect 567 19 619 71
rect 631 19 683 71
<< metal2 >>
rect 26 7538 229 8816
rect 26 7422 43 7538
rect 223 7422 229 7538
rect 26 7416 229 7422
rect 285 7538 511 8816
rect 285 7422 308 7538
rect 488 7422 511 7538
rect 0 7305 107 7357
rect 159 7305 171 7357
rect 223 7305 229 7357
rect 0 430 229 7305
rect 285 2378 511 7422
rect 567 8620 619 8816
rect 567 8556 619 8568
rect 567 8492 619 8504
rect 567 7538 619 8440
rect 675 8439 1057 8816
tri 675 8434 680 8439 ne
rect 680 8434 1057 8439
tri 680 8403 711 8434 ne
tri 680 7544 711 7575 se
rect 567 7474 619 7486
rect 567 2503 619 7422
tri 680 7385 711 7416 ne
rect 711 5620 1057 8434
rect 711 5568 1005 5620
rect 711 5556 1057 5568
rect 711 5504 1005 5556
rect 711 3804 1057 5504
rect 711 3752 1005 3804
rect 711 3740 1057 3752
rect 711 3688 1005 3740
tri 285 2333 330 2378 ne
rect 330 2333 511 2378
tri 330 2326 337 2333 ne
rect 257 2298 309 2304
rect 257 2234 309 2246
rect 257 689 309 2182
rect 337 852 511 2333
rect 567 2449 619 2455
rect 567 2385 619 2397
rect 567 2059 619 2333
rect 567 1995 619 2007
rect 567 925 619 1943
tri 699 925 711 937 se
rect 711 925 1057 3688
tri 675 901 699 925 se
rect 699 901 1057 925
tri 511 852 560 901 sw
tri 626 852 675 901 se
rect 675 852 1057 901
rect 337 705 1057 852
tri 337 693 349 705 ne
rect 349 693 1057 705
tri 309 689 313 693 sw
tri 349 689 353 693 ne
rect 353 689 1057 693
rect 257 671 313 689
tri 257 615 313 671 ne
tri 313 655 347 689 sw
tri 353 655 387 689 ne
rect 387 655 1057 689
rect 313 615 347 655
tri 347 615 387 655 sw
tri 387 615 427 655 ne
rect 427 615 1057 655
tri 313 541 387 615 ne
tri 387 581 421 615 sw
tri 427 581 461 615 ne
rect 461 581 1057 615
rect 387 541 421 581
tri 421 541 461 581 sw
tri 461 541 501 581 ne
rect 501 541 1057 581
tri 387 467 461 541 ne
tri 461 507 495 541 sw
tri 501 507 535 541 ne
rect 535 507 1057 541
rect 461 467 495 507
tri 495 467 535 507 sw
tri 535 467 575 507 ne
rect 575 467 1057 507
tri 461 430 498 467 ne
rect 498 433 535 467
tri 535 433 569 467 sw
tri 575 433 609 467 ne
rect 609 433 1057 467
rect 498 430 569 433
tri 569 430 572 433 sw
tri 609 430 612 433 ne
rect 612 430 1057 433
tri 498 393 535 430 ne
rect 535 393 572 430
tri 572 393 609 430 sw
tri 612 393 649 430 ne
rect 649 393 1057 430
tri 535 319 609 393 ne
tri 609 359 643 393 sw
tri 649 359 683 393 ne
rect 683 359 1057 393
rect 609 331 643 359
tri 643 331 671 359 sw
tri 683 331 711 359 ne
rect 609 319 671 331
tri 671 319 683 331 sw
tri 609 297 631 319 ne
rect 423 275 603 281
rect 423 153 603 159
rect 423 141 591 153
tri 591 141 603 153 nw
rect 423 117 567 141
tri 567 117 591 141 nw
tri 607 117 631 141 se
rect 631 117 683 319
rect 423 101 551 117
tri 551 101 567 117 nw
tri 591 101 607 117 se
rect 607 101 683 117
rect 711 101 1057 359
rect 1113 7061 1165 8816
rect 1113 6997 1165 7009
rect 1113 5983 1165 6945
rect 1221 6066 1467 8816
tri 1221 6039 1248 6066 ne
rect 1248 6039 1440 6066
tri 1440 6039 1467 6066 nw
rect 1523 7061 1575 8816
rect 1523 6997 1575 7009
tri 1165 5983 1192 6010 sw
rect 1113 5945 1429 5983
tri 1429 5945 1467 5983 sw
rect 1113 5939 1467 5945
rect 1113 5931 1415 5939
rect 1113 4677 1165 5931
tri 1165 5904 1192 5931 nw
tri 1388 5904 1415 5931 ne
rect 1415 5875 1467 5887
rect 1221 5869 1273 5875
rect 1415 5817 1467 5823
rect 1221 5805 1273 5817
tri 1273 5761 1300 5788 sw
tri 1496 5761 1523 5788 se
rect 1523 5761 1575 6945
rect 1273 5753 1575 5761
rect 1221 5747 1575 5753
tri 1221 5709 1259 5747 ne
rect 1259 5709 1575 5747
tri 1496 5682 1523 5709 ne
rect 1113 4613 1165 4625
rect 1113 3599 1165 4561
tri 1221 5626 1248 5653 se
rect 1248 5626 1440 5653
tri 1440 5626 1467 5653 sw
rect 1221 5620 1467 5626
rect 1273 5568 1415 5620
rect 1221 5556 1467 5568
rect 1273 5504 1415 5556
rect 1221 3804 1467 5504
rect 1273 3752 1415 3804
rect 1221 3740 1467 3752
rect 1273 3688 1415 3740
rect 1221 3682 1467 3688
tri 1221 3655 1248 3682 ne
rect 1248 3655 1440 3682
tri 1440 3655 1467 3682 nw
rect 1523 4677 1575 5709
rect 1523 4613 1575 4625
tri 1165 3599 1192 3626 sw
rect 1113 3561 1429 3599
tri 1429 3561 1467 3599 sw
rect 1113 3555 1467 3561
rect 1113 3547 1415 3555
rect 1113 101 1165 3547
tri 1165 3520 1192 3547 nw
tri 1388 3520 1415 3547 ne
rect 1415 3491 1467 3503
rect 1221 3485 1273 3491
rect 1415 3433 1467 3439
rect 1221 3421 1273 3433
tri 1273 3377 1300 3404 sw
tri 1496 3377 1523 3404 se
rect 1523 3377 1575 4561
rect 1273 3369 1575 3377
rect 1221 3363 1575 3369
tri 1221 3325 1259 3363 ne
rect 1259 3325 1575 3363
tri 1496 3298 1523 3325 ne
tri 1221 3242 1248 3269 se
rect 1248 3242 1440 3269
tri 1440 3242 1467 3269 sw
rect 1221 2334 1467 3242
rect 1221 2282 1286 2334
rect 1338 2282 1350 2334
rect 1402 2282 1467 2334
tri 1193 2089 1221 2117 se
rect 1221 2089 1467 2282
tri 1467 2089 1495 2117 sw
rect 1193 2087 1495 2089
rect 1193 101 1258 2087
tri 1258 2062 1283 2087 nw
tri 1405 2062 1430 2087 ne
rect 1286 101 1402 1531
rect 1430 101 1495 2087
rect 1523 101 1575 3325
rect 1631 5620 2013 8816
rect 1683 5568 2013 5620
rect 1631 5556 2013 5568
rect 1683 5504 2013 5556
rect 1631 3804 2013 5504
rect 1683 3752 2013 3804
rect 1631 3740 2013 3752
rect 1683 3688 2013 3740
rect 1631 101 2013 3688
rect 2069 2449 2121 8816
rect 2069 2385 2121 2397
rect 2069 2059 2121 2333
rect 2069 1995 2121 2007
rect 2069 101 2121 1943
rect 2177 7538 2403 7544
rect 2177 7422 2200 7538
rect 2380 7422 2403 7538
rect 2177 538 2403 7422
rect 2177 101 2310 538
tri 2310 445 2403 538 nw
rect 2459 7305 2465 7357
rect 2517 7305 2529 7357
rect 2581 7305 2688 7357
rect 2459 524 2688 7305
tri 2459 445 2538 524 ne
rect 2366 101 2482 167
rect 2538 101 2688 524
rect 423 89 539 101
tri 539 89 551 101 nw
tri 579 89 591 101 se
rect 591 89 683 101
tri 567 77 579 89 se
rect 579 77 683 89
rect 567 71 683 77
rect 619 19 631 71
rect 567 13 683 19
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_0
timestamp 1707688321
transform 0 -1 893 -1 0 1884
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_1
timestamp 1707688321
transform 0 1 1795 -1 0 1884
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_2
timestamp 1707688321
transform -1 0 2377 0 1 2288
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_3
timestamp 1707688321
transform 0 1 1405 1 0 1932
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_4
timestamp 1707688321
transform 0 1 1093 1 0 1932
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_5
timestamp 1707688321
transform 0 1 1249 1 0 1932
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_6
timestamp 1707688321
transform 0 1 1561 1 0 1932
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_7
timestamp 1707688321
transform 0 1 1483 1 0 1603
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_8
timestamp 1707688321
transform 0 -1 1205 1 0 1603
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_9
timestamp 1707688321
transform 1 0 2373 0 -1 130
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_10
timestamp 1707688321
transform 1 0 638 0 -1 130
box 0 0 1 1
use L1M1_CDNS_5246887918590  L1M1_CDNS_5246887918590_0
timestamp 1707688321
transform 0 1 1639 1 0 1661
box 0 0 1 1
use L1M1_CDNS_5246887918590  L1M1_CDNS_5246887918590_1
timestamp 1707688321
transform 0 -1 1049 1 0 1661
box 0 0 1 1
use L1M1_CDNS_52468879185191  L1M1_CDNS_52468879185191_0
timestamp 1707688321
transform 0 1 2360 -1 0 7047
box -12 -6 838 40
use L1M1_CDNS_52468879185195  L1M1_CDNS_52468879185195_0
timestamp 1707688321
transform -1 0 2009 0 1 2288
box -12 -6 550 40
use L1M1_CDNS_52468879185195  L1M1_CDNS_52468879185195_1
timestamp 1707688321
transform 1 0 679 0 1 2288
box -12 -6 550 40
use L1M1_CDNS_52468879185196  L1M1_CDNS_52468879185196_0
timestamp 1707688321
transform 0 -1 1361 1 0 1589
box 0 0 1 1
use L1M1_CDNS_52468879185307  L1M1_CDNS_52468879185307_0
timestamp 1707688321
transform 0 1 2536 1 0 201
box -12 -6 1414 40
use L1M1_CDNS_52468879185307  L1M1_CDNS_52468879185307_1
timestamp 1707688321
transform 0 -1 152 1 0 201
box -12 -6 1414 40
use L1M1_CDNS_52468879185308  L1M1_CDNS_52468879185308_0
timestamp 1707688321
transform 1 0 96 0 1 2099
box 0 0 1 1
use L1M1_CDNS_52468879185335  L1M1_CDNS_52468879185335_0
timestamp 1707688321
transform 1 0 61 0 1 7506
box -12 -6 1126 40
use L1M1_CDNS_52468879185381  L1M1_CDNS_52468879185381_0
timestamp 1707688321
transform 0 1 1171 -1 0 1242
box -12 -6 910 40
use L1M1_CDNS_52468879185381  L1M1_CDNS_52468879185381_1
timestamp 1707688321
transform 0 1 859 -1 0 1242
box -12 -6 910 40
use L1M1_CDNS_52468879185381  L1M1_CDNS_52468879185381_2
timestamp 1707688321
transform -1 0 2550 0 1 2099
box -12 -6 910 40
use L1M1_CDNS_52468879185381  L1M1_CDNS_52468879185381_3
timestamp 1707688321
transform -1 0 2339 0 1 7506
box -12 -6 910 40
use L1M1_CDNS_52468879185448  L1M1_CDNS_52468879185448_0
timestamp 1707688321
transform 0 1 2068 1 0 489
box -12 -6 1270 40
use L1M1_CDNS_52468879185448  L1M1_CDNS_52468879185448_1
timestamp 1707688321
transform 0 -1 620 1 0 489
box -12 -6 1270 40
use L1M1_CDNS_52468879185955  L1M1_CDNS_52468879185955_0
timestamp 1707688321
transform -1 0 1275 0 1 7106
box -12 -6 982 40
use L1M1_CDNS_52468879185955  L1M1_CDNS_52468879185955_1
timestamp 1707688321
transform 0 1 703 1 0 489
box -12 -6 982 40
use L1M1_CDNS_52468879185955  L1M1_CDNS_52468879185955_2
timestamp 1707688321
transform 0 1 1015 1 0 489
box -12 -6 982 40
use L1M1_CDNS_52468879185955  L1M1_CDNS_52468879185955_3
timestamp 1707688321
transform 0 -1 1985 1 0 489
box -12 -6 982 40
use L1M1_CDNS_52468879185955  L1M1_CDNS_52468879185955_4
timestamp 1707688321
transform 0 -1 1673 1 0 489
box -12 -6 982 40
use L1M1_CDNS_52468879185955  L1M1_CDNS_52468879185955_5
timestamp 1707688321
transform 0 -1 1361 1 0 489
box -12 -6 982 40
use L1M1_CDNS_52468879185955  L1M1_CDNS_52468879185955_6
timestamp 1707688321
transform 1 0 1413 0 1 7106
box -12 -6 982 40
use L1M1_CDNS_524688791851011  L1M1_CDNS_524688791851011_0
timestamp 1707688321
transform 0 -1 464 -1 0 1530
box -12 -6 1198 40
use L1M1_CDNS_524688791851011  L1M1_CDNS_524688791851011_1
timestamp 1707688321
transform -1 0 2599 0 1 7317
box -12 -6 1198 40
use L1M1_CDNS_524688791851011  L1M1_CDNS_524688791851011_2
timestamp 1707688321
transform 1 0 89 0 1 7317
box -12 -6 1198 40
use L1M1_CDNS_524688791851012  L1M1_CDNS_524688791851012_0
timestamp 1707688321
transform 0 1 2380 1 0 489
box -12 -6 1486 40
use L1M1_CDNS_524688791851012  L1M1_CDNS_524688791851012_1
timestamp 1707688321
transform 0 -1 308 1 0 489
box -12 -6 1486 40
use L1M1_CDNS_524688791851014  L1M1_CDNS_524688791851014_0
timestamp 1707688321
transform -1 0 289 0 -1 8393
box -12 -6 46 760
use L1M1_CDNS_524688791851014  L1M1_CDNS_524688791851014_1
timestamp 1707688321
transform -1 0 2337 0 -1 8393
box -12 -6 46 760
use L1M1_CDNS_524688791851015  L1M1_CDNS_524688791851015_0
timestamp 1707688321
transform -1 0 2490 0 -1 7113
box -12 -6 46 904
use L1M1_CDNS_524688791851016  L1M1_CDNS_524688791851016_0
timestamp 1707688321
transform -1 0 545 0 -1 8372
box -12 -6 46 616
use L1M1_CDNS_524688791851016  L1M1_CDNS_524688791851016_1
timestamp 1707688321
transform -1 0 1057 0 -1 8372
box -12 -6 46 616
use L1M1_CDNS_524688791851016  L1M1_CDNS_524688791851016_2
timestamp 1707688321
transform -1 0 1569 0 -1 8372
box -12 -6 46 616
use L1M1_CDNS_524688791851016  L1M1_CDNS_524688791851016_3
timestamp 1707688321
transform -1 0 2081 0 -1 8372
box -12 -6 46 616
use L1M1_CDNS_524688791851016  L1M1_CDNS_524688791851016_4
timestamp 1707688321
transform 0 1 1421 1 0 7021
box -12 -6 46 616
use L1M1_CDNS_524688791851016  L1M1_CDNS_524688791851016_5
timestamp 1707688321
transform 0 1 1421 1 0 4637
box -12 -6 46 616
use L1M1_CDNS_524688791851016  L1M1_CDNS_524688791851016_6
timestamp 1707688321
transform 0 1 1421 1 0 3445
box -12 -6 46 616
use L1M1_CDNS_524688791851016  L1M1_CDNS_524688791851016_7
timestamp 1707688321
transform 0 1 1421 1 0 5829
box -12 -6 46 616
use L1M1_CDNS_524688791851016  L1M1_CDNS_524688791851016_8
timestamp 1707688321
transform 0 -1 1267 1 0 7021
box -12 -6 46 616
use L1M1_CDNS_524688791851016  L1M1_CDNS_524688791851016_9
timestamp 1707688321
transform 0 -1 1267 1 0 3445
box -12 -6 46 616
use L1M1_CDNS_524688791851016  L1M1_CDNS_524688791851016_10
timestamp 1707688321
transform 0 -1 1267 1 0 5829
box -12 -6 46 616
use L1M1_CDNS_524688791851016  L1M1_CDNS_524688791851016_11
timestamp 1707688321
transform 0 -1 1267 1 0 4637
box -12 -6 46 616
use L1M1_CDNS_524688791851018  L1M1_CDNS_524688791851018_0
timestamp 1707688321
transform -1 0 801 0 1 7762
box -12 -6 46 832
use L1M1_CDNS_524688791851018  L1M1_CDNS_524688791851018_1
timestamp 1707688321
transform -1 0 1313 0 1 7762
box -12 -6 46 832
use L1M1_CDNS_524688791851018  L1M1_CDNS_524688791851018_2
timestamp 1707688321
transform -1 0 1825 0 1 7762
box -12 -6 46 832
use L1M1_CDNS_524688791851037  L1M1_CDNS_524688791851037_0
timestamp 1707688321
transform 0 1 2360 1 0 2393
box -12 -6 3646 40
use L1M1_CDNS_524688791851038  L1M1_CDNS_524688791851038_0
timestamp 1707688321
transform -1 0 2490 0 1 2321
box -12 -6 46 3712
use L1M1_CDNS_524688791851039  L1M1_CDNS_524688791851039_0
timestamp 1707688321
transform 0 -1 328 1 0 2393
box -12 -6 4654 40
use L1M1_CDNS_524688791851040  L1M1_CDNS_524688791851040_0
timestamp 1707688321
transform 0 -1 1829 1 0 201
box -12 -6 1054 40
use L1M1_CDNS_524688791851040  L1M1_CDNS_524688791851040_1
timestamp 1707688321
transform 0 -1 1517 1 0 201
box -12 -6 1054 40
use L1M1_CDNS_524688791851041  L1M1_CDNS_524688791851041_0
timestamp 1707688321
transform 1 0 2645 0 -1 7267
box -12 -6 46 7096
use L1M1_CDNS_524688791851042  L1M1_CDNS_524688791851042_0
timestamp 1707688321
transform 0 1 2224 1 0 200
box -12 -6 1342 40
use L1M1_CDNS_524688791851043  L1M1_CDNS_524688791851043_0
timestamp 1707688321
transform -1 0 232 0 -1 7107
box -12 -6 46 4720
use L1M1_CDNS_524688791851044  L1M1_CDNS_524688791851044_0
timestamp 1707688321
transform -1 0 43 0 -1 7260
box -12 -6 46 5008
use L1M1_CDNS_524688791851045  L1M1_CDNS_524688791851045_0
timestamp 1707688321
transform -1 0 43 0 1 515
box -12 -6 46 1624
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_0
timestamp 1707688321
transform 0 1 1415 -1 0 5945
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_1
timestamp 1707688321
transform 0 1 1415 -1 0 3561
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_2
timestamp 1707688321
transform -1 0 229 0 1 7305
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_3
timestamp 1707688321
transform 0 1 567 1 0 2327
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_4
timestamp 1707688321
transform 0 1 567 1 0 1937
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_5
timestamp 1707688321
transform 0 1 2069 1 0 2327
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_6
timestamp 1707688321
transform 0 1 2069 1 0 1937
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_7
timestamp 1707688321
transform 0 1 1523 1 0 6939
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_8
timestamp 1707688321
transform 0 1 1523 1 0 4555
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_9
timestamp 1707688321
transform 0 1 257 1 0 2176
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_10
timestamp 1707688321
transform 0 1 1221 1 0 5498
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_11
timestamp 1707688321
transform 0 1 1005 1 0 5498
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_12
timestamp 1707688321
transform 0 1 1221 1 0 3682
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_13
timestamp 1707688321
transform 0 1 1005 1 0 3682
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_14
timestamp 1707688321
transform 0 -1 1165 1 0 4555
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_15
timestamp 1707688321
transform 0 -1 1165 1 0 6939
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_16
timestamp 1707688321
transform 0 -1 1273 1 0 5747
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_17
timestamp 1707688321
transform 0 -1 1273 1 0 3363
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_18
timestamp 1707688321
transform 0 -1 619 1 0 7416
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_19
timestamp 1707688321
transform 0 -1 1683 1 0 5498
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_20
timestamp 1707688321
transform 0 -1 1467 1 0 5498
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_21
timestamp 1707688321
transform 0 -1 1683 1 0 3682
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_22
timestamp 1707688321
transform 0 -1 1467 1 0 3682
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_23
timestamp 1707688321
transform 1 0 1280 0 -1 2334
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_24
timestamp 1707688321
transform 1 0 2459 0 1 7305
box 0 0 1 1
use M1M2_CDNS_52468879185197  M1M2_CDNS_52468879185197_0
timestamp 1707688321
transform 0 1 2366 -1 0 423
box 0 0 256 116
use M1M2_CDNS_52468879185197  M1M2_CDNS_52468879185197_1
timestamp 1707688321
transform 0 1 1286 -1 0 423
box 0 0 256 116
use M1M2_CDNS_52468879185200  M1M2_CDNS_52468879185200_0
timestamp 1707688321
transform 0 1 2200 1 0 7416
box 0 0 1 1
use M1M2_CDNS_52468879185200  M1M2_CDNS_52468879185200_1
timestamp 1707688321
transform 0 1 423 1 0 153
box 0 0 1 1
use M1M2_CDNS_52468879185200  M1M2_CDNS_52468879185200_2
timestamp 1707688321
transform 0 -1 488 1 0 7416
box 0 0 1 1
use M1M2_CDNS_52468879185200  M1M2_CDNS_52468879185200_3
timestamp 1707688321
transform 0 -1 223 1 0 7416
box 0 0 1 1
use M1M2_CDNS_52468879185201  M1M2_CDNS_52468879185201_0
timestamp 1707688321
transform 0 1 1286 -1 0 1851
box 0 0 320 116
use M1M2_CDNS_52468879185203  M1M2_CDNS_52468879185203_0
timestamp 1707688321
transform 0 -1 619 -1 0 8626
box 0 0 1 1
use M1M2_CDNS_52468879185208  M1M2_CDNS_52468879185208_0
timestamp 1707688321
transform 0 -1 1466 -1 0 8626
box 0 0 192 244
use M1M2_CDNS_52468879185369  M1M2_CDNS_52468879185369_0
timestamp 1707688321
transform 0 1 567 1 0 13
box 0 0 1 1
use M1M2_CDNS_52468879185975  M1M2_CDNS_52468879185975_0
timestamp 1707688321
transform 0 -1 488 -1 0 8626
box 0 0 192 180
use M1M2_CDNS_524688791851023  M1M2_CDNS_524688791851023_0
timestamp 1707688321
transform 0 1 2351 -1 0 7050
box 0 0 832 52
use M1M2_CDNS_524688791851030  M1M2_CDNS_524688791851030_0
timestamp 1707688321
transform 0 1 2351 1 0 2378
box 0 0 3648 52
use M1M2_CDNS_524688791851031  M1M2_CDNS_524688791851031_0
timestamp 1707688321
transform 0 -1 1052 1 0 7416
box 0 0 128 372
use M1M2_CDNS_524688791851031  M1M2_CDNS_524688791851031_1
timestamp 1707688321
transform 0 -1 2008 1 0 7416
box 0 0 128 372
use M1M2_CDNS_524688791851032  M1M2_CDNS_524688791851032_0
timestamp 1707688321
transform 0 -1 2008 -1 0 8626
box 0 0 192 372
use M1M2_CDNS_524688791851032  M1M2_CDNS_524688791851032_1
timestamp 1707688321
transform 0 -1 1052 -1 0 8626
box 0 0 192 372
use M1M2_CDNS_524688791851033  M1M2_CDNS_524688791851033_0
timestamp 1707688321
transform 0 1 285 1 0 2378
box 0 0 4672 52
use M1M2_CDNS_524688791851034  M1M2_CDNS_524688791851034_0
timestamp 1707688321
transform 0 -1 2688 -1 0 7306
box 0 0 7104 52
use M1M2_CDNS_524688791851035  M1M2_CDNS_524688791851035_0
timestamp 1707688321
transform 0 1 0 -1 0 7306
box 0 0 5056 52
use M1M2_CDNS_524688791851036  M1M2_CDNS_524688791851036_0
timestamp 1707688321
transform 0 1 0 1 0 509
box 0 0 1600 52
use nfet_CDNS_524688791851024  nfet_CDNS_524688791851024_0
timestamp 1707688321
transform -1 0 756 0 1 7640
box -79 -52 535 1052
use nfet_CDNS_524688791851024  nfet_CDNS_524688791851024_1
timestamp 1707688321
transform -1 0 1268 0 1 7640
box -79 -52 535 1052
use nfet_CDNS_524688791851024  nfet_CDNS_524688791851024_2
timestamp 1707688321
transform -1 0 1780 0 1 7640
box -79 -52 535 1052
use nfet_CDNS_524688791851024  nfet_CDNS_524688791851024_3
timestamp 1707688321
transform -1 0 2292 0 1 7640
box -79 -52 535 1052
use nfet_CDNS_524688791851046  nfet_CDNS_524688791851046_0
timestamp 1707688321
transform -1 0 2172 0 1 3589
box -79 -52 879 1052
use nfet_CDNS_524688791851046  nfet_CDNS_524688791851046_1
timestamp 1707688321
transform -1 0 2172 0 1 5973
box -79 -52 879 1052
use nfet_CDNS_524688791851046  nfet_CDNS_524688791851046_2
timestamp 1707688321
transform -1 0 1316 0 1 3589
box -79 -52 879 1052
use nfet_CDNS_524688791851046  nfet_CDNS_524688791851046_3
timestamp 1707688321
transform -1 0 1316 0 1 5973
box -79 -52 879 1052
use nfet_CDNS_524688791851046  nfet_CDNS_524688791851046_4
timestamp 1707688321
transform 1 0 1372 0 1 2397
box -79 -52 879 1052
use nfet_CDNS_524688791851046  nfet_CDNS_524688791851046_5
timestamp 1707688321
transform 1 0 516 0 1 2397
box -79 -52 879 1052
use nfet_CDNS_524688791851046  nfet_CDNS_524688791851046_6
timestamp 1707688321
transform 1 0 516 0 1 4781
box -79 -52 879 1052
use nfet_CDNS_524688791851046  nfet_CDNS_524688791851046_7
timestamp 1707688321
transform 1 0 1372 0 1 4781
box -79 -52 879 1052
use nfet_CDNS_524688791851047  nfet_CDNS_524688791851047_0
timestamp 1707688321
transform -1 0 2328 0 1 5973
box -79 -52 182 1052
use nfet_CDNS_524688791851047  nfet_CDNS_524688791851047_1
timestamp 1707688321
transform -1 0 2328 0 1 4781
box -79 -52 182 1052
use nfet_CDNS_524688791851047  nfet_CDNS_524688791851047_2
timestamp 1707688321
transform -1 0 2328 0 1 3589
box -79 -52 182 1052
use nfet_CDNS_524688791851047  nfet_CDNS_524688791851047_3
timestamp 1707688321
transform -1 0 2328 0 1 2397
box -79 -52 182 1052
use nfet_CDNS_524688791851047  nfet_CDNS_524688791851047_4
timestamp 1707688321
transform 1 0 360 0 1 4781
box -79 -52 182 1052
use nfet_CDNS_524688791851047  nfet_CDNS_524688791851047_5
timestamp 1707688321
transform 1 0 360 0 1 3589
box -79 -52 182 1052
use nfet_CDNS_524688791851047  nfet_CDNS_524688791851047_6
timestamp 1707688321
transform 1 0 360 0 1 2397
box -79 -52 182 1052
use nfet_CDNS_524688791851047  nfet_CDNS_524688791851047_7
timestamp 1707688321
transform 1 0 360 0 1 5973
box -79 -52 182 1052
use pfet_CDNS_524688791851048  pfet_CDNS_524688791851048_0
timestamp 1707688321
transform -1 0 1004 0 1 1598
box -119 -66 219 366
use pfet_CDNS_524688791851048  pfet_CDNS_524688791851048_1
timestamp 1707688321
transform -1 0 1472 0 1 1598
box -119 -66 219 366
use pfet_CDNS_524688791851048  pfet_CDNS_524688791851048_2
timestamp 1707688321
transform -1 0 1160 0 1 1598
box -119 -66 219 366
use pfet_CDNS_524688791851048  pfet_CDNS_524688791851048_3
timestamp 1707688321
transform -1 0 1628 0 1 1598
box -119 -66 219 366
use pfet_CDNS_524688791851048  pfet_CDNS_524688791851048_4
timestamp 1707688321
transform -1 0 1316 0 1 1598
box -119 -66 219 366
use pfet_CDNS_524688791851048  pfet_CDNS_524688791851048_5
timestamp 1707688321
transform 1 0 1684 0 1 1598
box -119 -66 219 366
use pfet_CDNS_524688791851049  pfet_CDNS_524688791851049_0
timestamp 1707688321
transform -1 0 575 0 1 595
box -119 -66 531 1466
use pfet_CDNS_524688791851049  pfet_CDNS_524688791851049_1
timestamp 1707688321
transform 1 0 2113 0 1 595
box -119 -66 531 1466
use pfet_CDNS_524688791851050  pfet_CDNS_524688791851050_0
timestamp 1707688321
transform -1 0 1940 0 1 438
box -119 -66 1311 1066
use pfet_CDNS_524688791851051  pfet_CDNS_524688791851051_0
timestamp 1707688321
transform -1 0 1940 0 -1 378
box -119 -66 1311 266
use pfet_CDNS_524688791851052  pfet_CDNS_524688791851052_0
timestamp 1707688321
transform -1 0 575 0 1 178
box -119 -66 531 366
use pfet_CDNS_524688791851052  pfet_CDNS_524688791851052_1
timestamp 1707688321
transform -1 0 2525 0 1 178
box -119 -66 531 366
use PYL1_CDNS_5246887918526  PYL1_CDNS_5246887918526_0
timestamp 1707688321
transform 0 1 1701 -1 0 2064
box 0 0 1 1
use PYL1_CDNS_5246887918526  PYL1_CDNS_5246887918526_1
timestamp 1707688321
transform 0 1 921 -1 0 2064
box 0 0 1 1
use PYL1_CDNS_5246887918526  PYL1_CDNS_5246887918526_2
timestamp 1707688321
transform 0 1 1389 -1 0 2064
box 0 0 1 1
use PYL1_CDNS_5246887918526  PYL1_CDNS_5246887918526_3
timestamp 1707688321
transform 0 1 1545 -1 0 2064
box 0 0 1 1
use PYL1_CDNS_5246887918526  PYL1_CDNS_5246887918526_4
timestamp 1707688321
transform 0 1 1077 -1 0 2064
box 0 0 1 1
use PYL1_CDNS_5246887918526  PYL1_CDNS_5246887918526_5
timestamp 1707688321
transform 0 1 1233 -1 0 2064
box 0 0 1 1
use PYL1_CDNS_5246887918526  PYL1_CDNS_5246887918526_6
timestamp 1707688321
transform -1 0 460 0 -1 3495
box 0 0 1 1
use PYL1_CDNS_5246887918526  PYL1_CDNS_5246887918526_7
timestamp 1707688321
transform -1 0 460 0 -1 7071
box 0 0 1 1
use PYL1_CDNS_5246887918526  PYL1_CDNS_5246887918526_8
timestamp 1707688321
transform -1 0 460 0 -1 4687
box 0 0 1 1
use PYL1_CDNS_5246887918526  PYL1_CDNS_5246887918526_9
timestamp 1707688321
transform -1 0 2362 0 -1 3495
box 0 0 1 1
use PYL1_CDNS_5246887918526  PYL1_CDNS_5246887918526_10
timestamp 1707688321
transform -1 0 460 0 -1 5879
box 0 0 1 1
use PYL1_CDNS_5246887918526  PYL1_CDNS_5246887918526_11
timestamp 1707688321
transform -1 0 2362 0 -1 4687
box 0 0 1 1
use PYL1_CDNS_5246887918526  PYL1_CDNS_5246887918526_12
timestamp 1707688321
transform -1 0 2362 0 -1 5879
box 0 0 1 1
use PYL1_CDNS_5246887918526  PYL1_CDNS_5246887918526_13
timestamp 1707688321
transform -1 0 2362 0 -1 7071
box 0 0 1 1
use PYL1_CDNS_5246887918562  PYL1_CDNS_5246887918562_0
timestamp 1707688321
transform 0 1 1869 1 0 8672
box 0 0 1 1
use PYL1_CDNS_5246887918562  PYL1_CDNS_5246887918562_1
timestamp 1707688321
transform 0 1 1613 1 0 8672
box 0 0 1 1
use PYL1_CDNS_5246887918562  PYL1_CDNS_5246887918562_2
timestamp 1707688321
transform 0 1 1357 1 0 8672
box 0 0 1 1
use PYL1_CDNS_5246887918562  PYL1_CDNS_5246887918562_3
timestamp 1707688321
transform 0 1 1101 1 0 8672
box 0 0 1 1
use PYL1_CDNS_5246887918562  PYL1_CDNS_5246887918562_4
timestamp 1707688321
transform 0 1 845 1 0 8672
box 0 0 1 1
use PYL1_CDNS_5246887918562  PYL1_CDNS_5246887918562_5
timestamp 1707688321
transform 0 1 589 1 0 8672
box 0 0 1 1
use PYL1_CDNS_5246887918562  PYL1_CDNS_5246887918562_6
timestamp 1707688321
transform 0 1 333 1 0 8672
box 0 0 1 1
use PYL1_CDNS_5246887918562  PYL1_CDNS_5246887918562_7
timestamp 1707688321
transform 0 1 2125 1 0 8672
box 0 0 1 1
use PYL1_CDNS_524688791851028  PYL1_CDNS_524688791851028_0
timestamp 1707688321
transform -1 0 1289 0 -1 7071
box 0 0 746 66
use PYL1_CDNS_524688791851028  PYL1_CDNS_524688791851028_1
timestamp 1707688321
transform -1 0 2145 0 -1 7071
box 0 0 746 66
use PYL1_CDNS_524688791851028  PYL1_CDNS_524688791851028_2
timestamp 1707688321
transform -1 0 1289 0 -1 5879
box 0 0 746 66
use PYL1_CDNS_524688791851028  PYL1_CDNS_524688791851028_3
timestamp 1707688321
transform -1 0 2145 0 -1 5879
box 0 0 746 66
use PYL1_CDNS_524688791851028  PYL1_CDNS_524688791851028_4
timestamp 1707688321
transform -1 0 1289 0 -1 4687
box 0 0 746 66
use PYL1_CDNS_524688791851028  PYL1_CDNS_524688791851028_5
timestamp 1707688321
transform -1 0 2145 0 -1 4687
box 0 0 746 66
use PYL1_CDNS_524688791851028  PYL1_CDNS_524688791851028_6
timestamp 1707688321
transform -1 0 1289 0 -1 3495
box 0 0 746 66
use PYL1_CDNS_524688791851028  PYL1_CDNS_524688791851028_7
timestamp 1707688321
transform -1 0 2145 0 -1 3495
box 0 0 746 66
use PYL1_CDNS_524688791851029  PYL1_CDNS_524688791851029_0
timestamp 1707688321
transform 0 1 1405 1 0 80
box 0 0 66 1086
use PYL1_CDNS_524688791851029  PYL1_CDNS_524688791851029_1
timestamp 1707688321
transform 0 -1 1283 1 0 80
box 0 0 66 1086
use sky130_fd_io__tk_em1o_CDNS_52468879185340  sky130_fd_io__tk_em1o_CDNS_52468879185340_0
timestamp 1707688321
transform 0 1 1555 -1 0 2194
box 0 0 1 1
use sky130_fd_io__tk_em1o_CDNS_52468879185340  sky130_fd_io__tk_em1o_CDNS_52468879185340_1
timestamp 1707688321
transform 0 1 1243 -1 0 2194
box 0 0 1 1
use sky130_fd_io__tk_em1o_CDNS_52468879185985  sky130_fd_io__tk_em1o_CDNS_52468879185985_0
timestamp 1707688321
transform 0 1 499 -1 0 7802
box 0 0 1 1
use sky130_fd_io__tk_em1o_CDNS_52468879185985  sky130_fd_io__tk_em1o_CDNS_52468879185985_1
timestamp 1707688321
transform 0 1 1011 -1 0 7802
box 0 0 1 1
use sky130_fd_io__tk_em1o_CDNS_52468879185985  sky130_fd_io__tk_em1o_CDNS_52468879185985_2
timestamp 1707688321
transform 0 1 2035 -1 0 7802
box 0 0 1 1
use sky130_fd_io__tk_em1s_CDNS_52468879185341  sky130_fd_io__tk_em1s_CDNS_52468879185341_0
timestamp 1707688321
transform 0 1 1243 -1 0 1972
box 0 0 1 1
use sky130_fd_io__tk_em1s_CDNS_52468879185341  sky130_fd_io__tk_em1s_CDNS_52468879185341_1
timestamp 1707688321
transform 0 1 1555 -1 0 1972
box 0 0 1 1
<< labels >>
flabel comment s 494 7177 494 7177 0 FreeSans 1000 0 0 0 condiode
flabel metal1 s 70 2176 111 2222 3 FreeSans 200 0 0 0 ibuf_sel_h_n
port 4 nsew
flabel metal1 s 2670 90 2694 136 3 FreeSans 200 180 0 0 en_outop_h_n
port 2 nsew
flabel metal1 s -3 90 26 423 3 FreeSans 200 180 0 0 vcc_virt_i
port 3 nsew
flabel metal1 s 291 8682 345 8728 3 FreeSans 200 0 0 0 ngate
port 5 nsew
flabel metal2 s 0 430 229 455 3 FreeSans 200 0 0 0 vcc
port 6 nsew
flabel metal2 s 2538 101 2688 122 3 FreeSans 200 90 0 0 vcc
port 6 nsew
flabel metal2 s 2177 101 2310 122 3 FreeSans 200 90 0 0 vgnd
port 7 nsew
flabel metal2 s 1430 101 1495 122 3 FreeSans 200 90 0 0 vgnd
port 7 nsew
flabel metal2 s 1193 101 1258 122 3 FreeSans 200 90 0 0 vgnd
port 7 nsew
flabel metal2 s 1286 101 1402 122 3 FreeSans 200 90 0 0 vcc_virt_o
port 8 nsew
flabel metal2 s 2366 101 2482 122 3 FreeSans 200 90 0 0 vcc_virt_o
port 8 nsew
flabel metal2 s 567 13 683 34 3 FreeSans 200 90 0 0 ibuf_sel_h_n
port 4 nsew
flabel metal2 s 1523 101 1575 122 3 FreeSans 200 90 0 0 inn
port 9 nsew
flabel metal2 s 1113 101 1165 122 3 FreeSans 200 90 0 0 inp
port 10 nsew
flabel metal2 s 711 101 1057 122 3 FreeSans 200 90 0 0 vgnd
port 7 nsew
flabel metal2 s 2069 101 2121 122 3 FreeSans 200 90 0 0 out
port 11 nsew
flabel metal2 s 423 101 539 122 3 FreeSans 200 90 0 0 vcc_virt_o
port 8 nsew
flabel metal2 s 1631 101 2013 122 3 FreeSans 200 90 0 0 vgnd
port 7 nsew
<< properties >>
string GDS_END 80360890
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 80295898
string path 0.650 11.400 0.650 182.900 
<< end >>
