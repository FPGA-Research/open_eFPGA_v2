magic
tech sky130B
magscale 1 2
timestamp 1707688321
<< nwell >>
rect -91 1479 403 2319
rect 1573 2154 1879 2312
rect -91 61 340 739
rect 651 52 817 784
<< pwell >>
rect 463 1355 549 2253
rect 1427 1154 1513 2253
rect 2059 1208 2145 1460
rect 960 97 1046 749
<< psubdiff >>
rect 1453 2203 1487 2227
rect 1453 2135 1487 2169
rect 1453 2066 1487 2101
rect 1453 1997 1487 2032
rect 1453 1928 1487 1963
rect 1453 1859 1487 1894
rect 1453 1790 1487 1825
rect 1453 1721 1487 1756
rect 1453 1652 1487 1687
rect 1453 1583 1487 1618
rect 1453 1514 1487 1549
rect 1453 1445 1487 1480
rect 1453 1376 1487 1411
rect 1453 1307 1487 1342
rect 2085 1410 2119 1434
rect 1453 1238 1487 1273
rect 2085 1292 2119 1376
rect 2085 1234 2119 1258
rect 1453 1180 1487 1204
<< nsubdiff >>
rect 1609 2242 1633 2276
rect 1667 2242 1709 2276
rect 1743 2242 1785 2276
rect 1819 2242 1843 2276
<< mvpsubdiff >>
rect 489 2203 523 2227
rect 489 2134 523 2169
rect 489 2065 523 2100
rect 489 1996 523 2031
rect 489 1927 523 1962
rect 489 1858 523 1893
rect 489 1789 523 1824
rect 489 1719 523 1755
rect 489 1649 523 1685
rect 489 1579 523 1615
rect 489 1509 523 1545
rect 489 1439 523 1475
rect 489 1381 523 1405
rect 986 699 1020 723
rect 986 625 1020 665
rect 986 551 1020 591
rect 986 477 1020 517
rect 986 403 1020 443
rect 986 329 1020 369
rect 986 255 1020 295
rect 986 181 1020 221
rect 986 123 1020 147
<< mvnsubdiff >>
rect 0 2219 43 2253
rect 77 2219 121 2253
rect 155 2219 200 2253
rect 234 2219 279 2253
rect 313 2219 337 2253
rect 717 694 751 718
rect 717 620 751 660
rect 717 546 751 586
rect -17 469 153 493
rect -17 343 153 367
rect 717 472 751 512
rect 717 398 751 438
rect 717 324 751 364
rect 717 250 751 290
rect 717 176 751 216
rect 717 118 751 142
<< psubdiffcont >>
rect 1453 2169 1487 2203
rect 1453 2101 1487 2135
rect 1453 2032 1487 2066
rect 1453 1963 1487 1997
rect 1453 1894 1487 1928
rect 1453 1825 1487 1859
rect 1453 1756 1487 1790
rect 1453 1687 1487 1721
rect 1453 1618 1487 1652
rect 1453 1549 1487 1583
rect 1453 1480 1487 1514
rect 1453 1411 1487 1445
rect 1453 1342 1487 1376
rect 2085 1376 2119 1410
rect 1453 1273 1487 1307
rect 1453 1204 1487 1238
rect 2085 1258 2119 1292
<< nsubdiffcont >>
rect 1633 2242 1667 2276
rect 1709 2242 1743 2276
rect 1785 2242 1819 2276
<< mvpsubdiffcont >>
rect 489 2169 523 2203
rect 489 2100 523 2134
rect 489 2031 523 2065
rect 489 1962 523 1996
rect 489 1893 523 1927
rect 489 1824 523 1858
rect 489 1755 523 1789
rect 489 1685 523 1719
rect 489 1615 523 1649
rect 489 1545 523 1579
rect 489 1475 523 1509
rect 489 1405 523 1439
rect 986 665 1020 699
rect 986 591 1020 625
rect 986 517 1020 551
rect 986 443 1020 477
rect 986 369 1020 403
rect 986 295 1020 329
rect 986 221 1020 255
rect 986 147 1020 181
<< mvnsubdiffcont >>
rect 43 2219 77 2253
rect 121 2219 155 2253
rect 200 2219 234 2253
rect 279 2219 313 2253
rect 717 660 751 694
rect 717 586 751 620
rect 717 512 751 546
rect -17 367 153 469
rect 717 438 751 472
rect 717 364 751 398
rect 717 290 751 324
rect 717 216 751 250
rect 717 142 751 176
<< poly >>
rect 650 2253 1302 2319
rect 1754 2204 2009 2224
rect 1754 2188 1891 2204
rect 1875 2170 1891 2188
rect 1925 2170 1959 2204
rect 1993 2170 2009 2204
rect 1875 2154 2009 2170
rect 650 1632 830 2001
rect 909 1952 1043 2013
rect 909 1918 957 1952
rect 991 1918 1043 1952
rect 909 1884 1043 1918
rect 909 1850 957 1884
rect 991 1850 1043 1884
rect 909 1816 1043 1850
rect 909 1782 957 1816
rect 991 1782 1043 1816
rect 909 1672 1043 1782
rect 1122 1632 1302 2001
rect 28 1513 128 1519
rect 184 1513 284 1519
rect 28 1497 284 1513
rect 28 1463 44 1497
rect 78 1463 112 1497
rect 146 1463 180 1497
rect 214 1463 284 1497
rect 28 1447 284 1463
rect 1908 1593 1974 1609
rect 1908 1559 1924 1593
rect 1958 1559 1974 1593
rect 650 1383 1302 1443
rect 1662 1339 1698 1536
rect 1754 1336 1790 1536
rect 1908 1525 1974 1559
rect 1908 1496 1924 1525
rect 1846 1491 1924 1496
rect 1958 1491 1974 1525
rect 1846 1460 1974 1491
rect 86 999 206 1188
rect 28 983 207 999
rect 28 949 89 983
rect 123 949 157 983
rect 191 949 207 983
rect 262 976 382 1188
rect 1662 1166 1698 1208
rect 1662 1150 2050 1166
rect 1662 1116 1932 1150
rect 1966 1116 2000 1150
rect 2034 1116 2050 1150
rect 1662 1100 2050 1116
rect 682 1089 952 1093
rect 1023 1089 1293 1093
rect 670 1077 958 1089
rect 670 1043 698 1077
rect 732 1043 766 1077
rect 800 1043 834 1077
rect 868 1043 902 1077
rect 936 1043 958 1077
rect 670 1023 958 1043
rect 1014 1077 1302 1089
rect 1014 1043 1039 1077
rect 1073 1043 1107 1077
rect 1141 1043 1175 1077
rect 1209 1043 1243 1077
rect 1277 1043 1302 1077
rect 1014 1023 1302 1043
rect 262 972 414 976
rect 28 933 207 949
rect 264 956 414 972
rect 28 735 128 933
rect 264 922 280 956
rect 314 922 348 956
rect 382 922 414 956
rect 264 906 414 922
rect 294 744 414 906
rect 1545 854 1679 857
rect 1801 854 1935 857
rect 1486 841 1686 854
rect 456 800 590 816
rect 456 766 472 800
rect 506 766 540 800
rect 574 766 590 800
rect 1486 807 1561 841
rect 1595 807 1629 841
rect 1663 807 1686 841
rect 1486 791 1686 807
rect 1742 841 1942 854
rect 1742 807 1817 841
rect 1851 807 1885 841
rect 1919 807 1942 841
rect 1742 791 1942 807
rect 456 750 590 766
rect 470 744 590 750
rect 28 0 414 92
rect 470 66 590 92
rect 456 50 590 66
rect 456 16 472 50
rect 506 16 540 50
rect 574 16 590 50
rect 456 0 590 16
rect 1147 66 1267 97
rect 1433 66 1553 97
rect 1609 66 1729 97
rect 1147 50 1553 66
rect 1147 16 1163 50
rect 1197 16 1231 50
rect 1265 16 1299 50
rect 1333 16 1367 50
rect 1401 16 1435 50
rect 1469 16 1503 50
rect 1537 16 1553 50
rect 1147 0 1553 16
rect 1595 50 1729 66
rect 1595 16 1611 50
rect 1645 16 1679 50
rect 1713 16 1729 50
rect 1595 0 1729 16
rect 1785 66 1905 97
rect 1785 50 1919 66
rect 1785 16 1801 50
rect 1835 16 1869 50
rect 1903 16 1919 50
rect 1785 0 1919 16
<< polycont >>
rect 1891 2170 1925 2204
rect 1959 2170 1993 2204
rect 957 1918 991 1952
rect 957 1850 991 1884
rect 957 1782 991 1816
rect 44 1463 78 1497
rect 112 1463 146 1497
rect 180 1463 214 1497
rect 1924 1559 1958 1593
rect 1924 1491 1958 1525
rect 89 949 123 983
rect 157 949 191 983
rect 1932 1116 1966 1150
rect 2000 1116 2034 1150
rect 698 1043 732 1077
rect 766 1043 800 1077
rect 834 1043 868 1077
rect 902 1043 936 1077
rect 1039 1043 1073 1077
rect 1107 1043 1141 1077
rect 1175 1043 1209 1077
rect 1243 1043 1277 1077
rect 280 922 314 956
rect 348 922 382 956
rect 472 766 506 800
rect 540 766 574 800
rect 1561 807 1595 841
rect 1629 807 1663 841
rect 1817 807 1851 841
rect 1885 807 1919 841
rect 472 16 506 50
rect 540 16 574 50
rect 1163 16 1197 50
rect 1231 16 1265 50
rect 1299 16 1333 50
rect 1367 16 1401 50
rect 1435 16 1469 50
rect 1503 16 1537 50
rect 1611 16 1645 50
rect 1679 16 1713 50
rect 1801 16 1835 50
rect 1869 16 1903 50
<< locali >>
rect 841 2259 1419 2293
rect 0 2226 43 2253
rect 77 2226 121 2253
rect 155 2226 200 2253
rect 234 2226 279 2253
rect 17 2219 43 2226
rect 89 2219 121 2226
rect 17 2192 55 2219
rect 89 2192 127 2219
rect 161 2192 199 2226
rect 234 2219 271 2226
rect 313 2219 337 2253
rect 233 2192 271 2219
rect 489 2203 523 2227
rect 841 2225 875 2259
rect 1313 2225 1419 2259
rect 1549 2242 1633 2276
rect 1667 2242 1709 2276
rect 1743 2242 1785 2276
rect 1819 2242 2119 2276
rect 489 2134 523 2169
rect -17 2002 17 2040
rect -17 1930 17 1968
rect 295 2002 329 2040
rect 295 1930 329 1968
rect 489 2065 523 2100
rect 489 1996 523 2031
rect 605 1965 639 2059
rect 841 1965 875 2105
rect 957 2002 991 2040
rect 1111 2023 1251 2225
rect 1341 2023 1419 2225
rect 489 1927 523 1962
rect 957 1952 991 1968
rect 489 1858 523 1893
rect 941 1896 957 1952
rect 991 1896 1007 1952
rect 941 1884 1007 1896
rect 941 1850 957 1884
rect 991 1850 1007 1884
rect 489 1789 523 1824
rect 639 1816 677 1850
rect 941 1816 1007 1850
rect 1145 1850 1251 2023
rect 1179 1816 1217 1850
rect 941 1782 957 1816
rect 991 1782 1007 1816
rect 489 1719 523 1755
rect 1077 1735 1111 1763
rect 489 1649 523 1685
rect 605 1701 1111 1735
rect 605 1656 639 1701
rect 139 1589 173 1607
rect 139 1555 142 1589
rect 176 1555 214 1589
rect 489 1579 523 1615
rect 904 1605 942 1639
rect 1077 1638 1111 1701
rect 1313 1655 1347 1763
rect 1275 1605 1313 1639
rect 139 1549 173 1555
rect 489 1509 523 1545
rect 158 1497 196 1509
rect 28 1463 44 1497
rect 78 1463 112 1497
rect 158 1475 180 1497
rect 146 1463 180 1475
rect 214 1463 230 1475
rect 489 1439 523 1475
rect 217 1357 251 1395
rect 217 1285 251 1323
rect 217 1245 251 1251
rect 489 1357 523 1395
rect 605 1419 639 1471
rect 1381 1419 1419 2023
rect 605 1385 917 1419
rect 489 1285 523 1323
rect 489 1205 523 1251
rect 625 1279 659 1317
rect 711 1308 745 1385
rect 797 1279 831 1317
rect 883 1308 917 1385
rect 1055 1385 1419 1419
rect 1453 2203 1487 2227
rect 1453 2135 1487 2169
rect 1549 2226 1583 2242
rect 2085 2226 2119 2242
rect 1549 2154 1583 2192
rect 1875 2170 1891 2204
rect 1925 2170 1959 2204
rect 1993 2170 2026 2204
rect 1453 2066 1487 2101
rect 1453 1997 1487 2032
rect 1453 1928 1487 1963
rect 1453 1859 1487 1894
rect 1617 1850 1651 2118
rect 1453 1790 1487 1825
rect 1579 1816 1617 1850
rect 1453 1721 1487 1756
rect 1453 1652 1487 1687
rect 1453 1583 1487 1618
rect 1453 1514 1487 1549
rect 1453 1445 1487 1480
rect 1617 1432 1651 1816
rect 1777 1682 1835 2166
rect 1992 1850 2026 2170
rect 2085 2154 2119 2192
rect 1954 1816 1992 1850
rect 1777 1624 1885 1682
rect 1709 1583 1743 1624
rect 1719 1549 1757 1583
rect 1825 1497 1885 1624
rect 1777 1466 1885 1497
rect 1924 1593 1958 1609
rect 1924 1525 1958 1547
rect 969 1279 1003 1317
rect 1055 1308 1089 1385
rect 1141 1279 1175 1317
rect 1227 1308 1261 1385
rect 1453 1376 1487 1395
rect 1313 1279 1347 1317
rect 1453 1307 1487 1323
rect 1453 1238 1487 1251
rect 495 1171 533 1205
rect 1453 1202 1487 1204
rect 217 1089 251 1132
rect 75 1050 113 1084
rect 393 1053 450 1087
rect 121 983 159 1009
rect 73 975 87 983
rect 73 949 89 975
rect 123 949 157 983
rect 193 975 207 983
rect 191 949 207 975
rect 258 956 382 972
rect 258 922 280 956
rect 314 922 348 956
rect 258 906 382 922
rect 258 855 323 906
rect 416 872 450 1053
rect 484 935 546 1171
rect 1415 1168 1453 1202
rect 1521 1256 1651 1432
rect 1704 1429 1738 1432
rect 1704 1395 1709 1429
rect 1704 1357 1743 1395
rect 1704 1323 1709 1357
rect 1704 1285 1743 1323
rect 1521 1230 1627 1256
rect 1704 1251 1709 1285
rect 736 1077 774 1083
rect 808 1077 846 1083
rect 880 1077 918 1083
rect 1521 1078 1555 1230
rect 682 1043 698 1077
rect 736 1049 766 1077
rect 808 1049 834 1077
rect 880 1049 902 1077
rect 732 1043 766 1049
rect 800 1043 834 1049
rect 868 1043 902 1049
rect 936 1043 952 1049
rect 1023 1077 1555 1078
rect 1023 1043 1039 1077
rect 1073 1043 1107 1077
rect 1141 1043 1175 1077
rect 1209 1043 1243 1077
rect 1277 1044 1555 1077
rect 1277 1043 1293 1044
rect 1704 1010 1738 1251
rect 1777 1063 1859 1466
rect 1893 1357 1927 1395
rect 1893 1285 1927 1323
rect 1992 1230 2026 1816
rect 2085 1410 2119 1434
rect 2085 1292 2119 1376
rect 2085 1199 2119 1258
rect 1932 1150 2039 1166
rect 1966 1116 2000 1150
rect 2034 1116 2039 1150
rect 1932 1085 2039 1116
rect 1811 1029 1849 1063
rect 1932 1051 1933 1085
rect 1967 1051 2005 1085
rect 2085 1127 2119 1165
rect 614 975 652 1009
rect 518 901 556 935
rect 139 821 172 855
rect 206 821 244 855
rect 278 821 323 855
rect 357 838 450 872
rect 139 722 173 821
rect 357 722 391 838
rect 624 836 686 975
rect 1591 955 1629 989
rect 1441 855 1475 881
rect 493 802 686 836
rect 1064 821 1102 855
rect 1439 821 1477 855
rect 1564 841 1663 955
rect 1704 865 1747 1010
rect 1815 955 1853 989
rect 1887 955 1987 989
rect 493 800 590 802
rect 456 766 472 800
rect 506 766 540 800
rect 574 766 590 800
rect -17 493 105 722
rect 257 697 391 722
rect 257 663 283 697
rect 317 663 355 697
rect 389 663 391 697
rect 257 628 391 663
rect -17 469 153 493
rect -17 343 153 367
rect -17 280 105 343
rect 17 246 105 280
rect -17 208 105 246
rect 17 174 105 208
rect -17 136 105 174
rect 17 102 105 136
rect 139 68 215 272
rect 425 208 459 246
rect 425 136 459 174
rect 493 68 567 766
rect 624 696 658 734
rect 1102 727 1136 821
rect 1545 807 1561 841
rect 1595 807 1629 841
rect 1663 807 1679 841
rect 1278 775 1330 781
rect 1278 741 1296 775
rect 1278 727 1330 741
rect 624 180 658 662
rect 717 694 751 718
rect 717 620 751 660
rect 717 546 751 586
rect 717 472 751 512
rect 717 398 751 438
rect 717 324 751 364
rect 717 280 751 290
rect 717 208 751 216
rect 717 136 751 142
rect 986 699 1020 723
rect 986 625 1020 665
rect 986 551 1020 591
rect 986 477 1020 517
rect 986 438 1020 443
rect 986 403 1020 404
rect 986 366 1020 369
rect 986 329 1020 332
rect 986 255 1020 295
rect 986 181 1020 221
rect 1296 703 1330 727
rect 1296 185 1330 669
rect 1370 775 1422 781
rect 1404 741 1422 775
rect 1370 727 1422 741
rect 1564 727 1598 807
rect 1713 771 1747 865
rect 2085 929 2119 1093
rect 2085 857 2119 895
rect 1849 841 1887 855
rect 1801 821 1815 841
rect 1801 807 1817 821
rect 1851 807 1885 841
rect 1921 821 1950 841
rect 1919 807 1950 821
rect 1370 703 1404 727
rect 1370 185 1404 669
rect 1713 699 1747 737
rect 1916 727 1950 807
rect 1713 185 1747 665
rect 986 123 1020 147
rect 1102 151 1136 185
rect 1916 151 1950 185
rect 1102 117 1950 151
rect 139 50 567 68
rect 139 16 472 50
rect 506 16 540 50
rect 574 16 590 50
rect 1147 16 1163 50
rect 1197 16 1231 50
rect 1265 16 1299 50
rect 1333 16 1367 50
rect 1401 16 1435 50
rect 1469 16 1503 50
rect 1537 16 1553 50
rect 1595 16 1611 50
rect 1645 16 1679 50
rect 1713 16 1729 50
rect 1785 16 1801 50
rect 1835 16 1869 50
rect 1903 16 1919 50
<< viali >>
rect -17 2192 17 2226
rect 55 2219 77 2226
rect 77 2219 89 2226
rect 127 2219 155 2226
rect 155 2219 161 2226
rect 55 2192 89 2219
rect 127 2192 161 2219
rect 199 2219 200 2226
rect 200 2219 233 2226
rect 271 2219 279 2226
rect 279 2219 305 2226
rect 199 2192 233 2219
rect 271 2192 305 2219
rect -17 2040 17 2074
rect -17 1968 17 2002
rect -17 1896 17 1930
rect 295 2040 329 2074
rect 295 1968 329 2002
rect 295 1896 329 1930
rect 957 2040 991 2074
rect 957 1968 991 2002
rect 957 1918 991 1930
rect 957 1896 991 1918
rect 605 1816 639 1850
rect 677 1816 711 1850
rect 1145 1816 1179 1850
rect 1217 1816 1251 1850
rect 142 1555 176 1589
rect 214 1555 248 1589
rect 870 1605 904 1639
rect 942 1605 976 1639
rect 1241 1605 1275 1639
rect 1313 1605 1347 1639
rect 124 1497 158 1509
rect 196 1497 230 1509
rect 124 1475 146 1497
rect 146 1475 158 1497
rect 196 1475 214 1497
rect 214 1475 230 1497
rect 217 1395 251 1429
rect 217 1323 251 1357
rect 217 1251 251 1285
rect 489 1405 523 1429
rect 489 1395 523 1405
rect 489 1323 523 1357
rect 489 1251 523 1285
rect 625 1317 659 1351
rect 797 1317 831 1351
rect 625 1245 659 1279
rect 1549 2192 1583 2226
rect 1549 2120 1583 2154
rect 1545 1816 1579 1850
rect 1617 1816 1651 1850
rect 2085 2192 2119 2226
rect 2085 2120 2119 2154
rect 1920 1816 1954 1850
rect 1992 1816 2026 1850
rect 1685 1549 1719 1583
rect 1757 1549 1791 1583
rect 1924 1559 1958 1581
rect 1924 1547 1958 1559
rect 1924 1491 1958 1509
rect 1924 1475 1958 1491
rect 1453 1411 1487 1429
rect 1453 1395 1487 1411
rect 969 1317 1003 1351
rect 797 1245 831 1279
rect 1141 1317 1175 1351
rect 969 1245 1003 1279
rect 1313 1317 1347 1351
rect 1141 1245 1175 1279
rect 1313 1245 1347 1279
rect 1453 1342 1487 1357
rect 1453 1323 1487 1342
rect 1453 1273 1487 1285
rect 1453 1251 1487 1273
rect 461 1171 495 1205
rect 533 1171 567 1205
rect 41 1050 75 1084
rect 113 1050 147 1084
rect 87 983 121 1009
rect 159 983 193 1009
rect 87 975 89 983
rect 89 975 121 983
rect 159 975 191 983
rect 191 975 193 983
rect 1381 1168 1415 1202
rect 1453 1168 1487 1202
rect 1709 1395 1743 1429
rect 1709 1323 1743 1357
rect 1709 1251 1743 1285
rect 702 1077 736 1083
rect 774 1077 808 1083
rect 846 1077 880 1083
rect 918 1077 952 1083
rect 702 1049 732 1077
rect 732 1049 736 1077
rect 774 1049 800 1077
rect 800 1049 808 1077
rect 846 1049 868 1077
rect 868 1049 880 1077
rect 918 1049 936 1077
rect 936 1049 952 1077
rect 1893 1395 1927 1429
rect 1893 1323 1927 1357
rect 1893 1251 1927 1285
rect 1777 1029 1811 1063
rect 1849 1029 1883 1063
rect 1933 1051 1967 1085
rect 2005 1051 2039 1085
rect 2085 1165 2119 1199
rect 2085 1093 2119 1127
rect 580 975 614 1009
rect 652 975 686 1009
rect 484 901 518 935
rect 556 901 590 935
rect 172 821 206 855
rect 244 821 278 855
rect 1557 955 1591 989
rect 1629 955 1663 989
rect 1030 821 1064 855
rect 1102 821 1136 855
rect 1405 821 1439 855
rect 1477 821 1511 855
rect 1781 955 1815 989
rect 1853 955 1887 989
rect 283 663 317 697
rect 355 663 389 697
rect -17 246 17 280
rect -17 174 17 208
rect -17 102 17 136
rect 425 246 459 280
rect 425 174 459 208
rect 425 102 459 136
rect 624 734 658 768
rect 1296 741 1330 775
rect 624 662 658 696
rect 717 250 751 280
rect 717 246 751 250
rect 717 176 751 208
rect 717 174 751 176
rect 717 102 751 136
rect 986 404 1020 438
rect 986 332 1020 366
rect 1296 669 1330 703
rect 1370 741 1404 775
rect 2085 895 2119 929
rect 1815 841 1849 855
rect 1887 841 1921 855
rect 1815 821 1817 841
rect 1817 821 1849 841
rect 1887 821 1919 841
rect 1919 821 1921 841
rect 2085 823 2119 857
rect 1713 737 1747 771
rect 1370 669 1404 703
rect 1713 665 1747 699
<< metal1 >>
rect -31 2226 2131 2232
rect -31 2192 -17 2226
rect 17 2192 55 2226
rect 89 2192 127 2226
rect 161 2192 199 2226
rect 233 2192 271 2226
rect 305 2192 1549 2226
rect 1583 2192 2085 2226
rect 2119 2192 2131 2226
rect -31 2154 2131 2192
rect -31 2120 1549 2154
rect 1583 2120 2085 2154
rect 2119 2120 2131 2154
rect -31 2114 2131 2120
rect -39 2074 1917 2086
rect -39 2040 -17 2074
rect 17 2040 295 2074
rect 329 2040 957 2074
rect 991 2040 1917 2074
rect -39 2002 1917 2040
rect -39 1968 -17 2002
rect 17 1968 295 2002
rect 329 1968 957 2002
rect 991 1968 1917 2002
rect -39 1930 1917 1968
rect -39 1896 -17 1930
rect 17 1896 295 1930
rect 329 1896 957 1930
rect 991 1896 1917 1930
rect -39 1884 1917 1896
rect 593 1850 1290 1856
rect 593 1816 605 1850
rect 639 1816 677 1850
rect 711 1816 1145 1850
rect 1179 1816 1217 1850
rect 1251 1816 1290 1850
rect 593 1804 1290 1816
rect 1342 1804 1354 1856
rect 1406 1804 1412 1856
rect 1533 1850 2038 1856
rect 1533 1816 1545 1850
rect 1579 1816 1617 1850
rect 1651 1816 1920 1850
rect 1954 1816 1992 1850
rect 2026 1816 2038 1850
rect 1533 1810 2038 1816
tri 858 1645 864 1651 se
rect 864 1645 1370 1651
rect 858 1639 1370 1645
rect 858 1605 870 1639
rect 904 1605 942 1639
rect 976 1605 1241 1639
rect 1275 1605 1313 1639
rect 1347 1605 1370 1639
rect 858 1599 1370 1605
rect 1422 1599 1434 1651
rect 1486 1599 1492 1651
rect 130 1589 260 1595
tri 260 1589 266 1595 sw
rect 130 1555 142 1589
rect 176 1555 214 1589
rect 248 1583 266 1589
tri 266 1583 272 1589 sw
tri 1667 1583 1673 1589 se
rect 1673 1583 1803 1589
rect 248 1577 272 1583
tri 272 1577 278 1583 sw
tri 1661 1577 1667 1583 se
rect 1667 1577 1685 1583
rect 248 1571 725 1577
tri 725 1571 731 1577 sw
tri 1655 1571 1661 1577 se
rect 1661 1571 1685 1577
rect 248 1555 1685 1571
rect 130 1549 1685 1555
rect 1719 1549 1757 1583
rect 1791 1549 1803 1583
tri 695 1547 697 1549 ne
rect 697 1547 1803 1549
tri 697 1543 701 1547 ne
rect 701 1543 1803 1547
rect 1912 1581 1970 1587
rect 1912 1547 1924 1581
rect 1958 1547 1970 1581
tri 1887 1515 1912 1540 se
rect 1912 1515 1970 1547
rect 112 1509 1970 1515
rect 112 1475 124 1509
rect 158 1475 196 1509
rect 230 1475 1924 1509
rect 1958 1475 1970 1509
rect 112 1469 1970 1475
rect -25 1429 2102 1441
rect -25 1395 217 1429
rect 251 1395 489 1429
rect 523 1395 1453 1429
rect 1487 1395 1704 1429
rect 1756 1395 1893 1429
rect 1927 1395 2102 1429
rect -25 1377 1704 1395
rect 1756 1377 2102 1395
rect -25 1365 2102 1377
rect -25 1357 1704 1365
rect 1756 1357 2102 1365
rect -25 1323 217 1357
rect 251 1323 489 1357
rect 523 1351 1453 1357
rect 523 1323 625 1351
rect -25 1317 625 1323
rect 659 1317 797 1351
rect 831 1317 969 1351
rect 1003 1317 1141 1351
rect 1175 1317 1313 1351
rect 1347 1323 1453 1351
rect 1487 1323 1704 1357
rect 1756 1323 1893 1357
rect 1927 1323 2102 1357
rect 1347 1317 1704 1323
rect -25 1313 1704 1317
rect 1756 1313 2102 1323
rect -25 1301 2102 1313
rect -25 1285 1704 1301
rect 1756 1285 2102 1301
rect -25 1251 217 1285
rect 251 1251 489 1285
rect 523 1279 1453 1285
rect 523 1251 625 1279
rect -25 1245 625 1251
rect 659 1245 797 1279
rect 831 1245 969 1279
rect 1003 1245 1141 1279
rect 1175 1245 1313 1279
rect 1347 1251 1453 1279
rect 1487 1251 1704 1285
rect 1756 1251 1893 1285
rect 1927 1251 2102 1285
rect 1347 1249 1704 1251
rect 1756 1249 2102 1251
rect 1347 1245 2102 1249
rect -25 1239 2102 1245
rect 0 1159 456 1211
rect 508 1159 520 1211
rect 572 1202 2150 1211
rect 572 1168 1381 1202
rect 1415 1168 1453 1202
rect 1487 1199 2150 1202
rect 1487 1168 2085 1199
rect 572 1165 2085 1168
rect 2119 1165 2150 1199
rect 572 1159 2150 1165
tri 2054 1134 2079 1159 ne
rect 2079 1127 2125 1159
tri 2125 1134 2150 1159 nw
rect 29 1084 536 1095
rect 29 1050 41 1084
rect 75 1050 113 1084
rect 147 1050 536 1084
rect 29 1043 536 1050
rect 588 1043 600 1095
rect 652 1043 658 1095
rect 690 1085 965 1089
tri 965 1085 969 1089 sw
rect 1927 1085 2045 1097
rect 690 1083 969 1085
rect 690 1049 702 1083
rect 736 1049 774 1083
rect 808 1049 846 1083
rect 880 1049 918 1083
rect 952 1069 969 1083
tri 969 1069 985 1085 sw
rect 952 1063 985 1069
tri 985 1063 991 1069 sw
tri 1759 1063 1765 1069 se
rect 1765 1063 1895 1069
rect 952 1051 991 1063
tri 991 1051 1003 1063 sw
tri 1747 1051 1759 1063 se
rect 1759 1051 1777 1063
rect 952 1049 1777 1051
rect 690 1043 1777 1049
tri 891 1029 905 1043 ne
rect 905 1029 1777 1043
rect 1811 1029 1849 1063
rect 1883 1029 1895 1063
rect 1927 1051 1933 1085
rect 1967 1051 2005 1085
rect 2039 1051 2045 1085
rect 2079 1093 2085 1127
rect 2119 1093 2125 1127
rect 2079 1081 2125 1093
rect 1927 1039 2045 1051
tri 905 1023 911 1029 ne
rect 911 1023 1895 1029
rect 75 1009 737 1015
rect 75 975 87 1009
rect 121 975 159 1009
rect 193 975 580 1009
rect 614 975 652 1009
rect 686 995 737 1009
tri 737 995 757 1015 sw
rect 686 989 1899 995
rect 686 975 1557 989
rect 75 969 1557 975
tri 717 955 731 969 ne
rect 731 955 1557 969
rect 1591 955 1629 989
rect 1663 955 1781 989
rect 1815 955 1853 989
rect 1887 955 1899 989
tri 731 949 737 955 ne
rect 737 949 1899 955
rect 0 889 456 941
rect 508 935 520 941
rect 572 935 602 941
rect 518 901 520 935
rect 590 929 602 935
tri 602 929 614 941 sw
tri 1919 929 1931 941 se
rect 1931 929 2150 941
rect 590 921 614 929
tri 614 921 622 929 sw
tri 1911 921 1919 929 se
rect 1919 921 2085 929
rect 590 901 2085 921
rect 508 889 520 901
rect 572 895 2085 901
rect 2119 895 2150 929
rect 572 889 2150 895
tri 2054 864 2079 889 ne
rect 160 855 1933 861
rect 160 821 172 855
rect 206 821 244 855
rect 278 821 1030 855
rect 1064 821 1102 855
rect 1136 821 1405 855
rect 1439 821 1477 855
rect 1511 821 1815 855
rect 1849 821 1887 855
rect 1921 821 1933 855
rect 160 815 1933 821
rect 2079 857 2125 889
tri 2125 864 2150 889 nw
rect 2079 823 2085 857
rect 2119 823 2125 857
rect 2079 811 2125 823
rect 271 697 401 703
rect 271 663 283 697
rect 317 663 355 697
rect 389 663 401 697
rect 271 657 401 663
rect 530 671 536 787
rect 652 768 670 787
rect 658 734 670 768
rect 652 696 670 734
rect 530 662 624 671
rect 658 662 670 696
rect 530 656 670 662
rect 1284 781 1336 787
rect 1284 717 1336 729
rect 1284 657 1336 665
rect 1364 781 1416 787
rect 1364 717 1416 729
rect 1364 657 1416 665
rect 1701 781 1759 787
rect 1701 729 1704 781
rect 1756 729 1759 781
rect 1701 717 1759 729
rect 1701 665 1704 717
rect 1756 665 1759 717
rect 1701 659 1759 665
rect 0 442 2113 450
rect 0 390 450 442
rect 502 438 2113 442
rect 502 404 986 438
rect 1020 404 2113 438
rect 502 390 2113 404
rect 0 378 2113 390
rect 0 326 450 378
rect 502 366 2113 378
rect 502 332 986 366
rect 1020 332 2113 366
rect 502 326 2113 332
rect 0 320 2113 326
rect -23 280 2113 292
rect -23 246 -17 280
rect 17 246 425 280
rect 459 246 717 280
rect 751 246 2113 280
rect -23 208 2113 246
rect -23 174 -17 208
rect 17 174 425 208
rect 459 174 717 208
rect 751 174 2113 208
rect -23 136 2113 174
rect -23 102 -17 136
rect 17 102 425 136
rect 459 102 717 136
rect 751 102 2113 136
rect -23 90 2113 102
<< via1 >>
rect 1290 1804 1342 1856
rect 1354 1804 1406 1856
rect 1370 1599 1422 1651
rect 1434 1599 1486 1651
rect 1704 1395 1709 1429
rect 1709 1395 1743 1429
rect 1743 1395 1756 1429
rect 1704 1377 1756 1395
rect 1704 1357 1756 1365
rect 1704 1323 1709 1357
rect 1709 1323 1743 1357
rect 1743 1323 1756 1357
rect 1704 1313 1756 1323
rect 1704 1285 1756 1301
rect 1704 1251 1709 1285
rect 1709 1251 1743 1285
rect 1743 1251 1756 1285
rect 1704 1249 1756 1251
rect 456 1205 508 1211
rect 456 1171 461 1205
rect 461 1171 495 1205
rect 495 1171 508 1205
rect 456 1159 508 1171
rect 520 1205 572 1211
rect 520 1171 533 1205
rect 533 1171 567 1205
rect 567 1171 572 1205
rect 520 1159 572 1171
rect 536 1043 588 1095
rect 600 1043 652 1095
rect 456 935 508 941
rect 520 935 572 941
rect 456 901 484 935
rect 484 901 508 935
rect 520 901 556 935
rect 556 901 572 935
rect 456 889 508 901
rect 520 889 572 901
rect 536 768 652 787
rect 536 734 624 768
rect 624 734 652 768
rect 536 696 652 734
rect 536 671 624 696
rect 624 671 652 696
rect 1284 775 1336 781
rect 1284 741 1296 775
rect 1296 741 1330 775
rect 1330 741 1336 775
rect 1284 729 1336 741
rect 1284 703 1336 717
rect 1284 669 1296 703
rect 1296 669 1330 703
rect 1330 669 1336 703
rect 1284 665 1336 669
rect 1364 775 1416 781
rect 1364 741 1370 775
rect 1370 741 1404 775
rect 1404 741 1416 775
rect 1364 729 1416 741
rect 1364 703 1416 717
rect 1364 669 1370 703
rect 1370 669 1404 703
rect 1404 669 1416 703
rect 1364 665 1416 669
rect 1704 771 1756 781
rect 1704 737 1713 771
rect 1713 737 1747 771
rect 1747 737 1756 771
rect 1704 729 1756 737
rect 1704 699 1756 717
rect 1704 665 1713 699
rect 1713 665 1747 699
rect 1747 665 1756 699
rect 450 390 502 442
rect 450 326 502 378
<< metal2 >>
rect 1284 1804 1290 1856
rect 1342 1804 1354 1856
rect 1406 1804 1412 1856
rect 450 1159 456 1211
rect 508 1159 520 1211
rect 572 1159 578 1211
rect 450 941 502 1159
tri 502 1134 527 1159 nw
rect 530 1043 536 1095
rect 588 1043 600 1095
rect 652 1043 658 1095
tri 581 1018 606 1043 ne
tri 502 941 527 966 sw
rect 450 889 456 941
rect 508 889 520 941
rect 572 889 578 941
rect 450 442 502 889
tri 502 864 527 889 nw
tri 581 787 606 812 se
rect 606 787 658 1043
rect 530 671 536 787
rect 652 671 658 787
rect 1284 781 1336 1804
tri 1336 1779 1361 1804 nw
rect 1284 717 1336 729
rect 1284 659 1336 665
rect 1364 1599 1370 1651
rect 1422 1599 1434 1651
rect 1486 1599 1492 1651
rect 1364 781 1416 1599
tri 1416 1574 1441 1599 nw
rect 1364 717 1416 729
rect 1364 659 1416 665
rect 1704 1429 1756 1435
rect 1704 1365 1756 1377
rect 1704 1301 1756 1313
rect 1704 781 1756 1249
rect 1704 717 1756 729
rect 1704 659 1756 665
rect 450 378 502 390
rect 450 320 502 326
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_0
timestamp 1707688321
transform -1 0 1175 0 1 1245
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_1
timestamp 1707688321
transform -1 0 1003 0 1 1245
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_2
timestamp 1707688321
transform -1 0 831 0 1 1245
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_3
timestamp 1707688321
transform -1 0 659 0 1 1245
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_4
timestamp 1707688321
transform -1 0 1347 0 1 1245
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_5
timestamp 1707688321
transform 0 1 1933 1 0 1051
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_6
timestamp 1707688321
transform 1 0 1549 0 -1 2226
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_7
timestamp 1707688321
transform 1 0 624 0 -1 768
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_8
timestamp 1707688321
transform 1 0 1713 0 -1 771
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_9
timestamp 1707688321
transform 1 0 2085 0 -1 2226
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_10
timestamp 1707688321
transform 1 0 1924 0 1 1475
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_0
timestamp 1707688321
transform 0 -1 2119 -1 0 929
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_1
timestamp 1707688321
transform 0 -1 1020 -1 0 438
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_2
timestamp 1707688321
transform 0 -1 2119 -1 0 1199
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_3
timestamp 1707688321
transform 0 -1 1404 -1 0 775
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_4
timestamp 1707688321
transform 0 -1 1330 -1 0 775
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_5
timestamp 1707688321
transform -1 0 1487 0 1 1168
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_6
timestamp 1707688321
transform -1 0 278 0 1 821
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_7
timestamp 1707688321
transform -1 0 1887 0 1 955
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_8
timestamp 1707688321
transform -1 0 248 0 1 1555
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_9
timestamp 1707688321
transform -1 0 147 0 -1 1084
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_10
timestamp 1707688321
transform -1 0 1883 0 -1 1063
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_11
timestamp 1707688321
transform -1 0 193 0 -1 1009
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_12
timestamp 1707688321
transform -1 0 389 0 -1 697
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_13
timestamp 1707688321
transform -1 0 1663 0 -1 989
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_14
timestamp 1707688321
transform 1 0 1545 0 -1 1850
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_15
timestamp 1707688321
transform 1 0 1920 0 -1 1850
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_16
timestamp 1707688321
transform 1 0 1685 0 -1 1583
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_17
timestamp 1707688321
transform 1 0 484 0 -1 935
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_18
timestamp 1707688321
transform 1 0 461 0 -1 1205
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_19
timestamp 1707688321
transform 1 0 580 0 1 975
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_20
timestamp 1707688321
transform 1 0 870 0 1 1605
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_21
timestamp 1707688321
transform 1 0 1405 0 1 821
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_22
timestamp 1707688321
transform 1 0 124 0 1 1475
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_23
timestamp 1707688321
transform 1 0 1815 0 1 821
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_24
timestamp 1707688321
transform 1 0 1030 0 1 821
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_25
timestamp 1707688321
transform 1 0 1145 0 1 1816
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_26
timestamp 1707688321
transform 1 0 605 0 1 1816
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_27
timestamp 1707688321
transform 1 0 1241 0 1 1605
box 0 0 1 1
use L1M1_CDNS_5246887918590  L1M1_CDNS_5246887918590_0
timestamp 1707688321
transform 0 -1 251 -1 0 1429
box 0 0 1 1
use L1M1_CDNS_5246887918590  L1M1_CDNS_5246887918590_1
timestamp 1707688321
transform 0 -1 991 -1 0 2074
box 0 0 1 1
use L1M1_CDNS_5246887918590  L1M1_CDNS_5246887918590_2
timestamp 1707688321
transform 0 -1 523 -1 0 1429
box 0 0 1 1
use L1M1_CDNS_5246887918590  L1M1_CDNS_5246887918590_3
timestamp 1707688321
transform 0 -1 1487 -1 0 1429
box 0 0 1 1
use L1M1_CDNS_5246887918590  L1M1_CDNS_5246887918590_4
timestamp 1707688321
transform 0 1 295 1 0 1896
box 0 0 1 1
use L1M1_CDNS_5246887918590  L1M1_CDNS_5246887918590_5
timestamp 1707688321
transform 0 1 -17 1 0 1896
box 0 0 1 1
use L1M1_CDNS_5246887918590  L1M1_CDNS_5246887918590_6
timestamp 1707688321
transform 0 -1 1927 1 0 1251
box 0 0 1 1
use L1M1_CDNS_5246887918590  L1M1_CDNS_5246887918590_7
timestamp 1707688321
transform 0 -1 459 1 0 102
box 0 0 1 1
use L1M1_CDNS_5246887918590  L1M1_CDNS_5246887918590_8
timestamp 1707688321
transform 0 -1 17 1 0 102
box 0 0 1 1
use L1M1_CDNS_5246887918590  L1M1_CDNS_5246887918590_9
timestamp 1707688321
transform 0 -1 1743 1 0 1251
box 0 0 1 1
use L1M1_CDNS_5246887918590  L1M1_CDNS_5246887918590_10
timestamp 1707688321
transform 0 -1 751 1 0 102
box 0 0 1 1
use L1M1_CDNS_52468879185193  L1M1_CDNS_52468879185193_0
timestamp 1707688321
transform 1 0 -17 0 1 2192
box 0 0 1 1
use L1M1_CDNS_52468879185196  L1M1_CDNS_52468879185196_0
timestamp 1707688321
transform -1 0 952 0 1 1049
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_0
timestamp 1707688321
transform 0 -1 1756 -1 0 787
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_1
timestamp 1707688321
transform 0 -1 1336 -1 0 787
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_2
timestamp 1707688321
transform 0 -1 1416 -1 0 787
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_3
timestamp 1707688321
transform 0 1 450 -1 0 448
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_4
timestamp 1707688321
transform -1 0 658 0 -1 1095
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_5
timestamp 1707688321
transform -1 0 578 0 -1 1211
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_6
timestamp 1707688321
transform -1 0 578 0 -1 941
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_7
timestamp 1707688321
transform 1 0 1364 0 1 1599
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_8
timestamp 1707688321
transform 1 0 1284 0 1 1804
box 0 0 1 1
use M1M2_CDNS_52468879185199  M1M2_CDNS_52468879185199_0
timestamp 1707688321
transform -1 0 658 0 -1 787
box 0 0 1 1
use M1M2_CDNS_52468879185203  M1M2_CDNS_52468879185203_0
timestamp 1707688321
transform 0 -1 1756 -1 0 1435
box 0 0 1 1
use nfet_CDNS_52468879185411  nfet_CDNS_52468879185411_0
timestamp 1707688321
transform -1 0 206 0 -1 1268
box -79 -26 202 226
use nfet_CDNS_52468879185412  nfet_CDNS_52468879185412_0
timestamp 1707688321
transform 1 0 262 0 -1 1268
box -82 -26 202 226
use nfet_CDNS_52468879185413  nfet_CDNS_52468879185413_0
timestamp 1707688321
transform -1 0 1729 0 -1 723
box -82 -26 199 626
use nfet_CDNS_52468879185414  nfet_CDNS_52468879185414_0
timestamp 1707688321
transform 1 0 1785 0 -1 723
box -82 -26 199 626
use nfet_CDNS_52468879185415  nfet_CDNS_52468879185415_0
timestamp 1707688321
transform -1 0 958 0 -1 1315
box -79 -26 370 226
use nfet_CDNS_52468879185415  nfet_CDNS_52468879185415_1
timestamp 1707688321
transform -1 0 1302 0 -1 1315
box -79 -26 370 226
use nfet_CDNS_52468879185416  nfet_CDNS_52468879185416_0
timestamp 1707688321
transform -1 0 1553 0 -1 723
box -79 -26 199 626
use nfet_CDNS_52468879185417  nfet_CDNS_52468879185417_0
timestamp 1707688321
transform -1 0 1267 0 -1 723
box -79 -26 199 626
use nfet_CDNS_524688791851155  nfet_CDNS_524688791851155_0
timestamp 1707688321
transform -1 0 1942 0 1 880
box -79 -26 535 176
use nfet_CDNS_524688791851156  nfet_CDNS_524688791851156_0
timestamp 1707688321
transform 1 0 650 0 -1 1967
box -79 -26 259 226
use nfet_CDNS_524688791851156  nfet_CDNS_524688791851156_1
timestamp 1707688321
transform 1 0 1122 0 1 1767
box -79 -26 259 226
use nfet_CDNS_524688791851157  nfet_CDNS_524688791851157_0
timestamp 1707688321
transform 1 0 650 0 1 1469
box -79 -26 731 226
use nfet_CDNS_524688791851157  nfet_CDNS_524688791851157_1
timestamp 1707688321
transform 1 0 650 0 1 2027
box -79 -26 731 226
use nfet_CDNS_524688791851158  nfet_CDNS_524688791851158_0
timestamp 1707688321
transform -1 0 1974 0 1 1234
box -82 -26 394 226
use pfet_CDNS_52468879185420  pfet_CDNS_52468879185420_0
timestamp 1707688321
transform -1 0 414 0 -1 718
box -119 -66 239 666
use pfet_CDNS_52468879185421  pfet_CDNS_52468879185421_0
timestamp 1707688321
transform 1 0 470 0 -1 718
box -119 -66 239 666
use pfet_CDNS_52468879185422  pfet_CDNS_52468879185422_0
timestamp 1707688321
transform 1 0 28 0 -1 268
box -119 -66 219 216
use pfet_CDNS_52468879185424  pfet_CDNS_52468879185424_0
timestamp 1707688321
transform 1 0 28 0 -1 718
box -119 -66 219 216
use pfet_CDNS_52468879185442  pfet_CDNS_52468879185442_0
timestamp 1707688321
transform -1 0 284 0 -1 2145
box -119 -66 219 666
use pfet_CDNS_52468879185442  pfet_CDNS_52468879185442_1
timestamp 1707688321
transform 1 0 28 0 -1 2145
box -119 -66 219 666
use pfet_CDNS_524688791851159  pfet_CDNS_524688791851159_0
timestamp 1707688321
transform -1 0 1698 0 -1 2162
box -92 -36 125 636
use pfet_CDNS_524688791851159  pfet_CDNS_524688791851159_1
timestamp 1707688321
transform 1 0 1754 0 -1 2162
box -92 -36 125 636
use PYL1_CDNS_5246887918526  PYL1_CDNS_5246887918526_0
timestamp 1707688321
transform 1 0 1916 0 -1 1166
box 0 0 1 1
use PYL1_CDNS_5246887918526  PYL1_CDNS_5246887918526_1
timestamp 1707688321
transform 1 0 264 0 1 906
box 0 0 1 1
use PYL1_CDNS_5246887918562  PYL1_CDNS_5246887918562_0
timestamp 1707688321
transform 0 1 1875 1 0 2154
box 0 0 1 1
use PYL1_CDNS_5246887918562  PYL1_CDNS_5246887918562_1
timestamp 1707688321
transform 0 1 73 1 0 933
box 0 0 1 1
use PYL1_CDNS_5246887918562  PYL1_CDNS_5246887918562_2
timestamp 1707688321
transform 0 1 456 1 0 0
box 0 0 1 1
use PYL1_CDNS_5246887918562  PYL1_CDNS_5246887918562_3
timestamp 1707688321
transform 0 1 456 1 0 750
box 0 0 1 1
use PYL1_CDNS_5246887918562  PYL1_CDNS_5246887918562_4
timestamp 1707688321
transform 0 -1 1919 1 0 0
box 0 0 1 1
use PYL1_CDNS_5246887918562  PYL1_CDNS_5246887918562_5
timestamp 1707688321
transform 0 -1 1729 1 0 0
box 0 0 1 1
use PYL1_CDNS_5246887918562  PYL1_CDNS_5246887918562_6
timestamp 1707688321
transform 0 -1 1935 1 0 791
box 0 0 1 1
use PYL1_CDNS_5246887918562  PYL1_CDNS_5246887918562_7
timestamp 1707688321
transform 0 -1 1679 1 0 791
box 0 0 1 1
use PYL1_CDNS_5246887918562  PYL1_CDNS_5246887918562_8
timestamp 1707688321
transform 1 0 1908 0 1 1475
box 0 0 1 1
use PYL1_CDNS_52468879185136  PYL1_CDNS_52468879185136_0
timestamp 1707688321
transform 0 1 28 1 0 1447
box 0 0 1 1
use PYL1_CDNS_52468879185309  PYL1_CDNS_52468879185309_0
timestamp 1707688321
transform 0 -1 1293 -1 0 1093
box 0 0 1 1
use PYL1_CDNS_52468879185309  PYL1_CDNS_52468879185309_1
timestamp 1707688321
transform 0 -1 952 -1 0 1093
box 0 0 1 1
use PYL1_CDNS_52468879185327  PYL1_CDNS_52468879185327_0
timestamp 1707688321
transform 0 -1 1553 1 0 0
box 0 0 1 1
use PYL1_CDNS_52468879185444  PYL1_CDNS_52468879185444_0
timestamp 1707688321
transform 0 -1 1007 -1 0 1968
box 0 0 1 1
<< labels >>
flabel comment s 1481 1063 1481 1063 0 FreeSans 200 180 0 0 in_i_n
flabel comment s 824 1070 824 1070 0 FreeSans 200 180 0 0 in_i
flabel comment s 1728 886 1728 886 0 FreeSans 200 0 0 0 vgnd
flabel comment s 1932 628 1932 628 0 FreeSans 200 180 0 0 fbk
flabel comment s 1357 994 1357 994 0 FreeSans 200 0 0 0 fbk_n
flabel comment s 254 2193 254 2193 0 FreeSans 200 180 0 0 lv_net
flabel comment s 1770 1674 1770 1674 0 FreeSans 200 180 0 0 in_i
flabel comment s 626 1069 626 1069 0 FreeSans 200 0 0 0 out_h
flabel comment s 338 680 338 680 0 FreeSans 200 0 0 0 out_h_n
flabel comment s 1658 0 1658 0 0 FreeSans 200 0 0 0 set_h
flabel comment s 1867 0 1867 0 0 FreeSans 200 0 0 0 rst_h
flabel comment s 1738 630 1738 630 0 FreeSans 200 180 0 0 vgnd
flabel comment s 159 1459 159 1459 0 FreeSans 200 180 0 0 in_dis
flabel comment s 1579 628 1579 628 0 FreeSans 200 180 0 0 fbk_n
flabel comment s 1924 1824 1924 1824 0 FreeSans 200 0 0 0 in_i_n
flabel comment s 2024 1060 2024 1060 0 FreeSans 200 0 0 0 in
flabel comment s 1348 13 1348 13 0 FreeSans 200 180 0 0 hld_h_n
flabel comment s 428 1370 428 1370 0 FreeSans 200 180 0 0 vgnd
flabel comment s 1356 840 1356 840 0 FreeSans 200 0 0 0 fbk
flabel comment s 1562 1345 1562 1345 0 FreeSans 200 180 0 0 in_i_n
flabel comment s 398 1560 398 1560 0 FreeSans 200 0 0 0 virt_pwr
flabel metal1 s 0 1884 34 2086 3 FreeSans 400 0 0 0 vpwr
port 4 nsew
flabel metal1 s 1883 1884 1917 2086 3 FreeSans 400 180 0 0 vpwr
port 4 nsew
flabel metal1 s 0 320 34 450 3 FreeSans 400 0 0 0 vgnd
port 3 nsew
flabel metal1 s 196 1475 230 1509 0 FreeSans 400 0 0 0 in_dis
port 8 nsew
flabel metal1 s 2068 2114 2102 2232 7 FreeSans 400 0 0 0 vpb
port 2 nsew
flabel metal1 s 2068 1239 2102 1441 7 FreeSans 400 0 0 0 vgnd
port 3 nsew
flabel metal1 s 0 1239 34 1441 3 FreeSans 400 0 0 0 vgnd
port 3 nsew
flabel metal1 s 0 90 34 292 3 FreeSans 400 0 0 0 vcc_io
port 5 nsew
flabel metal1 s 321 663 355 697 0 FreeSans 200 0 0 0 out_h_n
port 6 nsew
flabel metal1 s 213 1492 213 1492 0 FreeSans 400 0 0 0 in_dis
flabel metal1 s 1969 1049 2004 1083 0 FreeSans 200 0 0 0 in
port 7 nsew
flabel metal1 s 0 2114 34 2232 3 FreeSans 400 0 0 0 vpb
port 2 nsew
flabel metal1 s 2068 90 2102 292 7 FreeSans 400 0 0 0 vcc_io
port 5 nsew
flabel locali s 1333 16 1367 49 0 FreeSans 200 180 0 0 hld_h_n
port 9 nsew
flabel locali s 1644 16 1678 50 0 FreeSans 400 180 0 0 set_h
port 10 nsew
flabel locali s 1835 16 1869 50 0 FreeSans 400 180 0 0 rst_h
port 11 nsew
flabel metal2 s 611 1054 641 1084 0 FreeSans 200 0 0 0 out_h
port 12 nsew
<< properties >>
string GDS_END 79640296
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 79615812
string path 9.075 55.900 -0.175 55.900 
<< end >>
