magic
tech sky130A
magscale 1 2
timestamp 1707688321
<< dnwell >>
rect 1900 26767 14000 39887
rect 4057 14468 14000 26767
rect 1931 8801 14000 14468
rect 10500 4585 14000 8801
rect 2365 235 14000 4585
<< nwell >>
rect 1767 39628 14086 40000
rect 1767 26975 2139 39628
rect 1767 26603 4265 26975
rect 3893 14629 4265 26603
rect 1767 14257 4265 14629
rect 1767 9007 2139 14257
rect 13714 9007 14086 39628
rect 1767 8635 14086 9007
rect 10364 8524 14086 8635
rect 10406 8224 14086 8524
rect 880 5785 9252 7586
rect 10406 6279 10706 8224
rect 13533 6279 14086 8224
rect 10406 5979 14086 6279
rect 10364 5623 14193 5979
rect 10364 4683 11073 5623
rect 2267 4379 11073 4683
rect 2267 441 2571 4379
rect 13794 441 14193 5623
rect 2267 137 14193 441
<< pwell >>
rect 2199 39346 13654 39568
rect 2199 27259 2421 39346
rect 2199 27037 4558 27259
rect 4336 14195 4558 27037
rect 2199 13973 4558 14195
rect 2199 9292 2421 13973
rect 13432 9292 13654 39346
rect 2199 9070 13654 9292
rect 594 7717 9662 7939
rect 594 5628 816 7717
rect 9440 5628 9662 7717
rect 10766 8056 13454 8142
rect 10766 6427 10852 8056
rect 13368 6427 13454 8056
rect 10766 6341 13454 6427
rect 594 5406 9662 5628
rect 11344 5477 12582 5563
rect 11344 4267 11430 5477
rect 12496 4267 12582 5477
<< mvpsubdiff >>
rect 2225 39508 2306 39542
rect 2340 39508 2374 39542
rect 2225 39474 2374 39508
rect 2327 39440 2374 39474
rect 13560 39458 13628 39542
rect 13560 39440 13594 39458
rect 2327 39406 2442 39440
rect 2395 39372 2442 39406
rect 13492 39424 13594 39440
rect 13492 39390 13628 39424
rect 13492 39372 13526 39390
rect 13458 39322 13526 39372
rect 2327 27233 2395 27268
rect 2327 27200 2361 27233
rect 2225 27166 2361 27200
rect 2259 27165 2361 27166
rect 4367 27199 4401 27233
rect 4435 27199 4532 27233
rect 4367 27165 4532 27199
rect 2259 27132 2293 27165
rect 2225 27063 2293 27132
rect 4367 27131 4430 27165
rect 4299 27097 4430 27131
rect 4299 27063 4362 27097
rect 4362 14169 4430 14211
rect 2225 14135 2322 14169
rect 2356 14135 2390 14169
rect 2225 14101 2390 14135
rect 4396 14143 4430 14169
rect 4396 14109 4532 14143
rect 4396 14101 4498 14109
rect 2327 14067 2390 14101
rect 4464 14075 4498 14101
rect 2327 14033 2458 14067
rect 2395 13999 2458 14033
rect 4464 13999 4532 14075
rect 2225 11659 2395 11755
rect 2327 9266 2395 9313
rect 2327 9245 2361 9266
rect 2225 9211 2361 9245
rect 2259 9198 2361 9211
rect 13411 9232 13458 9266
rect 13411 9198 13526 9232
rect 2259 9177 2293 9198
rect 2225 9096 2293 9177
rect 13479 9164 13526 9198
rect 13479 9130 13628 9164
rect 13479 9096 13513 9130
rect 13547 9096 13628 9130
rect 620 7879 694 7913
rect 728 7879 762 7913
rect 620 7845 762 7879
rect 722 7811 762 7845
rect 9568 7811 9636 7913
rect 722 7777 830 7811
rect 790 7743 830 7777
rect 9500 7778 9636 7811
rect 9500 7744 9602 7778
rect 9500 7743 9636 7744
rect 9466 7710 9636 7743
rect 9466 7642 9534 7710
rect 620 5631 790 5703
rect 654 5597 688 5631
rect 722 5602 790 5631
rect 722 5597 756 5602
rect 620 5563 756 5597
rect 654 5534 756 5563
rect 9426 5568 9466 5602
rect 10792 8082 10878 8116
rect 10912 8082 10946 8116
rect 10980 8082 11014 8116
rect 11048 8082 11082 8116
rect 11116 8082 11150 8116
rect 11184 8082 11218 8116
rect 11252 8082 11286 8116
rect 11320 8082 11354 8116
rect 11388 8082 11422 8116
rect 11456 8082 11490 8116
rect 11524 8082 11558 8116
rect 11592 8082 11626 8116
rect 11660 8082 11694 8116
rect 11728 8082 11762 8116
rect 11796 8082 11830 8116
rect 11864 8082 11898 8116
rect 11932 8082 11966 8116
rect 12000 8082 12034 8116
rect 12068 8082 12102 8116
rect 12136 8082 12170 8116
rect 12204 8082 12238 8116
rect 12272 8082 12306 8116
rect 12340 8082 12374 8116
rect 12408 8082 12442 8116
rect 12476 8082 12510 8116
rect 12544 8082 12578 8116
rect 12612 8082 12646 8116
rect 12680 8082 12714 8116
rect 12748 8082 12782 8116
rect 12816 8082 12850 8116
rect 12884 8082 12918 8116
rect 12952 8082 12986 8116
rect 13020 8082 13054 8116
rect 13088 8082 13122 8116
rect 13156 8082 13190 8116
rect 13224 8082 13258 8116
rect 13292 8082 13326 8116
rect 13360 8082 13428 8116
rect 10792 8048 10826 8082
rect 10792 7980 10826 8014
rect 13394 8033 13428 8082
rect 10792 7912 10826 7946
rect 13394 7965 13428 7999
rect 10792 7844 10826 7878
rect 10792 7776 10826 7810
rect 10792 7708 10826 7742
rect 10792 7640 10826 7674
rect 10792 7572 10826 7606
rect 10792 7504 10826 7538
rect 10792 7436 10826 7470
rect 10792 7368 10826 7402
rect 10792 7300 10826 7334
rect 10792 7232 10826 7266
rect 10792 7164 10826 7198
rect 10792 7096 10826 7130
rect 10792 7028 10826 7062
rect 10792 6960 10826 6994
rect 10792 6892 10826 6926
rect 10792 6824 10826 6858
rect 10792 6756 10826 6790
rect 10792 6688 10826 6722
rect 10792 6620 10826 6654
rect 10792 6552 10826 6586
rect 10792 6401 10826 6518
rect 13394 7897 13428 7931
rect 13394 7829 13428 7863
rect 13394 7761 13428 7795
rect 13394 7693 13428 7727
rect 13394 7625 13428 7659
rect 13394 7557 13428 7591
rect 13394 7489 13428 7523
rect 13394 7421 13428 7455
rect 13394 7353 13428 7387
rect 13394 7285 13428 7319
rect 13394 7217 13428 7251
rect 13394 7149 13428 7183
rect 13394 7081 13428 7115
rect 13394 7013 13428 7047
rect 13394 6945 13428 6979
rect 13394 6877 13428 6911
rect 13394 6809 13428 6843
rect 13394 6741 13428 6775
rect 13394 6673 13428 6707
rect 13394 6605 13428 6639
rect 13394 6537 13428 6571
rect 13394 6469 13428 6503
rect 13394 6401 13428 6435
rect 10792 6367 10860 6401
rect 10894 6367 10928 6401
rect 10962 6367 10996 6401
rect 11030 6367 11064 6401
rect 11098 6367 11132 6401
rect 11166 6367 11200 6401
rect 11234 6367 11268 6401
rect 11302 6367 11336 6401
rect 11370 6367 11404 6401
rect 11438 6367 11472 6401
rect 11506 6367 11540 6401
rect 11574 6367 11608 6401
rect 11642 6367 11676 6401
rect 11710 6367 11744 6401
rect 11778 6367 11812 6401
rect 11846 6367 11880 6401
rect 11914 6367 11948 6401
rect 11982 6367 12016 6401
rect 12050 6367 12084 6401
rect 12118 6367 12152 6401
rect 12186 6367 12220 6401
rect 12254 6367 12288 6401
rect 12322 6367 12356 6401
rect 12390 6367 12424 6401
rect 12458 6367 12492 6401
rect 12526 6367 12560 6401
rect 12594 6367 12628 6401
rect 12662 6367 12696 6401
rect 12730 6367 12764 6401
rect 12798 6367 12832 6401
rect 12866 6367 12900 6401
rect 12934 6367 12968 6401
rect 13002 6367 13036 6401
rect 13070 6367 13104 6401
rect 13138 6367 13172 6401
rect 13206 6367 13240 6401
rect 13274 6367 13308 6401
rect 13342 6367 13428 6401
rect 9426 5534 9534 5568
rect 654 5529 688 5534
rect 620 5432 688 5529
rect 9494 5500 9534 5534
rect 9494 5466 9636 5500
rect 9494 5432 9528 5466
rect 9562 5432 9636 5466
rect 11370 5503 11468 5537
rect 11502 5503 11536 5537
rect 11570 5503 11604 5537
rect 11638 5503 11672 5537
rect 11706 5503 11740 5537
rect 11774 5503 11808 5537
rect 11842 5503 11876 5537
rect 11910 5503 11944 5537
rect 11978 5503 12012 5537
rect 12046 5503 12080 5537
rect 12114 5503 12148 5537
rect 12182 5503 12216 5537
rect 12250 5503 12284 5537
rect 12318 5503 12352 5537
rect 12386 5503 12420 5537
rect 12454 5503 12488 5537
rect 11370 5449 11404 5503
rect 11370 5381 11404 5415
rect 11370 5313 11404 5347
rect 11370 5245 11404 5279
rect 11370 5177 11404 5211
rect 11370 5109 11404 5143
rect 11370 5041 11404 5075
rect 11370 4973 11404 5007
rect 11370 4905 11404 4939
rect 11370 4837 11404 4871
rect 11370 4769 11404 4803
rect 11370 4701 11404 4735
rect 11370 4633 11404 4667
rect 11370 4565 11404 4599
rect 11370 4497 11404 4531
rect 11370 4429 11404 4463
rect 12522 5449 12556 5537
rect 12522 5381 12556 5415
rect 12522 5313 12556 5347
rect 12522 5245 12556 5279
rect 12522 5177 12556 5211
rect 12522 5109 12556 5143
rect 12522 5041 12556 5075
rect 12522 4973 12556 5007
rect 12522 4905 12556 4939
rect 12522 4837 12556 4871
rect 12522 4769 12556 4803
rect 12522 4701 12556 4735
rect 12522 4633 12556 4667
rect 12522 4565 12556 4599
rect 12522 4497 12556 4531
rect 12522 4429 12556 4463
rect 11370 4361 11404 4395
rect 12522 4361 12556 4395
rect 11370 4293 11404 4327
rect 12522 4293 12556 4327
<< mvnsubdiff >>
rect 1834 39899 1949 39933
rect 1983 39899 2017 39933
rect 1834 39865 2017 39899
rect 1936 39831 2017 39865
rect 13951 39831 14019 39933
rect 1936 39797 2085 39831
rect 2004 39763 2085 39797
rect 13883 39812 14019 39831
rect 13883 39778 13985 39812
rect 13883 39763 14019 39778
rect 2004 39729 2153 39763
rect 2072 39695 2153 39729
rect 13815 39744 14019 39763
rect 13815 39695 13917 39744
rect 13781 39676 13917 39695
rect 13781 39608 13849 39676
rect 2004 26911 2072 26979
rect 1936 26908 2072 26911
rect 1936 26843 2038 26908
rect 1834 26840 2038 26843
rect 4044 26874 4078 26908
rect 4112 26874 4198 26908
rect 4044 26840 4198 26874
rect 1834 26809 1970 26840
rect 1868 26775 1970 26809
rect 4044 26806 4096 26840
rect 1834 26772 1970 26775
rect 3976 26772 4096 26806
rect 1834 26670 1902 26772
rect 3976 26738 4028 26772
rect 3908 26704 4028 26738
rect 3908 26670 3960 26704
rect 3960 14566 4028 14634
rect 3960 14562 4096 14566
rect 1834 14528 1920 14562
rect 1954 14528 1988 14562
rect 1834 14494 1988 14528
rect 3994 14498 4096 14562
rect 3994 14494 4198 14498
rect 1936 14460 1988 14494
rect 4062 14464 4198 14494
rect 1936 14426 2056 14460
rect 4062 14430 4164 14464
rect 4062 14426 4198 14430
rect 2004 14392 2056 14426
rect 2004 14358 2124 14392
rect 2072 14324 2124 14358
rect 4130 14324 4198 14426
rect 1834 10746 2072 10856
rect 2004 8944 2072 9012
rect 1936 8940 2072 8944
rect 1936 8876 2038 8940
rect 1834 8872 2038 8876
rect 13700 8906 13781 8940
rect 13700 8872 13849 8906
rect 1834 8842 1970 8872
rect 1868 8808 1970 8842
rect 1834 8804 1970 8808
rect 13768 8838 13849 8872
rect 13768 8804 13917 8838
rect 1834 8702 1902 8804
rect 13836 8770 13917 8804
rect 13836 8736 14019 8770
rect 13836 8702 13870 8736
rect 13904 8702 14019 8736
rect 10473 8423 10604 8457
rect 10638 8423 10672 8457
rect 10706 8423 10740 8457
rect 10774 8423 10808 8457
rect 10842 8423 10876 8457
rect 10910 8423 10944 8457
rect 10978 8423 11012 8457
rect 11046 8423 11080 8457
rect 11114 8423 11148 8457
rect 11182 8423 11216 8457
rect 11250 8423 11284 8457
rect 11318 8423 11352 8457
rect 11386 8423 11420 8457
rect 11454 8423 11488 8457
rect 11522 8423 11556 8457
rect 11590 8423 11624 8457
rect 11658 8423 11692 8457
rect 11726 8423 11760 8457
rect 11794 8423 11828 8457
rect 11862 8423 11896 8457
rect 11930 8423 11964 8457
rect 11998 8423 12032 8457
rect 12066 8423 12100 8457
rect 12134 8423 12168 8457
rect 12202 8423 12236 8457
rect 12270 8423 12304 8457
rect 12338 8423 12372 8457
rect 12406 8423 12440 8457
rect 12474 8423 12508 8457
rect 12542 8423 12576 8457
rect 12610 8423 12644 8457
rect 12678 8423 12712 8457
rect 12746 8423 12780 8457
rect 12814 8423 12848 8457
rect 12882 8423 12916 8457
rect 12950 8423 12984 8457
rect 13018 8423 13052 8457
rect 13086 8423 13120 8457
rect 13154 8423 13188 8457
rect 13222 8423 13256 8457
rect 13290 8423 13324 8457
rect 13358 8423 13392 8457
rect 13426 8423 13460 8457
rect 13494 8423 13528 8457
rect 13562 8423 13596 8457
rect 13630 8423 13664 8457
rect 13698 8423 13766 8457
rect 10473 8389 13766 8423
rect 10507 8355 13766 8389
rect 10473 8325 13766 8355
rect 10473 8321 10605 8325
rect 10507 8291 10605 8321
rect 10639 8291 10676 8325
rect 10710 8291 10744 8325
rect 10778 8291 10812 8325
rect 10846 8291 10880 8325
rect 10914 8291 10948 8325
rect 10982 8291 11016 8325
rect 11050 8291 11084 8325
rect 11118 8291 11152 8325
rect 11186 8291 11220 8325
rect 11254 8291 11288 8325
rect 11322 8291 11356 8325
rect 11390 8291 11424 8325
rect 11458 8291 11492 8325
rect 11526 8291 11560 8325
rect 11594 8291 11628 8325
rect 11662 8291 11696 8325
rect 11730 8291 11764 8325
rect 11798 8291 11832 8325
rect 11866 8291 11900 8325
rect 11934 8291 11968 8325
rect 12002 8291 12036 8325
rect 12070 8291 12104 8325
rect 12138 8291 12172 8325
rect 12206 8291 12240 8325
rect 12274 8291 12308 8325
rect 12342 8291 12376 8325
rect 12410 8291 12444 8325
rect 12478 8291 12512 8325
rect 12546 8291 12580 8325
rect 12614 8291 12648 8325
rect 12682 8291 12716 8325
rect 12750 8291 12784 8325
rect 12818 8291 12852 8325
rect 12886 8291 12920 8325
rect 12954 8291 12988 8325
rect 13022 8291 13056 8325
rect 13090 8291 13124 8325
rect 13158 8291 13192 8325
rect 13226 8291 13260 8325
rect 13294 8291 13328 8325
rect 13362 8291 13396 8325
rect 13430 8291 13464 8325
rect 13498 8291 13532 8325
rect 13566 8291 13600 8325
rect 13634 8324 13766 8325
rect 13634 8291 13732 8324
rect 10507 8287 10639 8291
rect 10473 8257 10639 8287
rect 10473 8253 10605 8257
rect 10507 8223 10605 8253
rect 10507 8219 10639 8223
rect 10473 8189 10639 8219
rect 10473 8185 10605 8189
rect 10507 8155 10605 8185
rect 10507 8151 10639 8155
rect 10473 8121 10639 8151
rect 10473 8117 10605 8121
rect 10507 8087 10605 8117
rect 13600 8290 13732 8291
rect 13600 8256 13766 8290
rect 13600 8252 13732 8256
rect 13634 8222 13732 8252
rect 13634 8218 13766 8222
rect 13600 8188 13766 8218
rect 13600 8184 13732 8188
rect 13634 8154 13732 8184
rect 13634 8150 13766 8154
rect 13600 8120 13766 8150
rect 13600 8116 13732 8120
rect 10507 8083 10639 8087
rect 10473 8053 10639 8083
rect 10473 8049 10605 8053
rect 10507 8019 10605 8049
rect 10507 8015 10639 8019
rect 10473 7985 10639 8015
rect 10473 7981 10605 7985
rect 10507 7951 10605 7981
rect 10507 7947 10639 7951
rect 10473 7917 10639 7947
rect 10473 7913 10605 7917
rect 947 7485 1059 7519
rect 1093 7485 1127 7519
rect 1161 7485 1195 7519
rect 1229 7485 1263 7519
rect 1297 7485 1331 7519
rect 1365 7485 1399 7519
rect 1433 7485 1467 7519
rect 1501 7485 1535 7519
rect 1569 7485 1603 7519
rect 1637 7485 1671 7519
rect 1705 7485 1739 7519
rect 1773 7485 1807 7519
rect 1841 7485 1875 7519
rect 1909 7485 1943 7519
rect 1977 7485 2011 7519
rect 2045 7485 2079 7519
rect 2113 7485 2147 7519
rect 2181 7485 2215 7519
rect 2249 7485 2283 7519
rect 2317 7485 2351 7519
rect 2385 7485 2419 7519
rect 2453 7485 2487 7519
rect 2521 7485 2555 7519
rect 2589 7485 2623 7519
rect 2657 7485 2691 7519
rect 2725 7485 2759 7519
rect 2793 7485 2827 7519
rect 2861 7485 2895 7519
rect 2929 7485 2963 7519
rect 2997 7485 3031 7519
rect 3065 7485 3099 7519
rect 3133 7485 3167 7519
rect 3201 7485 3235 7519
rect 3269 7485 3303 7519
rect 3337 7485 3371 7519
rect 3405 7485 3439 7519
rect 3473 7485 3507 7519
rect 3541 7485 3575 7519
rect 3609 7485 3643 7519
rect 3677 7485 3711 7519
rect 3745 7485 3779 7519
rect 3813 7485 3847 7519
rect 3881 7485 3915 7519
rect 3949 7485 3983 7519
rect 4017 7485 4051 7519
rect 4085 7485 4119 7519
rect 4153 7485 4187 7519
rect 4221 7485 4255 7519
rect 4289 7485 4323 7519
rect 4357 7485 4391 7519
rect 4425 7485 4459 7519
rect 4493 7485 4527 7519
rect 4561 7485 4595 7519
rect 4629 7485 4663 7519
rect 4697 7485 4731 7519
rect 4765 7485 4799 7519
rect 4833 7485 4867 7519
rect 4901 7485 4935 7519
rect 4969 7485 5003 7519
rect 5037 7485 5071 7519
rect 5105 7485 5139 7519
rect 5173 7485 5207 7519
rect 5241 7485 5275 7519
rect 5309 7485 5343 7519
rect 5377 7485 5411 7519
rect 5445 7485 5479 7519
rect 5513 7485 5547 7519
rect 5581 7485 5615 7519
rect 5649 7485 5683 7519
rect 5717 7485 5751 7519
rect 5785 7485 5819 7519
rect 5853 7485 5887 7519
rect 5921 7485 5955 7519
rect 5989 7485 6023 7519
rect 6057 7485 6091 7519
rect 6125 7485 6159 7519
rect 6193 7485 6227 7519
rect 6261 7485 6295 7519
rect 6329 7485 6363 7519
rect 6397 7485 6431 7519
rect 6465 7485 6499 7519
rect 6533 7485 6567 7519
rect 6601 7485 6635 7519
rect 6669 7485 6703 7519
rect 6737 7485 6771 7519
rect 6805 7485 6839 7519
rect 6873 7485 6907 7519
rect 6941 7485 6975 7519
rect 7009 7485 7043 7519
rect 7077 7485 7111 7519
rect 7145 7485 7179 7519
rect 7213 7485 7247 7519
rect 7281 7485 7315 7519
rect 7349 7485 7383 7519
rect 7417 7485 7451 7519
rect 7485 7485 7519 7519
rect 7553 7485 7587 7519
rect 7621 7485 7655 7519
rect 7689 7485 7723 7519
rect 7757 7485 7791 7519
rect 7825 7485 7859 7519
rect 7893 7485 7927 7519
rect 7961 7485 7995 7519
rect 8029 7485 8063 7519
rect 8097 7485 8131 7519
rect 8165 7485 8199 7519
rect 8233 7485 8267 7519
rect 8301 7485 8335 7519
rect 8369 7485 8403 7519
rect 8437 7485 8471 7519
rect 8505 7485 8539 7519
rect 8573 7485 8607 7519
rect 8641 7485 8675 7519
rect 8709 7485 8743 7519
rect 8777 7485 8811 7519
rect 8845 7485 8879 7519
rect 8913 7485 8947 7519
rect 8981 7485 9015 7519
rect 9049 7485 9083 7519
rect 9117 7485 9185 7519
rect 947 7451 981 7485
rect 947 7383 981 7417
rect 9151 7450 9185 7485
rect 947 7315 981 7349
rect 947 7247 981 7281
rect 947 7179 981 7213
rect 947 7111 981 7145
rect 947 7043 981 7077
rect 947 6975 981 7009
rect 947 6907 981 6941
rect 947 6839 981 6873
rect 947 6771 981 6805
rect 947 6703 981 6737
rect 947 6635 981 6669
rect 947 6567 981 6601
rect 947 6499 981 6533
rect 947 6431 981 6465
rect 947 6363 981 6397
rect 947 6295 981 6329
rect 947 6227 981 6261
rect 947 6159 981 6193
rect 947 6091 981 6125
rect 947 6023 981 6057
rect 947 5886 981 5989
rect 9151 7382 9185 7416
rect 9151 7314 9185 7348
rect 9151 7246 9185 7280
rect 9151 7178 9185 7212
rect 9151 7110 9185 7144
rect 9151 7042 9185 7076
rect 9151 6974 9185 7008
rect 9151 6906 9185 6940
rect 9151 6838 9185 6872
rect 9151 6770 9185 6804
rect 9151 6702 9185 6736
rect 9151 6634 9185 6668
rect 9151 6566 9185 6600
rect 9151 6498 9185 6532
rect 9151 6430 9185 6464
rect 9151 6362 9185 6396
rect 9151 6294 9185 6328
rect 9151 6226 9185 6260
rect 9151 6158 9185 6192
rect 9151 6090 9185 6124
rect 9151 6022 9185 6056
rect 9151 5954 9185 5988
rect 9151 5886 9185 5920
rect 947 5852 1015 5886
rect 1049 5852 1083 5886
rect 1117 5852 1151 5886
rect 1185 5852 1219 5886
rect 1253 5852 1287 5886
rect 1321 5852 1355 5886
rect 1389 5852 1423 5886
rect 1457 5852 1491 5886
rect 1525 5852 1559 5886
rect 1593 5852 1627 5886
rect 1661 5852 1695 5886
rect 1729 5852 1763 5886
rect 1797 5852 1831 5886
rect 1865 5852 1899 5886
rect 1933 5852 1967 5886
rect 2001 5852 2035 5886
rect 2069 5852 2103 5886
rect 2137 5852 2171 5886
rect 2205 5852 2239 5886
rect 2273 5852 2307 5886
rect 2341 5852 2375 5886
rect 2409 5852 2443 5886
rect 2477 5852 2511 5886
rect 2545 5852 2579 5886
rect 2613 5852 2647 5886
rect 2681 5852 2715 5886
rect 2749 5852 2783 5886
rect 2817 5852 2851 5886
rect 2885 5852 2919 5886
rect 2953 5852 2987 5886
rect 3021 5852 3055 5886
rect 3089 5852 3123 5886
rect 3157 5852 3191 5886
rect 3225 5852 3259 5886
rect 3293 5852 3327 5886
rect 3361 5852 3395 5886
rect 3429 5852 3463 5886
rect 3497 5852 3531 5886
rect 3565 5852 3599 5886
rect 3633 5852 3667 5886
rect 3701 5852 3735 5886
rect 3769 5852 3803 5886
rect 3837 5852 3871 5886
rect 3905 5852 3939 5886
rect 3973 5852 4007 5886
rect 4041 5852 4075 5886
rect 4109 5852 4143 5886
rect 4177 5852 4211 5886
rect 4245 5852 4279 5886
rect 4313 5852 4347 5886
rect 4381 5852 4415 5886
rect 4449 5852 4483 5886
rect 4517 5852 4551 5886
rect 4585 5852 4619 5886
rect 4653 5852 4687 5886
rect 4721 5852 4755 5886
rect 4789 5852 4823 5886
rect 4857 5852 4891 5886
rect 4925 5852 4959 5886
rect 4993 5852 5027 5886
rect 5061 5852 5095 5886
rect 5129 5852 5163 5886
rect 5197 5852 5231 5886
rect 5265 5852 5299 5886
rect 5333 5852 5367 5886
rect 5401 5852 5435 5886
rect 5469 5852 5503 5886
rect 5537 5852 5571 5886
rect 5605 5852 5639 5886
rect 5673 5852 5707 5886
rect 5741 5852 5775 5886
rect 5809 5852 5843 5886
rect 5877 5852 5911 5886
rect 5945 5852 5979 5886
rect 6013 5852 6047 5886
rect 6081 5852 6115 5886
rect 6149 5852 6183 5886
rect 6217 5852 6251 5886
rect 6285 5852 6319 5886
rect 6353 5852 6387 5886
rect 6421 5852 6455 5886
rect 6489 5852 6523 5886
rect 6557 5852 6591 5886
rect 6625 5852 6659 5886
rect 6693 5852 6727 5886
rect 6761 5852 6795 5886
rect 6829 5852 6863 5886
rect 6897 5852 6931 5886
rect 6965 5852 6999 5886
rect 7033 5852 7067 5886
rect 7101 5852 7135 5886
rect 7169 5852 7203 5886
rect 7237 5852 7271 5886
rect 7305 5852 7339 5886
rect 7373 5852 7407 5886
rect 7441 5852 7475 5886
rect 7509 5852 7543 5886
rect 7577 5852 7611 5886
rect 7645 5852 7679 5886
rect 7713 5852 7747 5886
rect 7781 5852 7815 5886
rect 7849 5852 7883 5886
rect 7917 5852 7951 5886
rect 7985 5852 8019 5886
rect 8053 5852 8087 5886
rect 8121 5852 8155 5886
rect 8189 5852 8223 5886
rect 8257 5852 8291 5886
rect 8325 5852 8359 5886
rect 8393 5852 8427 5886
rect 8461 5852 8495 5886
rect 8529 5852 8563 5886
rect 8597 5852 8631 5886
rect 8665 5852 8699 5886
rect 8733 5852 8767 5886
rect 8801 5852 8835 5886
rect 8869 5852 8903 5886
rect 8937 5852 8971 5886
rect 9005 5852 9039 5886
rect 9073 5852 9185 5886
rect 10507 7883 10605 7913
rect 10507 7879 10639 7883
rect 10473 7849 10639 7879
rect 10473 7845 10605 7849
rect 10507 7815 10605 7845
rect 10507 7811 10639 7815
rect 10473 7781 10639 7811
rect 10473 7777 10605 7781
rect 10507 7747 10605 7777
rect 10507 7743 10639 7747
rect 10473 7713 10639 7743
rect 10473 7709 10605 7713
rect 10507 7679 10605 7709
rect 10507 7675 10639 7679
rect 10473 7645 10639 7675
rect 10473 7641 10605 7645
rect 10507 7611 10605 7641
rect 10507 7607 10639 7611
rect 10473 7577 10639 7607
rect 10473 7573 10605 7577
rect 10507 7543 10605 7573
rect 10507 7539 10639 7543
rect 10473 7509 10639 7539
rect 10473 7505 10605 7509
rect 10507 7475 10605 7505
rect 10507 7471 10639 7475
rect 10473 7441 10639 7471
rect 10473 7437 10605 7441
rect 10507 7407 10605 7437
rect 10507 7403 10639 7407
rect 10473 7373 10639 7403
rect 10473 7369 10605 7373
rect 10507 7339 10605 7369
rect 10507 7335 10639 7339
rect 10473 7305 10639 7335
rect 10473 7301 10605 7305
rect 10507 7271 10605 7301
rect 10507 7267 10639 7271
rect 10473 7237 10639 7267
rect 10473 7233 10605 7237
rect 10507 7203 10605 7233
rect 10507 7199 10639 7203
rect 10473 7169 10639 7199
rect 10473 7165 10605 7169
rect 10507 7135 10605 7165
rect 10507 7131 10639 7135
rect 10473 7101 10639 7131
rect 10473 7097 10605 7101
rect 10507 7067 10605 7097
rect 10507 7063 10639 7067
rect 10473 7033 10639 7063
rect 10473 7029 10605 7033
rect 10507 6999 10605 7029
rect 10507 6995 10639 6999
rect 10473 6965 10639 6995
rect 10473 6961 10605 6965
rect 10507 6931 10605 6961
rect 10507 6927 10639 6931
rect 10473 6897 10639 6927
rect 10473 6893 10605 6897
rect 10507 6863 10605 6893
rect 10507 6859 10639 6863
rect 10473 6829 10639 6859
rect 10473 6825 10605 6829
rect 10507 6795 10605 6825
rect 10507 6791 10639 6795
rect 10473 6761 10639 6791
rect 10473 6757 10605 6761
rect 10507 6727 10605 6757
rect 10507 6723 10639 6727
rect 10473 6693 10639 6723
rect 10473 6689 10605 6693
rect 10507 6659 10605 6689
rect 10507 6655 10639 6659
rect 10473 6625 10639 6655
rect 10473 6621 10605 6625
rect 10507 6591 10605 6621
rect 10507 6587 10639 6591
rect 10473 6557 10639 6587
rect 10473 6553 10605 6557
rect 10507 6523 10605 6553
rect 10507 6519 10639 6523
rect 10473 6489 10639 6519
rect 10473 6485 10605 6489
rect 10507 6455 10605 6485
rect 10507 6451 10639 6455
rect 10473 6329 10639 6451
rect 13634 8086 13732 8116
rect 13634 8082 13766 8086
rect 13600 8052 13766 8082
rect 13600 8048 13732 8052
rect 13634 8018 13732 8048
rect 13634 8014 13766 8018
rect 13600 7984 13766 8014
rect 13600 7980 13732 7984
rect 13634 7950 13732 7980
rect 13634 7946 13766 7950
rect 13600 7916 13766 7946
rect 13600 7912 13732 7916
rect 13634 7882 13732 7912
rect 13634 7878 13766 7882
rect 13600 7848 13766 7878
rect 13600 7844 13732 7848
rect 13634 7814 13732 7844
rect 13634 7810 13766 7814
rect 13600 7780 13766 7810
rect 13600 7776 13732 7780
rect 13634 7746 13732 7776
rect 13634 7742 13766 7746
rect 13600 7712 13766 7742
rect 13600 7708 13732 7712
rect 13634 7678 13732 7708
rect 13634 7674 13766 7678
rect 13600 7644 13766 7674
rect 13600 7640 13732 7644
rect 13634 7610 13732 7640
rect 13634 7606 13766 7610
rect 13600 7576 13766 7606
rect 13600 7572 13732 7576
rect 13634 7542 13732 7572
rect 13634 7538 13766 7542
rect 13600 7508 13766 7538
rect 13600 7504 13732 7508
rect 13634 7474 13732 7504
rect 13634 7470 13766 7474
rect 13600 7440 13766 7470
rect 13600 7436 13732 7440
rect 13634 7406 13732 7436
rect 13634 7402 13766 7406
rect 13600 7372 13766 7402
rect 13600 7368 13732 7372
rect 13634 7338 13732 7368
rect 13634 7334 13766 7338
rect 13600 7304 13766 7334
rect 13600 7300 13732 7304
rect 13634 7270 13732 7300
rect 13634 7266 13766 7270
rect 13600 7236 13766 7266
rect 13600 7232 13732 7236
rect 13634 7202 13732 7232
rect 13634 7198 13766 7202
rect 13600 7168 13766 7198
rect 13600 7164 13732 7168
rect 13634 7134 13732 7164
rect 13634 7130 13766 7134
rect 13600 7100 13766 7130
rect 13600 7096 13732 7100
rect 13634 7066 13732 7096
rect 13634 7062 13766 7066
rect 13600 7032 13766 7062
rect 13600 7028 13732 7032
rect 13634 6998 13732 7028
rect 13634 6994 13766 6998
rect 13600 6964 13766 6994
rect 13600 6960 13732 6964
rect 13634 6930 13732 6960
rect 13634 6926 13766 6930
rect 13600 6896 13766 6926
rect 13600 6892 13732 6896
rect 13634 6862 13732 6892
rect 13634 6858 13766 6862
rect 13600 6828 13766 6858
rect 13600 6824 13732 6828
rect 13634 6794 13732 6824
rect 13634 6790 13766 6794
rect 13600 6760 13766 6790
rect 13600 6756 13732 6760
rect 13634 6726 13732 6756
rect 13634 6722 13766 6726
rect 13600 6692 13766 6722
rect 13600 6688 13732 6692
rect 13634 6658 13732 6688
rect 13634 6654 13766 6658
rect 13600 6624 13766 6654
rect 13600 6620 13732 6624
rect 13634 6590 13732 6620
rect 13634 6586 13766 6590
rect 13600 6556 13766 6586
rect 13600 6552 13732 6556
rect 13634 6522 13732 6552
rect 13634 6518 13766 6522
rect 13600 6488 13766 6518
rect 13600 6484 13732 6488
rect 13634 6454 13732 6484
rect 13634 6450 13766 6454
rect 13600 6420 13766 6450
rect 13600 6416 13732 6420
rect 13634 6386 13732 6416
rect 13634 6382 13766 6386
rect 10507 6295 10605 6329
rect 10473 6261 10639 6295
rect 10507 6227 10639 6261
rect 10473 6212 10639 6227
rect 13600 6352 13766 6382
rect 13600 6348 13732 6352
rect 13634 6318 13732 6348
rect 13634 6314 13766 6318
rect 13600 6284 13766 6314
rect 13600 6280 13732 6284
rect 13634 6250 13732 6280
rect 13634 6246 13766 6250
rect 13600 6216 13766 6246
rect 13600 6212 13732 6216
rect 10473 6193 10605 6212
rect 10507 6178 10605 6193
rect 10639 6178 10673 6212
rect 10707 6178 10741 6212
rect 10775 6178 10809 6212
rect 10843 6178 10877 6212
rect 10911 6178 10945 6212
rect 10979 6178 11013 6212
rect 11047 6178 11081 6212
rect 11115 6178 11149 6212
rect 11183 6178 11217 6212
rect 11251 6178 11285 6212
rect 11319 6178 11353 6212
rect 11387 6178 11421 6212
rect 11455 6178 11489 6212
rect 11523 6178 11557 6212
rect 11591 6178 11625 6212
rect 11659 6178 11693 6212
rect 11727 6178 11761 6212
rect 11795 6178 11829 6212
rect 11863 6178 11897 6212
rect 11931 6178 11965 6212
rect 11999 6178 12033 6212
rect 12067 6178 12101 6212
rect 12135 6178 12169 6212
rect 12203 6178 12237 6212
rect 12271 6178 12305 6212
rect 12339 6178 12373 6212
rect 12407 6178 12441 6212
rect 12475 6178 12509 6212
rect 12543 6178 12577 6212
rect 12611 6178 12645 6212
rect 12679 6178 12713 6212
rect 12747 6178 12781 6212
rect 12815 6178 12849 6212
rect 12883 6178 12917 6212
rect 12951 6178 12985 6212
rect 13019 6178 13053 6212
rect 13087 6178 13121 6212
rect 13155 6178 13189 6212
rect 13223 6178 13257 6212
rect 13291 6178 13325 6212
rect 13359 6178 13393 6212
rect 13427 6178 13461 6212
rect 13495 6178 13529 6212
rect 13563 6178 13600 6212
rect 13634 6182 13732 6212
rect 13634 6178 13766 6182
rect 10507 6159 13766 6178
rect 10473 6148 13766 6159
rect 10473 6114 13732 6148
rect 10473 6080 13766 6114
rect 10473 6046 10541 6080
rect 10575 6046 10609 6080
rect 10643 6046 10677 6080
rect 10711 6046 10745 6080
rect 10779 6046 10813 6080
rect 10847 6046 10881 6080
rect 10915 6046 10949 6080
rect 10983 6046 11017 6080
rect 11051 6046 11085 6080
rect 11119 6046 11153 6080
rect 11187 6046 11221 6080
rect 11255 6046 11289 6080
rect 11323 6046 11357 6080
rect 11391 6046 11425 6080
rect 11459 6046 11493 6080
rect 11527 6046 11561 6080
rect 11595 6046 11629 6080
rect 11663 6046 11697 6080
rect 11731 6046 11765 6080
rect 11799 6046 11833 6080
rect 11867 6046 11901 6080
rect 11935 6046 11969 6080
rect 12003 6046 12037 6080
rect 12071 6046 12105 6080
rect 12139 6046 12173 6080
rect 12207 6046 12241 6080
rect 12275 6046 12309 6080
rect 12343 6046 12377 6080
rect 12411 6046 12445 6080
rect 12479 6046 12513 6080
rect 12547 6046 12581 6080
rect 12615 6046 12649 6080
rect 12683 6046 12717 6080
rect 12751 6046 12785 6080
rect 12819 6046 12853 6080
rect 12887 6046 12921 6080
rect 12955 6046 12989 6080
rect 13023 6046 13057 6080
rect 13091 6046 13125 6080
rect 13159 6046 13193 6080
rect 13227 6046 13261 6080
rect 13295 6046 13329 6080
rect 13363 6046 13397 6080
rect 13431 6046 13465 6080
rect 13499 6046 13533 6080
rect 13567 6046 13601 6080
rect 13635 6046 13766 6080
rect 10473 5860 13766 6046
rect 10836 5826 10964 5860
rect 10998 5826 11032 5860
rect 10836 5792 11032 5826
rect 10938 5758 11032 5792
rect 14058 5758 14126 5860
rect 10938 5724 11100 5758
rect 11006 5690 11100 5724
rect 13990 5746 14126 5758
rect 13990 5712 14092 5746
rect 13990 5690 14126 5712
rect 13956 5678 14126 5690
rect 13956 5610 14024 5678
rect 10836 4616 10904 4670
rect 2334 4582 2404 4616
rect 2438 4582 2472 4616
rect 2334 4548 2472 4582
rect 10870 4602 10904 4616
rect 10870 4568 11006 4602
rect 10870 4548 10972 4568
rect 2436 4514 2472 4548
rect 10938 4534 10972 4548
rect 2436 4480 2540 4514
rect 2504 4446 2540 4480
rect 10938 4446 11006 4534
rect 2334 390 2504 502
rect 2368 356 2402 390
rect 2436 374 2504 390
rect 2436 356 2470 374
rect 2334 322 2470 356
rect 2368 306 2470 322
rect 13860 340 13956 374
rect 13860 306 14024 340
rect 2368 288 2402 306
rect 2334 204 2402 288
rect 13928 272 14024 306
rect 13928 238 14126 272
rect 13928 204 13962 238
rect 13996 204 14126 238
<< mvpsubdiffcont >>
rect 2306 39508 2340 39542
rect 2225 39406 2327 39474
rect 2374 39440 13560 39542
rect 2225 27268 2395 39406
rect 2442 39372 13492 39440
rect 13594 39424 13628 39458
rect 13526 39322 13628 39390
rect 2225 27200 2327 27268
rect 2225 27132 2259 27166
rect 2361 27165 4367 27233
rect 4401 27199 4435 27233
rect 2293 27131 4367 27165
rect 2293 27063 4299 27131
rect 4430 27097 4532 27165
rect 4362 14211 4532 27097
rect 2322 14135 2356 14169
rect 2390 14101 4396 14169
rect 4430 14143 4532 14211
rect 2225 14033 2327 14101
rect 2390 14067 4464 14101
rect 4498 14075 4532 14109
rect 2225 11755 2395 14033
rect 2458 13999 4464 14067
rect 2225 9313 2395 11659
rect 2225 9245 2327 9313
rect 2225 9177 2259 9211
rect 2361 9198 13411 9266
rect 13458 9232 13628 39322
rect 2293 9096 13479 9198
rect 13526 9164 13628 9232
rect 13513 9096 13547 9130
rect 694 7879 728 7913
rect 620 7777 722 7845
rect 762 7811 9568 7913
rect 620 5703 790 7777
rect 830 7743 9500 7811
rect 9602 7744 9636 7778
rect 9534 7642 9636 7710
rect 620 5597 654 5631
rect 688 5597 722 5631
rect 620 5529 654 5563
rect 756 5534 9426 5602
rect 9466 5568 9636 7642
rect 10878 8082 10912 8116
rect 10946 8082 10980 8116
rect 11014 8082 11048 8116
rect 11082 8082 11116 8116
rect 11150 8082 11184 8116
rect 11218 8082 11252 8116
rect 11286 8082 11320 8116
rect 11354 8082 11388 8116
rect 11422 8082 11456 8116
rect 11490 8082 11524 8116
rect 11558 8082 11592 8116
rect 11626 8082 11660 8116
rect 11694 8082 11728 8116
rect 11762 8082 11796 8116
rect 11830 8082 11864 8116
rect 11898 8082 11932 8116
rect 11966 8082 12000 8116
rect 12034 8082 12068 8116
rect 12102 8082 12136 8116
rect 12170 8082 12204 8116
rect 12238 8082 12272 8116
rect 12306 8082 12340 8116
rect 12374 8082 12408 8116
rect 12442 8082 12476 8116
rect 12510 8082 12544 8116
rect 12578 8082 12612 8116
rect 12646 8082 12680 8116
rect 12714 8082 12748 8116
rect 12782 8082 12816 8116
rect 12850 8082 12884 8116
rect 12918 8082 12952 8116
rect 12986 8082 13020 8116
rect 13054 8082 13088 8116
rect 13122 8082 13156 8116
rect 13190 8082 13224 8116
rect 13258 8082 13292 8116
rect 13326 8082 13360 8116
rect 10792 8014 10826 8048
rect 10792 7946 10826 7980
rect 13394 7999 13428 8033
rect 10792 7878 10826 7912
rect 10792 7810 10826 7844
rect 10792 7742 10826 7776
rect 10792 7674 10826 7708
rect 10792 7606 10826 7640
rect 10792 7538 10826 7572
rect 10792 7470 10826 7504
rect 10792 7402 10826 7436
rect 10792 7334 10826 7368
rect 10792 7266 10826 7300
rect 10792 7198 10826 7232
rect 10792 7130 10826 7164
rect 10792 7062 10826 7096
rect 10792 6994 10826 7028
rect 10792 6926 10826 6960
rect 10792 6858 10826 6892
rect 10792 6790 10826 6824
rect 10792 6722 10826 6756
rect 10792 6654 10826 6688
rect 10792 6586 10826 6620
rect 10792 6518 10826 6552
rect 13394 7931 13428 7965
rect 13394 7863 13428 7897
rect 13394 7795 13428 7829
rect 13394 7727 13428 7761
rect 13394 7659 13428 7693
rect 13394 7591 13428 7625
rect 13394 7523 13428 7557
rect 13394 7455 13428 7489
rect 13394 7387 13428 7421
rect 13394 7319 13428 7353
rect 13394 7251 13428 7285
rect 13394 7183 13428 7217
rect 13394 7115 13428 7149
rect 13394 7047 13428 7081
rect 13394 6979 13428 7013
rect 13394 6911 13428 6945
rect 13394 6843 13428 6877
rect 13394 6775 13428 6809
rect 13394 6707 13428 6741
rect 13394 6639 13428 6673
rect 13394 6571 13428 6605
rect 13394 6503 13428 6537
rect 13394 6435 13428 6469
rect 10860 6367 10894 6401
rect 10928 6367 10962 6401
rect 10996 6367 11030 6401
rect 11064 6367 11098 6401
rect 11132 6367 11166 6401
rect 11200 6367 11234 6401
rect 11268 6367 11302 6401
rect 11336 6367 11370 6401
rect 11404 6367 11438 6401
rect 11472 6367 11506 6401
rect 11540 6367 11574 6401
rect 11608 6367 11642 6401
rect 11676 6367 11710 6401
rect 11744 6367 11778 6401
rect 11812 6367 11846 6401
rect 11880 6367 11914 6401
rect 11948 6367 11982 6401
rect 12016 6367 12050 6401
rect 12084 6367 12118 6401
rect 12152 6367 12186 6401
rect 12220 6367 12254 6401
rect 12288 6367 12322 6401
rect 12356 6367 12390 6401
rect 12424 6367 12458 6401
rect 12492 6367 12526 6401
rect 12560 6367 12594 6401
rect 12628 6367 12662 6401
rect 12696 6367 12730 6401
rect 12764 6367 12798 6401
rect 12832 6367 12866 6401
rect 12900 6367 12934 6401
rect 12968 6367 13002 6401
rect 13036 6367 13070 6401
rect 13104 6367 13138 6401
rect 13172 6367 13206 6401
rect 13240 6367 13274 6401
rect 13308 6367 13342 6401
rect 688 5432 9494 5534
rect 9534 5500 9636 5568
rect 9528 5432 9562 5466
rect 11468 5503 11502 5537
rect 11536 5503 11570 5537
rect 11604 5503 11638 5537
rect 11672 5503 11706 5537
rect 11740 5503 11774 5537
rect 11808 5503 11842 5537
rect 11876 5503 11910 5537
rect 11944 5503 11978 5537
rect 12012 5503 12046 5537
rect 12080 5503 12114 5537
rect 12148 5503 12182 5537
rect 12216 5503 12250 5537
rect 12284 5503 12318 5537
rect 12352 5503 12386 5537
rect 12420 5503 12454 5537
rect 12488 5503 12522 5537
rect 11370 5415 11404 5449
rect 11370 5347 11404 5381
rect 11370 5279 11404 5313
rect 11370 5211 11404 5245
rect 11370 5143 11404 5177
rect 11370 5075 11404 5109
rect 11370 5007 11404 5041
rect 11370 4939 11404 4973
rect 11370 4871 11404 4905
rect 11370 4803 11404 4837
rect 11370 4735 11404 4769
rect 11370 4667 11404 4701
rect 11370 4599 11404 4633
rect 11370 4531 11404 4565
rect 11370 4463 11404 4497
rect 11370 4395 11404 4429
rect 12522 5415 12556 5449
rect 12522 5347 12556 5381
rect 12522 5279 12556 5313
rect 12522 5211 12556 5245
rect 12522 5143 12556 5177
rect 12522 5075 12556 5109
rect 12522 5007 12556 5041
rect 12522 4939 12556 4973
rect 12522 4871 12556 4905
rect 12522 4803 12556 4837
rect 12522 4735 12556 4769
rect 12522 4667 12556 4701
rect 12522 4599 12556 4633
rect 12522 4531 12556 4565
rect 12522 4463 12556 4497
rect 11370 4327 11404 4361
rect 12522 4395 12556 4429
rect 12522 4327 12556 4361
<< mvnsubdiffcont >>
rect 1949 39899 1983 39933
rect 1834 39797 1936 39865
rect 2017 39831 13951 39933
rect 1834 39729 2004 39797
rect 2085 39763 13883 39831
rect 13985 39778 14019 39812
rect 1834 26979 2072 39729
rect 2153 39695 13815 39763
rect 13917 39676 14019 39744
rect 13849 39608 14019 39676
rect 1834 26911 2004 26979
rect 1834 26843 1936 26911
rect 2038 26840 4044 26908
rect 4078 26874 4112 26908
rect 1834 26775 1868 26809
rect 1970 26806 4044 26840
rect 1970 26772 3976 26806
rect 4096 26772 4198 26840
rect 1902 26738 3976 26772
rect 1902 26670 3908 26738
rect 4028 26704 4198 26772
rect 3960 14634 4198 26704
rect 4028 14566 4198 14634
rect 1920 14528 1954 14562
rect 1988 14494 3994 14562
rect 4096 14498 4198 14566
rect 1834 14426 1936 14494
rect 1988 14460 4062 14494
rect 2056 14426 4062 14460
rect 4164 14430 4198 14464
rect 1834 14358 2004 14426
rect 2056 14392 4130 14426
rect 1834 10856 2072 14358
rect 2124 14324 4130 14392
rect 1834 9012 2072 10746
rect 1834 8944 2004 9012
rect 1834 8876 1936 8944
rect 2038 8872 13700 8940
rect 13781 8906 14019 39608
rect 1834 8808 1868 8842
rect 1970 8804 13768 8872
rect 13849 8838 14019 8906
rect 1902 8702 13836 8804
rect 13917 8770 14019 8838
rect 13870 8702 13904 8736
rect 10604 8423 10638 8457
rect 10672 8423 10706 8457
rect 10740 8423 10774 8457
rect 10808 8423 10842 8457
rect 10876 8423 10910 8457
rect 10944 8423 10978 8457
rect 11012 8423 11046 8457
rect 11080 8423 11114 8457
rect 11148 8423 11182 8457
rect 11216 8423 11250 8457
rect 11284 8423 11318 8457
rect 11352 8423 11386 8457
rect 11420 8423 11454 8457
rect 11488 8423 11522 8457
rect 11556 8423 11590 8457
rect 11624 8423 11658 8457
rect 11692 8423 11726 8457
rect 11760 8423 11794 8457
rect 11828 8423 11862 8457
rect 11896 8423 11930 8457
rect 11964 8423 11998 8457
rect 12032 8423 12066 8457
rect 12100 8423 12134 8457
rect 12168 8423 12202 8457
rect 12236 8423 12270 8457
rect 12304 8423 12338 8457
rect 12372 8423 12406 8457
rect 12440 8423 12474 8457
rect 12508 8423 12542 8457
rect 12576 8423 12610 8457
rect 12644 8423 12678 8457
rect 12712 8423 12746 8457
rect 12780 8423 12814 8457
rect 12848 8423 12882 8457
rect 12916 8423 12950 8457
rect 12984 8423 13018 8457
rect 13052 8423 13086 8457
rect 13120 8423 13154 8457
rect 13188 8423 13222 8457
rect 13256 8423 13290 8457
rect 13324 8423 13358 8457
rect 13392 8423 13426 8457
rect 13460 8423 13494 8457
rect 13528 8423 13562 8457
rect 13596 8423 13630 8457
rect 13664 8423 13698 8457
rect 10473 8355 10507 8389
rect 10473 8287 10507 8321
rect 10605 8291 10639 8325
rect 10676 8291 10710 8325
rect 10744 8291 10778 8325
rect 10812 8291 10846 8325
rect 10880 8291 10914 8325
rect 10948 8291 10982 8325
rect 11016 8291 11050 8325
rect 11084 8291 11118 8325
rect 11152 8291 11186 8325
rect 11220 8291 11254 8325
rect 11288 8291 11322 8325
rect 11356 8291 11390 8325
rect 11424 8291 11458 8325
rect 11492 8291 11526 8325
rect 11560 8291 11594 8325
rect 11628 8291 11662 8325
rect 11696 8291 11730 8325
rect 11764 8291 11798 8325
rect 11832 8291 11866 8325
rect 11900 8291 11934 8325
rect 11968 8291 12002 8325
rect 12036 8291 12070 8325
rect 12104 8291 12138 8325
rect 12172 8291 12206 8325
rect 12240 8291 12274 8325
rect 12308 8291 12342 8325
rect 12376 8291 12410 8325
rect 12444 8291 12478 8325
rect 12512 8291 12546 8325
rect 12580 8291 12614 8325
rect 12648 8291 12682 8325
rect 12716 8291 12750 8325
rect 12784 8291 12818 8325
rect 12852 8291 12886 8325
rect 12920 8291 12954 8325
rect 12988 8291 13022 8325
rect 13056 8291 13090 8325
rect 13124 8291 13158 8325
rect 13192 8291 13226 8325
rect 13260 8291 13294 8325
rect 13328 8291 13362 8325
rect 13396 8291 13430 8325
rect 13464 8291 13498 8325
rect 13532 8291 13566 8325
rect 13600 8291 13634 8325
rect 10473 8219 10507 8253
rect 10605 8223 10639 8257
rect 10473 8151 10507 8185
rect 10605 8155 10639 8189
rect 10473 8083 10507 8117
rect 10605 8087 10639 8121
rect 13732 8290 13766 8324
rect 13600 8218 13634 8252
rect 13732 8222 13766 8256
rect 13600 8150 13634 8184
rect 13732 8154 13766 8188
rect 10473 8015 10507 8049
rect 10605 8019 10639 8053
rect 10473 7947 10507 7981
rect 10605 7951 10639 7985
rect 1059 7485 1093 7519
rect 1127 7485 1161 7519
rect 1195 7485 1229 7519
rect 1263 7485 1297 7519
rect 1331 7485 1365 7519
rect 1399 7485 1433 7519
rect 1467 7485 1501 7519
rect 1535 7485 1569 7519
rect 1603 7485 1637 7519
rect 1671 7485 1705 7519
rect 1739 7485 1773 7519
rect 1807 7485 1841 7519
rect 1875 7485 1909 7519
rect 1943 7485 1977 7519
rect 2011 7485 2045 7519
rect 2079 7485 2113 7519
rect 2147 7485 2181 7519
rect 2215 7485 2249 7519
rect 2283 7485 2317 7519
rect 2351 7485 2385 7519
rect 2419 7485 2453 7519
rect 2487 7485 2521 7519
rect 2555 7485 2589 7519
rect 2623 7485 2657 7519
rect 2691 7485 2725 7519
rect 2759 7485 2793 7519
rect 2827 7485 2861 7519
rect 2895 7485 2929 7519
rect 2963 7485 2997 7519
rect 3031 7485 3065 7519
rect 3099 7485 3133 7519
rect 3167 7485 3201 7519
rect 3235 7485 3269 7519
rect 3303 7485 3337 7519
rect 3371 7485 3405 7519
rect 3439 7485 3473 7519
rect 3507 7485 3541 7519
rect 3575 7485 3609 7519
rect 3643 7485 3677 7519
rect 3711 7485 3745 7519
rect 3779 7485 3813 7519
rect 3847 7485 3881 7519
rect 3915 7485 3949 7519
rect 3983 7485 4017 7519
rect 4051 7485 4085 7519
rect 4119 7485 4153 7519
rect 4187 7485 4221 7519
rect 4255 7485 4289 7519
rect 4323 7485 4357 7519
rect 4391 7485 4425 7519
rect 4459 7485 4493 7519
rect 4527 7485 4561 7519
rect 4595 7485 4629 7519
rect 4663 7485 4697 7519
rect 4731 7485 4765 7519
rect 4799 7485 4833 7519
rect 4867 7485 4901 7519
rect 4935 7485 4969 7519
rect 5003 7485 5037 7519
rect 5071 7485 5105 7519
rect 5139 7485 5173 7519
rect 5207 7485 5241 7519
rect 5275 7485 5309 7519
rect 5343 7485 5377 7519
rect 5411 7485 5445 7519
rect 5479 7485 5513 7519
rect 5547 7485 5581 7519
rect 5615 7485 5649 7519
rect 5683 7485 5717 7519
rect 5751 7485 5785 7519
rect 5819 7485 5853 7519
rect 5887 7485 5921 7519
rect 5955 7485 5989 7519
rect 6023 7485 6057 7519
rect 6091 7485 6125 7519
rect 6159 7485 6193 7519
rect 6227 7485 6261 7519
rect 6295 7485 6329 7519
rect 6363 7485 6397 7519
rect 6431 7485 6465 7519
rect 6499 7485 6533 7519
rect 6567 7485 6601 7519
rect 6635 7485 6669 7519
rect 6703 7485 6737 7519
rect 6771 7485 6805 7519
rect 6839 7485 6873 7519
rect 6907 7485 6941 7519
rect 6975 7485 7009 7519
rect 7043 7485 7077 7519
rect 7111 7485 7145 7519
rect 7179 7485 7213 7519
rect 7247 7485 7281 7519
rect 7315 7485 7349 7519
rect 7383 7485 7417 7519
rect 7451 7485 7485 7519
rect 7519 7485 7553 7519
rect 7587 7485 7621 7519
rect 7655 7485 7689 7519
rect 7723 7485 7757 7519
rect 7791 7485 7825 7519
rect 7859 7485 7893 7519
rect 7927 7485 7961 7519
rect 7995 7485 8029 7519
rect 8063 7485 8097 7519
rect 8131 7485 8165 7519
rect 8199 7485 8233 7519
rect 8267 7485 8301 7519
rect 8335 7485 8369 7519
rect 8403 7485 8437 7519
rect 8471 7485 8505 7519
rect 8539 7485 8573 7519
rect 8607 7485 8641 7519
rect 8675 7485 8709 7519
rect 8743 7485 8777 7519
rect 8811 7485 8845 7519
rect 8879 7485 8913 7519
rect 8947 7485 8981 7519
rect 9015 7485 9049 7519
rect 9083 7485 9117 7519
rect 947 7417 981 7451
rect 9151 7416 9185 7450
rect 947 7349 981 7383
rect 947 7281 981 7315
rect 947 7213 981 7247
rect 947 7145 981 7179
rect 947 7077 981 7111
rect 947 7009 981 7043
rect 947 6941 981 6975
rect 947 6873 981 6907
rect 947 6805 981 6839
rect 947 6737 981 6771
rect 947 6669 981 6703
rect 947 6601 981 6635
rect 947 6533 981 6567
rect 947 6465 981 6499
rect 947 6397 981 6431
rect 947 6329 981 6363
rect 947 6261 981 6295
rect 947 6193 981 6227
rect 947 6125 981 6159
rect 947 6057 981 6091
rect 947 5989 981 6023
rect 9151 7348 9185 7382
rect 9151 7280 9185 7314
rect 9151 7212 9185 7246
rect 9151 7144 9185 7178
rect 9151 7076 9185 7110
rect 9151 7008 9185 7042
rect 9151 6940 9185 6974
rect 9151 6872 9185 6906
rect 9151 6804 9185 6838
rect 9151 6736 9185 6770
rect 9151 6668 9185 6702
rect 9151 6600 9185 6634
rect 9151 6532 9185 6566
rect 9151 6464 9185 6498
rect 9151 6396 9185 6430
rect 9151 6328 9185 6362
rect 9151 6260 9185 6294
rect 9151 6192 9185 6226
rect 9151 6124 9185 6158
rect 9151 6056 9185 6090
rect 9151 5988 9185 6022
rect 9151 5920 9185 5954
rect 1015 5852 1049 5886
rect 1083 5852 1117 5886
rect 1151 5852 1185 5886
rect 1219 5852 1253 5886
rect 1287 5852 1321 5886
rect 1355 5852 1389 5886
rect 1423 5852 1457 5886
rect 1491 5852 1525 5886
rect 1559 5852 1593 5886
rect 1627 5852 1661 5886
rect 1695 5852 1729 5886
rect 1763 5852 1797 5886
rect 1831 5852 1865 5886
rect 1899 5852 1933 5886
rect 1967 5852 2001 5886
rect 2035 5852 2069 5886
rect 2103 5852 2137 5886
rect 2171 5852 2205 5886
rect 2239 5852 2273 5886
rect 2307 5852 2341 5886
rect 2375 5852 2409 5886
rect 2443 5852 2477 5886
rect 2511 5852 2545 5886
rect 2579 5852 2613 5886
rect 2647 5852 2681 5886
rect 2715 5852 2749 5886
rect 2783 5852 2817 5886
rect 2851 5852 2885 5886
rect 2919 5852 2953 5886
rect 2987 5852 3021 5886
rect 3055 5852 3089 5886
rect 3123 5852 3157 5886
rect 3191 5852 3225 5886
rect 3259 5852 3293 5886
rect 3327 5852 3361 5886
rect 3395 5852 3429 5886
rect 3463 5852 3497 5886
rect 3531 5852 3565 5886
rect 3599 5852 3633 5886
rect 3667 5852 3701 5886
rect 3735 5852 3769 5886
rect 3803 5852 3837 5886
rect 3871 5852 3905 5886
rect 3939 5852 3973 5886
rect 4007 5852 4041 5886
rect 4075 5852 4109 5886
rect 4143 5852 4177 5886
rect 4211 5852 4245 5886
rect 4279 5852 4313 5886
rect 4347 5852 4381 5886
rect 4415 5852 4449 5886
rect 4483 5852 4517 5886
rect 4551 5852 4585 5886
rect 4619 5852 4653 5886
rect 4687 5852 4721 5886
rect 4755 5852 4789 5886
rect 4823 5852 4857 5886
rect 4891 5852 4925 5886
rect 4959 5852 4993 5886
rect 5027 5852 5061 5886
rect 5095 5852 5129 5886
rect 5163 5852 5197 5886
rect 5231 5852 5265 5886
rect 5299 5852 5333 5886
rect 5367 5852 5401 5886
rect 5435 5852 5469 5886
rect 5503 5852 5537 5886
rect 5571 5852 5605 5886
rect 5639 5852 5673 5886
rect 5707 5852 5741 5886
rect 5775 5852 5809 5886
rect 5843 5852 5877 5886
rect 5911 5852 5945 5886
rect 5979 5852 6013 5886
rect 6047 5852 6081 5886
rect 6115 5852 6149 5886
rect 6183 5852 6217 5886
rect 6251 5852 6285 5886
rect 6319 5852 6353 5886
rect 6387 5852 6421 5886
rect 6455 5852 6489 5886
rect 6523 5852 6557 5886
rect 6591 5852 6625 5886
rect 6659 5852 6693 5886
rect 6727 5852 6761 5886
rect 6795 5852 6829 5886
rect 6863 5852 6897 5886
rect 6931 5852 6965 5886
rect 6999 5852 7033 5886
rect 7067 5852 7101 5886
rect 7135 5852 7169 5886
rect 7203 5852 7237 5886
rect 7271 5852 7305 5886
rect 7339 5852 7373 5886
rect 7407 5852 7441 5886
rect 7475 5852 7509 5886
rect 7543 5852 7577 5886
rect 7611 5852 7645 5886
rect 7679 5852 7713 5886
rect 7747 5852 7781 5886
rect 7815 5852 7849 5886
rect 7883 5852 7917 5886
rect 7951 5852 7985 5886
rect 8019 5852 8053 5886
rect 8087 5852 8121 5886
rect 8155 5852 8189 5886
rect 8223 5852 8257 5886
rect 8291 5852 8325 5886
rect 8359 5852 8393 5886
rect 8427 5852 8461 5886
rect 8495 5852 8529 5886
rect 8563 5852 8597 5886
rect 8631 5852 8665 5886
rect 8699 5852 8733 5886
rect 8767 5852 8801 5886
rect 8835 5852 8869 5886
rect 8903 5852 8937 5886
rect 8971 5852 9005 5886
rect 9039 5852 9073 5886
rect 10473 7879 10507 7913
rect 10605 7883 10639 7917
rect 10473 7811 10507 7845
rect 10605 7815 10639 7849
rect 10473 7743 10507 7777
rect 10605 7747 10639 7781
rect 10473 7675 10507 7709
rect 10605 7679 10639 7713
rect 10473 7607 10507 7641
rect 10605 7611 10639 7645
rect 10473 7539 10507 7573
rect 10605 7543 10639 7577
rect 10473 7471 10507 7505
rect 10605 7475 10639 7509
rect 10473 7403 10507 7437
rect 10605 7407 10639 7441
rect 10473 7335 10507 7369
rect 10605 7339 10639 7373
rect 10473 7267 10507 7301
rect 10605 7271 10639 7305
rect 10473 7199 10507 7233
rect 10605 7203 10639 7237
rect 10473 7131 10507 7165
rect 10605 7135 10639 7169
rect 10473 7063 10507 7097
rect 10605 7067 10639 7101
rect 10473 6995 10507 7029
rect 10605 6999 10639 7033
rect 10473 6927 10507 6961
rect 10605 6931 10639 6965
rect 10473 6859 10507 6893
rect 10605 6863 10639 6897
rect 10473 6791 10507 6825
rect 10605 6795 10639 6829
rect 10473 6723 10507 6757
rect 10605 6727 10639 6761
rect 10473 6655 10507 6689
rect 10605 6659 10639 6693
rect 10473 6587 10507 6621
rect 10605 6591 10639 6625
rect 10473 6519 10507 6553
rect 10605 6523 10639 6557
rect 10473 6451 10507 6485
rect 10605 6455 10639 6489
rect 13600 8082 13634 8116
rect 13732 8086 13766 8120
rect 13600 8014 13634 8048
rect 13732 8018 13766 8052
rect 13600 7946 13634 7980
rect 13732 7950 13766 7984
rect 13600 7878 13634 7912
rect 13732 7882 13766 7916
rect 13600 7810 13634 7844
rect 13732 7814 13766 7848
rect 13600 7742 13634 7776
rect 13732 7746 13766 7780
rect 13600 7674 13634 7708
rect 13732 7678 13766 7712
rect 13600 7606 13634 7640
rect 13732 7610 13766 7644
rect 13600 7538 13634 7572
rect 13732 7542 13766 7576
rect 13600 7470 13634 7504
rect 13732 7474 13766 7508
rect 13600 7402 13634 7436
rect 13732 7406 13766 7440
rect 13600 7334 13634 7368
rect 13732 7338 13766 7372
rect 13600 7266 13634 7300
rect 13732 7270 13766 7304
rect 13600 7198 13634 7232
rect 13732 7202 13766 7236
rect 13600 7130 13634 7164
rect 13732 7134 13766 7168
rect 13600 7062 13634 7096
rect 13732 7066 13766 7100
rect 13600 6994 13634 7028
rect 13732 6998 13766 7032
rect 13600 6926 13634 6960
rect 13732 6930 13766 6964
rect 13600 6858 13634 6892
rect 13732 6862 13766 6896
rect 13600 6790 13634 6824
rect 13732 6794 13766 6828
rect 13600 6722 13634 6756
rect 13732 6726 13766 6760
rect 13600 6654 13634 6688
rect 13732 6658 13766 6692
rect 13600 6586 13634 6620
rect 13732 6590 13766 6624
rect 13600 6518 13634 6552
rect 13732 6522 13766 6556
rect 13600 6450 13634 6484
rect 13732 6454 13766 6488
rect 13600 6382 13634 6416
rect 13732 6386 13766 6420
rect 10473 6295 10507 6329
rect 10605 6295 10639 6329
rect 10473 6227 10507 6261
rect 13600 6314 13634 6348
rect 13732 6318 13766 6352
rect 13600 6246 13634 6280
rect 13732 6250 13766 6284
rect 10473 6159 10507 6193
rect 10605 6178 10639 6212
rect 10673 6178 10707 6212
rect 10741 6178 10775 6212
rect 10809 6178 10843 6212
rect 10877 6178 10911 6212
rect 10945 6178 10979 6212
rect 11013 6178 11047 6212
rect 11081 6178 11115 6212
rect 11149 6178 11183 6212
rect 11217 6178 11251 6212
rect 11285 6178 11319 6212
rect 11353 6178 11387 6212
rect 11421 6178 11455 6212
rect 11489 6178 11523 6212
rect 11557 6178 11591 6212
rect 11625 6178 11659 6212
rect 11693 6178 11727 6212
rect 11761 6178 11795 6212
rect 11829 6178 11863 6212
rect 11897 6178 11931 6212
rect 11965 6178 11999 6212
rect 12033 6178 12067 6212
rect 12101 6178 12135 6212
rect 12169 6178 12203 6212
rect 12237 6178 12271 6212
rect 12305 6178 12339 6212
rect 12373 6178 12407 6212
rect 12441 6178 12475 6212
rect 12509 6178 12543 6212
rect 12577 6178 12611 6212
rect 12645 6178 12679 6212
rect 12713 6178 12747 6212
rect 12781 6178 12815 6212
rect 12849 6178 12883 6212
rect 12917 6178 12951 6212
rect 12985 6178 13019 6212
rect 13053 6178 13087 6212
rect 13121 6178 13155 6212
rect 13189 6178 13223 6212
rect 13257 6178 13291 6212
rect 13325 6178 13359 6212
rect 13393 6178 13427 6212
rect 13461 6178 13495 6212
rect 13529 6178 13563 6212
rect 13600 6178 13634 6212
rect 13732 6182 13766 6216
rect 13732 6114 13766 6148
rect 10541 6046 10575 6080
rect 10609 6046 10643 6080
rect 10677 6046 10711 6080
rect 10745 6046 10779 6080
rect 10813 6046 10847 6080
rect 10881 6046 10915 6080
rect 10949 6046 10983 6080
rect 11017 6046 11051 6080
rect 11085 6046 11119 6080
rect 11153 6046 11187 6080
rect 11221 6046 11255 6080
rect 11289 6046 11323 6080
rect 11357 6046 11391 6080
rect 11425 6046 11459 6080
rect 11493 6046 11527 6080
rect 11561 6046 11595 6080
rect 11629 6046 11663 6080
rect 11697 6046 11731 6080
rect 11765 6046 11799 6080
rect 11833 6046 11867 6080
rect 11901 6046 11935 6080
rect 11969 6046 12003 6080
rect 12037 6046 12071 6080
rect 12105 6046 12139 6080
rect 12173 6046 12207 6080
rect 12241 6046 12275 6080
rect 12309 6046 12343 6080
rect 12377 6046 12411 6080
rect 12445 6046 12479 6080
rect 12513 6046 12547 6080
rect 12581 6046 12615 6080
rect 12649 6046 12683 6080
rect 12717 6046 12751 6080
rect 12785 6046 12819 6080
rect 12853 6046 12887 6080
rect 12921 6046 12955 6080
rect 12989 6046 13023 6080
rect 13057 6046 13091 6080
rect 13125 6046 13159 6080
rect 13193 6046 13227 6080
rect 13261 6046 13295 6080
rect 13329 6046 13363 6080
rect 13397 6046 13431 6080
rect 13465 6046 13499 6080
rect 13533 6046 13567 6080
rect 13601 6046 13635 6080
rect 10964 5826 10998 5860
rect 10836 5724 10938 5792
rect 11032 5758 14058 5860
rect 10836 4670 11006 5724
rect 11100 5690 13990 5758
rect 14092 5712 14126 5746
rect 14024 5610 14126 5678
rect 2404 4582 2438 4616
rect 2472 4548 10870 4616
rect 10904 4602 11006 4670
rect 2334 4480 2436 4548
rect 2472 4514 10938 4548
rect 10972 4534 11006 4568
rect 2334 502 2504 4480
rect 2540 4446 10938 4514
rect 2334 356 2368 390
rect 2402 356 2436 390
rect 2334 288 2368 322
rect 2470 306 13860 374
rect 13956 340 14126 5610
rect 2402 204 13928 306
rect 14024 272 14126 340
rect 13962 204 13996 238
<< poly >>
rect 3156 39108 3298 39124
rect 3156 39074 3176 39108
rect 3210 39074 3244 39108
rect 3278 39074 3298 39108
rect 3156 39058 3298 39074
rect 3558 39108 3700 39124
rect 3558 39074 3578 39108
rect 3612 39074 3646 39108
rect 3680 39074 3700 39108
rect 3558 39058 3700 39074
rect 4076 39108 4218 39124
rect 4076 39074 4096 39108
rect 4130 39074 4164 39108
rect 4198 39074 4218 39108
rect 4076 39058 4218 39074
rect 4478 39108 4620 39124
rect 4478 39074 4498 39108
rect 4532 39074 4566 39108
rect 4600 39074 4620 39108
rect 4478 39058 4620 39074
rect 4996 39108 5138 39124
rect 4996 39074 5016 39108
rect 5050 39074 5084 39108
rect 5118 39074 5138 39108
rect 4996 39058 5138 39074
rect 5398 39108 5540 39124
rect 5398 39074 5418 39108
rect 5452 39074 5486 39108
rect 5520 39074 5540 39108
rect 5398 39058 5540 39074
rect 5916 39108 6058 39124
rect 5916 39074 5936 39108
rect 5970 39074 6004 39108
rect 6038 39074 6058 39108
rect 5916 39058 6058 39074
rect 6318 39108 6460 39124
rect 6318 39074 6338 39108
rect 6372 39074 6406 39108
rect 6440 39074 6460 39108
rect 6318 39058 6460 39074
rect 6836 39108 6978 39124
rect 6836 39074 6856 39108
rect 6890 39074 6924 39108
rect 6958 39074 6978 39108
rect 6836 39058 6978 39074
rect 7238 39108 7380 39124
rect 7238 39074 7258 39108
rect 7292 39074 7326 39108
rect 7360 39074 7380 39108
rect 7238 39058 7380 39074
rect 7756 39108 7898 39124
rect 7756 39074 7776 39108
rect 7810 39074 7844 39108
rect 7878 39074 7898 39108
rect 7756 39058 7898 39074
rect 8158 39108 8300 39124
rect 8158 39074 8178 39108
rect 8212 39074 8246 39108
rect 8280 39074 8300 39108
rect 8158 39058 8300 39074
rect 8676 39108 8818 39124
rect 8676 39074 8696 39108
rect 8730 39074 8764 39108
rect 8798 39074 8818 39108
rect 8676 39058 8818 39074
rect 9078 39108 9220 39124
rect 9078 39074 9098 39108
rect 9132 39074 9166 39108
rect 9200 39074 9220 39108
rect 9078 39058 9220 39074
rect 9596 39108 9738 39124
rect 9596 39074 9616 39108
rect 9650 39074 9684 39108
rect 9718 39074 9738 39108
rect 9596 39058 9738 39074
rect 9998 39108 10140 39124
rect 9998 39074 10018 39108
rect 10052 39074 10086 39108
rect 10120 39074 10140 39108
rect 9998 39058 10140 39074
rect 10516 39108 10658 39124
rect 10516 39074 10536 39108
rect 10570 39074 10604 39108
rect 10638 39074 10658 39108
rect 10516 39058 10658 39074
rect 10918 39108 11060 39124
rect 10918 39074 10938 39108
rect 10972 39074 11006 39108
rect 11040 39074 11060 39108
rect 10918 39058 11060 39074
rect 11436 39108 11578 39124
rect 11436 39074 11456 39108
rect 11490 39074 11524 39108
rect 11558 39074 11578 39108
rect 11436 39058 11578 39074
rect 11838 39108 11980 39124
rect 11838 39074 11858 39108
rect 11892 39074 11926 39108
rect 11960 39074 11980 39108
rect 11838 39058 11980 39074
rect 12356 39108 12498 39124
rect 12356 39074 12376 39108
rect 12410 39074 12444 39108
rect 12478 39074 12498 39108
rect 12356 39058 12498 39074
rect 12758 39108 12900 39124
rect 12758 39074 12778 39108
rect 12812 39074 12846 39108
rect 12880 39074 12900 39108
rect 12758 39058 12900 39074
rect 3156 36998 3298 37014
rect 3156 36964 3176 36998
rect 3210 36964 3244 36998
rect 3278 36964 3298 36998
rect 3156 36948 3298 36964
rect 3558 36998 3700 37014
rect 3558 36964 3578 36998
rect 3612 36964 3646 36998
rect 3680 36964 3700 36998
rect 3558 36948 3700 36964
rect 4076 36998 4218 37014
rect 4076 36964 4096 36998
rect 4130 36964 4164 36998
rect 4198 36964 4218 36998
rect 4076 36948 4218 36964
rect 4478 36998 4620 37014
rect 4478 36964 4498 36998
rect 4532 36964 4566 36998
rect 4600 36964 4620 36998
rect 4478 36948 4620 36964
rect 4996 36998 5138 37014
rect 4996 36964 5016 36998
rect 5050 36964 5084 36998
rect 5118 36964 5138 36998
rect 4996 36948 5138 36964
rect 5398 36998 5540 37014
rect 5398 36964 5418 36998
rect 5452 36964 5486 36998
rect 5520 36964 5540 36998
rect 5398 36948 5540 36964
rect 5916 36998 6058 37014
rect 5916 36964 5936 36998
rect 5970 36964 6004 36998
rect 6038 36964 6058 36998
rect 5916 36948 6058 36964
rect 6318 36998 6460 37014
rect 6318 36964 6338 36998
rect 6372 36964 6406 36998
rect 6440 36964 6460 36998
rect 6318 36948 6460 36964
rect 6836 36998 6978 37014
rect 6836 36964 6856 36998
rect 6890 36964 6924 36998
rect 6958 36964 6978 36998
rect 6836 36948 6978 36964
rect 7238 36998 7380 37014
rect 7238 36964 7258 36998
rect 7292 36964 7326 36998
rect 7360 36964 7380 36998
rect 7238 36948 7380 36964
rect 7756 36998 7898 37014
rect 7756 36964 7776 36998
rect 7810 36964 7844 36998
rect 7878 36964 7898 36998
rect 7756 36948 7898 36964
rect 8158 36998 8300 37014
rect 8158 36964 8178 36998
rect 8212 36964 8246 36998
rect 8280 36964 8300 36998
rect 8158 36948 8300 36964
rect 8676 36998 8818 37014
rect 8676 36964 8696 36998
rect 8730 36964 8764 36998
rect 8798 36964 8818 36998
rect 8676 36948 8818 36964
rect 9078 36998 9220 37014
rect 9078 36964 9098 36998
rect 9132 36964 9166 36998
rect 9200 36964 9220 36998
rect 9078 36948 9220 36964
rect 9596 36998 9738 37014
rect 9596 36964 9616 36998
rect 9650 36964 9684 36998
rect 9718 36964 9738 36998
rect 9596 36948 9738 36964
rect 9998 36998 10140 37014
rect 9998 36964 10018 36998
rect 10052 36964 10086 36998
rect 10120 36964 10140 36998
rect 9998 36948 10140 36964
rect 10516 36998 10658 37014
rect 10516 36964 10536 36998
rect 10570 36964 10604 36998
rect 10638 36964 10658 36998
rect 10516 36948 10658 36964
rect 10918 36998 11060 37014
rect 10918 36964 10938 36998
rect 10972 36964 11006 36998
rect 11040 36964 11060 36998
rect 10918 36948 11060 36964
rect 11436 36998 11578 37014
rect 11436 36964 11456 36998
rect 11490 36964 11524 36998
rect 11558 36964 11578 36998
rect 11436 36948 11578 36964
rect 11838 36998 11980 37014
rect 11838 36964 11858 36998
rect 11892 36964 11926 36998
rect 11960 36964 11980 36998
rect 11838 36948 11980 36964
rect 12356 36998 12498 37014
rect 12356 36964 12376 36998
rect 12410 36964 12444 36998
rect 12478 36964 12498 36998
rect 12356 36948 12498 36964
rect 12758 36998 12900 37014
rect 12758 36964 12778 36998
rect 12812 36964 12846 36998
rect 12880 36964 12900 36998
rect 12758 36948 12900 36964
rect 3156 36508 3298 36524
rect 3156 36474 3176 36508
rect 3210 36474 3244 36508
rect 3278 36474 3298 36508
rect 3156 36458 3298 36474
rect 3558 36508 3700 36524
rect 3558 36474 3578 36508
rect 3612 36474 3646 36508
rect 3680 36474 3700 36508
rect 3558 36458 3700 36474
rect 4076 36508 4218 36524
rect 4076 36474 4096 36508
rect 4130 36474 4164 36508
rect 4198 36474 4218 36508
rect 4076 36458 4218 36474
rect 4478 36508 4620 36524
rect 4478 36474 4498 36508
rect 4532 36474 4566 36508
rect 4600 36474 4620 36508
rect 4478 36458 4620 36474
rect 4996 36508 5138 36524
rect 4996 36474 5016 36508
rect 5050 36474 5084 36508
rect 5118 36474 5138 36508
rect 4996 36458 5138 36474
rect 5398 36508 5540 36524
rect 5398 36474 5418 36508
rect 5452 36474 5486 36508
rect 5520 36474 5540 36508
rect 5398 36458 5540 36474
rect 5916 36508 6058 36524
rect 5916 36474 5936 36508
rect 5970 36474 6004 36508
rect 6038 36474 6058 36508
rect 5916 36458 6058 36474
rect 6318 36508 6460 36524
rect 6318 36474 6338 36508
rect 6372 36474 6406 36508
rect 6440 36474 6460 36508
rect 6318 36458 6460 36474
rect 6836 36508 6978 36524
rect 6836 36474 6856 36508
rect 6890 36474 6924 36508
rect 6958 36474 6978 36508
rect 6836 36458 6978 36474
rect 7238 36508 7380 36524
rect 7238 36474 7258 36508
rect 7292 36474 7326 36508
rect 7360 36474 7380 36508
rect 7238 36458 7380 36474
rect 7756 36508 7898 36524
rect 7756 36474 7776 36508
rect 7810 36474 7844 36508
rect 7878 36474 7898 36508
rect 7756 36458 7898 36474
rect 8158 36508 8300 36524
rect 8158 36474 8178 36508
rect 8212 36474 8246 36508
rect 8280 36474 8300 36508
rect 8158 36458 8300 36474
rect 8676 36508 8818 36524
rect 8676 36474 8696 36508
rect 8730 36474 8764 36508
rect 8798 36474 8818 36508
rect 8676 36458 8818 36474
rect 9078 36508 9220 36524
rect 9078 36474 9098 36508
rect 9132 36474 9166 36508
rect 9200 36474 9220 36508
rect 9078 36458 9220 36474
rect 9596 36508 9738 36524
rect 9596 36474 9616 36508
rect 9650 36474 9684 36508
rect 9718 36474 9738 36508
rect 9596 36458 9738 36474
rect 9998 36508 10140 36524
rect 9998 36474 10018 36508
rect 10052 36474 10086 36508
rect 10120 36474 10140 36508
rect 9998 36458 10140 36474
rect 10516 36508 10658 36524
rect 10516 36474 10536 36508
rect 10570 36474 10604 36508
rect 10638 36474 10658 36508
rect 10516 36458 10658 36474
rect 10918 36508 11060 36524
rect 10918 36474 10938 36508
rect 10972 36474 11006 36508
rect 11040 36474 11060 36508
rect 10918 36458 11060 36474
rect 11436 36508 11578 36524
rect 11436 36474 11456 36508
rect 11490 36474 11524 36508
rect 11558 36474 11578 36508
rect 11436 36458 11578 36474
rect 11838 36508 11980 36524
rect 11838 36474 11858 36508
rect 11892 36474 11926 36508
rect 11960 36474 11980 36508
rect 11838 36458 11980 36474
rect 12356 36508 12498 36524
rect 12356 36474 12376 36508
rect 12410 36474 12444 36508
rect 12478 36474 12498 36508
rect 12356 36458 12498 36474
rect 12758 36508 12900 36524
rect 12758 36474 12778 36508
rect 12812 36474 12846 36508
rect 12880 36474 12900 36508
rect 12758 36458 12900 36474
rect 3156 32398 3298 32414
rect 3156 32364 3176 32398
rect 3210 32364 3244 32398
rect 3278 32364 3298 32398
rect 3156 32348 3298 32364
rect 3558 32398 3700 32414
rect 3558 32364 3578 32398
rect 3612 32364 3646 32398
rect 3680 32364 3700 32398
rect 3558 32348 3700 32364
rect 4076 32398 4218 32414
rect 4076 32364 4096 32398
rect 4130 32364 4164 32398
rect 4198 32364 4218 32398
rect 4076 32348 4218 32364
rect 4478 32398 4620 32414
rect 4478 32364 4498 32398
rect 4532 32364 4566 32398
rect 4600 32364 4620 32398
rect 4478 32348 4620 32364
rect 4996 32398 5138 32414
rect 4996 32364 5016 32398
rect 5050 32364 5084 32398
rect 5118 32364 5138 32398
rect 4996 32348 5138 32364
rect 5398 32398 5540 32414
rect 5398 32364 5418 32398
rect 5452 32364 5486 32398
rect 5520 32364 5540 32398
rect 5398 32348 5540 32364
rect 5916 32398 6058 32414
rect 5916 32364 5936 32398
rect 5970 32364 6004 32398
rect 6038 32364 6058 32398
rect 5916 32348 6058 32364
rect 6318 32398 6460 32414
rect 6318 32364 6338 32398
rect 6372 32364 6406 32398
rect 6440 32364 6460 32398
rect 6318 32348 6460 32364
rect 6836 32398 6978 32414
rect 6836 32364 6856 32398
rect 6890 32364 6924 32398
rect 6958 32364 6978 32398
rect 6836 32348 6978 32364
rect 7238 32398 7380 32414
rect 7238 32364 7258 32398
rect 7292 32364 7326 32398
rect 7360 32364 7380 32398
rect 7238 32348 7380 32364
rect 7756 32398 7898 32414
rect 7756 32364 7776 32398
rect 7810 32364 7844 32398
rect 7878 32364 7898 32398
rect 7756 32348 7898 32364
rect 8158 32398 8300 32414
rect 8158 32364 8178 32398
rect 8212 32364 8246 32398
rect 8280 32364 8300 32398
rect 8158 32348 8300 32364
rect 8676 32398 8818 32414
rect 8676 32364 8696 32398
rect 8730 32364 8764 32398
rect 8798 32364 8818 32398
rect 8676 32348 8818 32364
rect 9078 32398 9220 32414
rect 9078 32364 9098 32398
rect 9132 32364 9166 32398
rect 9200 32364 9220 32398
rect 9078 32348 9220 32364
rect 9596 32398 9738 32414
rect 9596 32364 9616 32398
rect 9650 32364 9684 32398
rect 9718 32364 9738 32398
rect 9596 32348 9738 32364
rect 9998 32398 10140 32414
rect 9998 32364 10018 32398
rect 10052 32364 10086 32398
rect 10120 32364 10140 32398
rect 9998 32348 10140 32364
rect 10516 32398 10658 32414
rect 10516 32364 10536 32398
rect 10570 32364 10604 32398
rect 10638 32364 10658 32398
rect 10516 32348 10658 32364
rect 10918 32398 11060 32414
rect 10918 32364 10938 32398
rect 10972 32364 11006 32398
rect 11040 32364 11060 32398
rect 10918 32348 11060 32364
rect 11436 32398 11578 32414
rect 11436 32364 11456 32398
rect 11490 32364 11524 32398
rect 11558 32364 11578 32398
rect 11436 32348 11578 32364
rect 11838 32398 11980 32414
rect 11838 32364 11858 32398
rect 11892 32364 11926 32398
rect 11960 32364 11980 32398
rect 11838 32348 11980 32364
rect 12356 32398 12498 32414
rect 12356 32364 12376 32398
rect 12410 32364 12444 32398
rect 12478 32364 12498 32398
rect 12356 32348 12498 32364
rect 12758 32398 12900 32414
rect 12758 32364 12778 32398
rect 12812 32364 12846 32398
rect 12880 32364 12900 32398
rect 12758 32348 12900 32364
rect 3156 31908 3298 31924
rect 3156 31874 3176 31908
rect 3210 31874 3244 31908
rect 3278 31874 3298 31908
rect 3156 31858 3298 31874
rect 3558 31908 3700 31924
rect 3558 31874 3578 31908
rect 3612 31874 3646 31908
rect 3680 31874 3700 31908
rect 3558 31858 3700 31874
rect 4076 31908 4218 31924
rect 4076 31874 4096 31908
rect 4130 31874 4164 31908
rect 4198 31874 4218 31908
rect 4076 31858 4218 31874
rect 4478 31908 4620 31924
rect 4478 31874 4498 31908
rect 4532 31874 4566 31908
rect 4600 31874 4620 31908
rect 4478 31858 4620 31874
rect 4996 31908 5138 31924
rect 4996 31874 5016 31908
rect 5050 31874 5084 31908
rect 5118 31874 5138 31908
rect 4996 31858 5138 31874
rect 5398 31908 5540 31924
rect 5398 31874 5418 31908
rect 5452 31874 5486 31908
rect 5520 31874 5540 31908
rect 5398 31858 5540 31874
rect 5916 31908 6058 31924
rect 5916 31874 5936 31908
rect 5970 31874 6004 31908
rect 6038 31874 6058 31908
rect 5916 31858 6058 31874
rect 6318 31908 6460 31924
rect 6318 31874 6338 31908
rect 6372 31874 6406 31908
rect 6440 31874 6460 31908
rect 6318 31858 6460 31874
rect 6836 31908 6978 31924
rect 6836 31874 6856 31908
rect 6890 31874 6924 31908
rect 6958 31874 6978 31908
rect 6836 31858 6978 31874
rect 7238 31908 7380 31924
rect 7238 31874 7258 31908
rect 7292 31874 7326 31908
rect 7360 31874 7380 31908
rect 7238 31858 7380 31874
rect 7756 31908 7898 31924
rect 7756 31874 7776 31908
rect 7810 31874 7844 31908
rect 7878 31874 7898 31908
rect 7756 31858 7898 31874
rect 8158 31908 8300 31924
rect 8158 31874 8178 31908
rect 8212 31874 8246 31908
rect 8280 31874 8300 31908
rect 8158 31858 8300 31874
rect 8676 31908 8818 31924
rect 8676 31874 8696 31908
rect 8730 31874 8764 31908
rect 8798 31874 8818 31908
rect 8676 31858 8818 31874
rect 9078 31908 9220 31924
rect 9078 31874 9098 31908
rect 9132 31874 9166 31908
rect 9200 31874 9220 31908
rect 9078 31858 9220 31874
rect 9596 31908 9738 31924
rect 9596 31874 9616 31908
rect 9650 31874 9684 31908
rect 9718 31874 9738 31908
rect 9596 31858 9738 31874
rect 9998 31908 10140 31924
rect 9998 31874 10018 31908
rect 10052 31874 10086 31908
rect 10120 31874 10140 31908
rect 9998 31858 10140 31874
rect 10516 31908 10658 31924
rect 10516 31874 10536 31908
rect 10570 31874 10604 31908
rect 10638 31874 10658 31908
rect 10516 31858 10658 31874
rect 10918 31908 11060 31924
rect 10918 31874 10938 31908
rect 10972 31874 11006 31908
rect 11040 31874 11060 31908
rect 10918 31858 11060 31874
rect 11436 31908 11578 31924
rect 11436 31874 11456 31908
rect 11490 31874 11524 31908
rect 11558 31874 11578 31908
rect 11436 31858 11578 31874
rect 11838 31908 11980 31924
rect 11838 31874 11858 31908
rect 11892 31874 11926 31908
rect 11960 31874 11980 31908
rect 11838 31858 11980 31874
rect 12356 31908 12498 31924
rect 12356 31874 12376 31908
rect 12410 31874 12444 31908
rect 12478 31874 12498 31908
rect 12356 31858 12498 31874
rect 12758 31908 12900 31924
rect 12758 31874 12778 31908
rect 12812 31874 12846 31908
rect 12880 31874 12900 31908
rect 12758 31858 12900 31874
rect 3156 27798 3298 27814
rect 3156 27764 3176 27798
rect 3210 27764 3244 27798
rect 3278 27764 3298 27798
rect 3156 27748 3298 27764
rect 3558 27798 3700 27814
rect 3558 27764 3578 27798
rect 3612 27764 3646 27798
rect 3680 27764 3700 27798
rect 3558 27748 3700 27764
rect 4076 27798 4218 27814
rect 4076 27764 4096 27798
rect 4130 27764 4164 27798
rect 4198 27764 4218 27798
rect 4076 27748 4218 27764
rect 4478 27798 4620 27814
rect 4478 27764 4498 27798
rect 4532 27764 4566 27798
rect 4600 27764 4620 27798
rect 4478 27748 4620 27764
rect 4996 27798 5138 27814
rect 4996 27764 5016 27798
rect 5050 27764 5084 27798
rect 5118 27764 5138 27798
rect 4996 27748 5138 27764
rect 5398 27798 5540 27814
rect 5398 27764 5418 27798
rect 5452 27764 5486 27798
rect 5520 27764 5540 27798
rect 5398 27748 5540 27764
rect 5916 27798 6058 27814
rect 5916 27764 5936 27798
rect 5970 27764 6004 27798
rect 6038 27764 6058 27798
rect 5916 27748 6058 27764
rect 6318 27798 6460 27814
rect 6318 27764 6338 27798
rect 6372 27764 6406 27798
rect 6440 27764 6460 27798
rect 6318 27748 6460 27764
rect 6836 27798 6978 27814
rect 6836 27764 6856 27798
rect 6890 27764 6924 27798
rect 6958 27764 6978 27798
rect 6836 27748 6978 27764
rect 7238 27798 7380 27814
rect 7238 27764 7258 27798
rect 7292 27764 7326 27798
rect 7360 27764 7380 27798
rect 7238 27748 7380 27764
rect 7756 27798 7898 27814
rect 7756 27764 7776 27798
rect 7810 27764 7844 27798
rect 7878 27764 7898 27798
rect 7756 27748 7898 27764
rect 8158 27798 8300 27814
rect 8158 27764 8178 27798
rect 8212 27764 8246 27798
rect 8280 27764 8300 27798
rect 8158 27748 8300 27764
rect 8676 27798 8818 27814
rect 8676 27764 8696 27798
rect 8730 27764 8764 27798
rect 8798 27764 8818 27798
rect 8676 27748 8818 27764
rect 9078 27798 9220 27814
rect 9078 27764 9098 27798
rect 9132 27764 9166 27798
rect 9200 27764 9220 27798
rect 9078 27748 9220 27764
rect 9596 27798 9738 27814
rect 9596 27764 9616 27798
rect 9650 27764 9684 27798
rect 9718 27764 9738 27798
rect 9596 27748 9738 27764
rect 9998 27798 10140 27814
rect 9998 27764 10018 27798
rect 10052 27764 10086 27798
rect 10120 27764 10140 27798
rect 9998 27748 10140 27764
rect 10516 27798 10658 27814
rect 10516 27764 10536 27798
rect 10570 27764 10604 27798
rect 10638 27764 10658 27798
rect 10516 27748 10658 27764
rect 10918 27798 11060 27814
rect 10918 27764 10938 27798
rect 10972 27764 11006 27798
rect 11040 27764 11060 27798
rect 10918 27748 11060 27764
rect 11436 27798 11578 27814
rect 11436 27764 11456 27798
rect 11490 27764 11524 27798
rect 11558 27764 11578 27798
rect 11436 27748 11578 27764
rect 11838 27798 11980 27814
rect 11838 27764 11858 27798
rect 11892 27764 11926 27798
rect 11960 27764 11980 27798
rect 11838 27748 11980 27764
rect 12356 27798 12498 27814
rect 12356 27764 12376 27798
rect 12410 27764 12444 27798
rect 12478 27764 12498 27798
rect 12356 27748 12498 27764
rect 12758 27798 12900 27814
rect 12758 27764 12778 27798
rect 12812 27764 12846 27798
rect 12880 27764 12900 27798
rect 12758 27748 12900 27764
rect 4996 27308 5138 27324
rect 4996 27274 5016 27308
rect 5050 27274 5084 27308
rect 5118 27274 5138 27308
rect 4996 27258 5138 27274
rect 5398 27308 5540 27324
rect 5398 27274 5418 27308
rect 5452 27274 5486 27308
rect 5520 27274 5540 27308
rect 5398 27258 5540 27274
rect 5916 27308 6058 27324
rect 5916 27274 5936 27308
rect 5970 27274 6004 27308
rect 6038 27274 6058 27308
rect 5916 27258 6058 27274
rect 6318 27308 6460 27324
rect 6318 27274 6338 27308
rect 6372 27274 6406 27308
rect 6440 27274 6460 27308
rect 6318 27258 6460 27274
rect 6836 27308 6978 27324
rect 6836 27274 6856 27308
rect 6890 27274 6924 27308
rect 6958 27274 6978 27308
rect 6836 27258 6978 27274
rect 7238 27308 7380 27324
rect 7238 27274 7258 27308
rect 7292 27274 7326 27308
rect 7360 27274 7380 27308
rect 7238 27258 7380 27274
rect 7756 27308 7898 27324
rect 7756 27274 7776 27308
rect 7810 27274 7844 27308
rect 7878 27274 7898 27308
rect 7756 27258 7898 27274
rect 8158 27308 8300 27324
rect 8158 27274 8178 27308
rect 8212 27274 8246 27308
rect 8280 27274 8300 27308
rect 8158 27258 8300 27274
rect 8676 27308 8818 27324
rect 8676 27274 8696 27308
rect 8730 27274 8764 27308
rect 8798 27274 8818 27308
rect 8676 27258 8818 27274
rect 9078 27308 9220 27324
rect 9078 27274 9098 27308
rect 9132 27274 9166 27308
rect 9200 27274 9220 27308
rect 9078 27258 9220 27274
rect 9596 27308 9738 27324
rect 9596 27274 9616 27308
rect 9650 27274 9684 27308
rect 9718 27274 9738 27308
rect 9596 27258 9738 27274
rect 9998 27308 10140 27324
rect 9998 27274 10018 27308
rect 10052 27274 10086 27308
rect 10120 27274 10140 27308
rect 9998 27258 10140 27274
rect 10516 27308 10658 27324
rect 10516 27274 10536 27308
rect 10570 27274 10604 27308
rect 10638 27274 10658 27308
rect 10516 27258 10658 27274
rect 10918 27308 11060 27324
rect 10918 27274 10938 27308
rect 10972 27274 11006 27308
rect 11040 27274 11060 27308
rect 10918 27258 11060 27274
rect 11436 27308 11578 27324
rect 11436 27274 11456 27308
rect 11490 27274 11524 27308
rect 11558 27274 11578 27308
rect 11436 27258 11578 27274
rect 11838 27308 11980 27324
rect 11838 27274 11858 27308
rect 11892 27274 11926 27308
rect 11960 27274 11980 27308
rect 11838 27258 11980 27274
rect 12356 27308 12498 27324
rect 12356 27274 12376 27308
rect 12410 27274 12444 27308
rect 12478 27274 12498 27308
rect 12356 27258 12498 27274
rect 12758 27308 12900 27324
rect 12758 27274 12778 27308
rect 12812 27274 12846 27308
rect 12880 27274 12900 27308
rect 12758 27258 12900 27274
rect 4996 23198 5138 23214
rect 4996 23164 5016 23198
rect 5050 23164 5084 23198
rect 5118 23164 5138 23198
rect 4996 23148 5138 23164
rect 5398 23198 5540 23214
rect 5398 23164 5418 23198
rect 5452 23164 5486 23198
rect 5520 23164 5540 23198
rect 5398 23148 5540 23164
rect 5916 23198 6058 23214
rect 5916 23164 5936 23198
rect 5970 23164 6004 23198
rect 6038 23164 6058 23198
rect 5916 23148 6058 23164
rect 6318 23198 6460 23214
rect 6318 23164 6338 23198
rect 6372 23164 6406 23198
rect 6440 23164 6460 23198
rect 6318 23148 6460 23164
rect 6836 23198 6978 23214
rect 6836 23164 6856 23198
rect 6890 23164 6924 23198
rect 6958 23164 6978 23198
rect 6836 23148 6978 23164
rect 7238 23198 7380 23214
rect 7238 23164 7258 23198
rect 7292 23164 7326 23198
rect 7360 23164 7380 23198
rect 7238 23148 7380 23164
rect 7756 23198 7898 23214
rect 7756 23164 7776 23198
rect 7810 23164 7844 23198
rect 7878 23164 7898 23198
rect 7756 23148 7898 23164
rect 8158 23198 8300 23214
rect 8158 23164 8178 23198
rect 8212 23164 8246 23198
rect 8280 23164 8300 23198
rect 8158 23148 8300 23164
rect 8676 23198 8818 23214
rect 8676 23164 8696 23198
rect 8730 23164 8764 23198
rect 8798 23164 8818 23198
rect 8676 23148 8818 23164
rect 9078 23198 9220 23214
rect 9078 23164 9098 23198
rect 9132 23164 9166 23198
rect 9200 23164 9220 23198
rect 9078 23148 9220 23164
rect 9596 23198 9738 23214
rect 9596 23164 9616 23198
rect 9650 23164 9684 23198
rect 9718 23164 9738 23198
rect 9596 23148 9738 23164
rect 9998 23198 10140 23214
rect 9998 23164 10018 23198
rect 10052 23164 10086 23198
rect 10120 23164 10140 23198
rect 9998 23148 10140 23164
rect 10516 23198 10658 23214
rect 10516 23164 10536 23198
rect 10570 23164 10604 23198
rect 10638 23164 10658 23198
rect 10516 23148 10658 23164
rect 10918 23198 11060 23214
rect 10918 23164 10938 23198
rect 10972 23164 11006 23198
rect 11040 23164 11060 23198
rect 10918 23148 11060 23164
rect 11436 23198 11578 23214
rect 11436 23164 11456 23198
rect 11490 23164 11524 23198
rect 11558 23164 11578 23198
rect 11436 23148 11578 23164
rect 11838 23198 11980 23214
rect 11838 23164 11858 23198
rect 11892 23164 11926 23198
rect 11960 23164 11980 23198
rect 11838 23148 11980 23164
rect 12356 23198 12498 23214
rect 12356 23164 12376 23198
rect 12410 23164 12444 23198
rect 12478 23164 12498 23198
rect 12356 23148 12498 23164
rect 12758 23198 12900 23214
rect 12758 23164 12778 23198
rect 12812 23164 12846 23198
rect 12880 23164 12900 23198
rect 12758 23148 12900 23164
rect 4996 22708 5138 22724
rect 4996 22674 5016 22708
rect 5050 22674 5084 22708
rect 5118 22674 5138 22708
rect 4996 22658 5138 22674
rect 5398 22708 5540 22724
rect 5398 22674 5418 22708
rect 5452 22674 5486 22708
rect 5520 22674 5540 22708
rect 5398 22658 5540 22674
rect 5916 22708 6058 22724
rect 5916 22674 5936 22708
rect 5970 22674 6004 22708
rect 6038 22674 6058 22708
rect 5916 22658 6058 22674
rect 6318 22708 6460 22724
rect 6318 22674 6338 22708
rect 6372 22674 6406 22708
rect 6440 22674 6460 22708
rect 6318 22658 6460 22674
rect 6836 22708 6978 22724
rect 6836 22674 6856 22708
rect 6890 22674 6924 22708
rect 6958 22674 6978 22708
rect 6836 22658 6978 22674
rect 7238 22708 7380 22724
rect 7238 22674 7258 22708
rect 7292 22674 7326 22708
rect 7360 22674 7380 22708
rect 7238 22658 7380 22674
rect 7756 22708 7898 22724
rect 7756 22674 7776 22708
rect 7810 22674 7844 22708
rect 7878 22674 7898 22708
rect 7756 22658 7898 22674
rect 8158 22708 8300 22724
rect 8158 22674 8178 22708
rect 8212 22674 8246 22708
rect 8280 22674 8300 22708
rect 8158 22658 8300 22674
rect 8676 22708 8818 22724
rect 8676 22674 8696 22708
rect 8730 22674 8764 22708
rect 8798 22674 8818 22708
rect 8676 22658 8818 22674
rect 9078 22708 9220 22724
rect 9078 22674 9098 22708
rect 9132 22674 9166 22708
rect 9200 22674 9220 22708
rect 9078 22658 9220 22674
rect 9596 22708 9738 22724
rect 9596 22674 9616 22708
rect 9650 22674 9684 22708
rect 9718 22674 9738 22708
rect 9596 22658 9738 22674
rect 9998 22708 10140 22724
rect 9998 22674 10018 22708
rect 10052 22674 10086 22708
rect 10120 22674 10140 22708
rect 9998 22658 10140 22674
rect 10516 22708 10658 22724
rect 10516 22674 10536 22708
rect 10570 22674 10604 22708
rect 10638 22674 10658 22708
rect 10516 22658 10658 22674
rect 10918 22708 11060 22724
rect 10918 22674 10938 22708
rect 10972 22674 11006 22708
rect 11040 22674 11060 22708
rect 10918 22658 11060 22674
rect 11436 22708 11578 22724
rect 11436 22674 11456 22708
rect 11490 22674 11524 22708
rect 11558 22674 11578 22708
rect 11436 22658 11578 22674
rect 11838 22708 11980 22724
rect 11838 22674 11858 22708
rect 11892 22674 11926 22708
rect 11960 22674 11980 22708
rect 11838 22658 11980 22674
rect 12356 22708 12498 22724
rect 12356 22674 12376 22708
rect 12410 22674 12444 22708
rect 12478 22674 12498 22708
rect 12356 22658 12498 22674
rect 12758 22708 12900 22724
rect 12758 22674 12778 22708
rect 12812 22674 12846 22708
rect 12880 22674 12900 22708
rect 12758 22658 12900 22674
rect 4996 18598 5138 18614
rect 4996 18564 5016 18598
rect 5050 18564 5084 18598
rect 5118 18564 5138 18598
rect 4996 18548 5138 18564
rect 5398 18598 5540 18614
rect 5398 18564 5418 18598
rect 5452 18564 5486 18598
rect 5520 18564 5540 18598
rect 5398 18548 5540 18564
rect 5916 18598 6058 18614
rect 5916 18564 5936 18598
rect 5970 18564 6004 18598
rect 6038 18564 6058 18598
rect 5916 18548 6058 18564
rect 6318 18598 6460 18614
rect 6318 18564 6338 18598
rect 6372 18564 6406 18598
rect 6440 18564 6460 18598
rect 6318 18548 6460 18564
rect 6836 18598 6978 18614
rect 6836 18564 6856 18598
rect 6890 18564 6924 18598
rect 6958 18564 6978 18598
rect 6836 18548 6978 18564
rect 7238 18598 7380 18614
rect 7238 18564 7258 18598
rect 7292 18564 7326 18598
rect 7360 18564 7380 18598
rect 7238 18548 7380 18564
rect 7756 18598 7898 18614
rect 7756 18564 7776 18598
rect 7810 18564 7844 18598
rect 7878 18564 7898 18598
rect 7756 18548 7898 18564
rect 8158 18598 8300 18614
rect 8158 18564 8178 18598
rect 8212 18564 8246 18598
rect 8280 18564 8300 18598
rect 8158 18548 8300 18564
rect 8676 18598 8818 18614
rect 8676 18564 8696 18598
rect 8730 18564 8764 18598
rect 8798 18564 8818 18598
rect 8676 18548 8818 18564
rect 9078 18598 9220 18614
rect 9078 18564 9098 18598
rect 9132 18564 9166 18598
rect 9200 18564 9220 18598
rect 9078 18548 9220 18564
rect 9596 18598 9738 18614
rect 9596 18564 9616 18598
rect 9650 18564 9684 18598
rect 9718 18564 9738 18598
rect 9596 18548 9738 18564
rect 9998 18598 10140 18614
rect 9998 18564 10018 18598
rect 10052 18564 10086 18598
rect 10120 18564 10140 18598
rect 9998 18548 10140 18564
rect 10516 18598 10658 18614
rect 10516 18564 10536 18598
rect 10570 18564 10604 18598
rect 10638 18564 10658 18598
rect 10516 18548 10658 18564
rect 10918 18598 11060 18614
rect 10918 18564 10938 18598
rect 10972 18564 11006 18598
rect 11040 18564 11060 18598
rect 10918 18548 11060 18564
rect 11436 18598 11578 18614
rect 11436 18564 11456 18598
rect 11490 18564 11524 18598
rect 11558 18564 11578 18598
rect 11436 18548 11578 18564
rect 11838 18598 11980 18614
rect 11838 18564 11858 18598
rect 11892 18564 11926 18598
rect 11960 18564 11980 18598
rect 11838 18548 11980 18564
rect 12356 18598 12498 18614
rect 12356 18564 12376 18598
rect 12410 18564 12444 18598
rect 12478 18564 12498 18598
rect 12356 18548 12498 18564
rect 12758 18598 12900 18614
rect 12758 18564 12778 18598
rect 12812 18564 12846 18598
rect 12880 18564 12900 18598
rect 12758 18548 12900 18564
rect 4996 18108 5138 18124
rect 4996 18074 5016 18108
rect 5050 18074 5084 18108
rect 5118 18074 5138 18108
rect 4996 18058 5138 18074
rect 5398 18108 5540 18124
rect 5398 18074 5418 18108
rect 5452 18074 5486 18108
rect 5520 18074 5540 18108
rect 5398 18058 5540 18074
rect 5916 18108 6058 18124
rect 5916 18074 5936 18108
rect 5970 18074 6004 18108
rect 6038 18074 6058 18108
rect 5916 18058 6058 18074
rect 6318 18108 6460 18124
rect 6318 18074 6338 18108
rect 6372 18074 6406 18108
rect 6440 18074 6460 18108
rect 6318 18058 6460 18074
rect 6836 18108 6978 18124
rect 6836 18074 6856 18108
rect 6890 18074 6924 18108
rect 6958 18074 6978 18108
rect 6836 18058 6978 18074
rect 7238 18108 7380 18124
rect 7238 18074 7258 18108
rect 7292 18074 7326 18108
rect 7360 18074 7380 18108
rect 7238 18058 7380 18074
rect 7756 18108 7898 18124
rect 7756 18074 7776 18108
rect 7810 18074 7844 18108
rect 7878 18074 7898 18108
rect 7756 18058 7898 18074
rect 8158 18108 8300 18124
rect 8158 18074 8178 18108
rect 8212 18074 8246 18108
rect 8280 18074 8300 18108
rect 8158 18058 8300 18074
rect 8676 18108 8818 18124
rect 8676 18074 8696 18108
rect 8730 18074 8764 18108
rect 8798 18074 8818 18108
rect 8676 18058 8818 18074
rect 9078 18108 9220 18124
rect 9078 18074 9098 18108
rect 9132 18074 9166 18108
rect 9200 18074 9220 18108
rect 9078 18058 9220 18074
rect 9596 18108 9738 18124
rect 9596 18074 9616 18108
rect 9650 18074 9684 18108
rect 9718 18074 9738 18108
rect 9596 18058 9738 18074
rect 9998 18108 10140 18124
rect 9998 18074 10018 18108
rect 10052 18074 10086 18108
rect 10120 18074 10140 18108
rect 9998 18058 10140 18074
rect 10516 18108 10658 18124
rect 10516 18074 10536 18108
rect 10570 18074 10604 18108
rect 10638 18074 10658 18108
rect 10516 18058 10658 18074
rect 10918 18108 11060 18124
rect 10918 18074 10938 18108
rect 10972 18074 11006 18108
rect 11040 18074 11060 18108
rect 10918 18058 11060 18074
rect 11436 18108 11578 18124
rect 11436 18074 11456 18108
rect 11490 18074 11524 18108
rect 11558 18074 11578 18108
rect 11436 18058 11578 18074
rect 11838 18108 11980 18124
rect 11838 18074 11858 18108
rect 11892 18074 11926 18108
rect 11960 18074 11980 18108
rect 11838 18058 11980 18074
rect 12356 18108 12498 18124
rect 12356 18074 12376 18108
rect 12410 18074 12444 18108
rect 12478 18074 12498 18108
rect 12356 18058 12498 18074
rect 12758 18108 12900 18124
rect 12758 18074 12778 18108
rect 12812 18074 12846 18108
rect 12880 18074 12900 18108
rect 12758 18058 12900 18074
rect 4996 13998 5138 14014
rect 4996 13964 5016 13998
rect 5050 13964 5084 13998
rect 5118 13964 5138 13998
rect 4996 13948 5138 13964
rect 5398 13998 5540 14014
rect 5398 13964 5418 13998
rect 5452 13964 5486 13998
rect 5520 13964 5540 13998
rect 5398 13948 5540 13964
rect 5916 13998 6058 14014
rect 5916 13964 5936 13998
rect 5970 13964 6004 13998
rect 6038 13964 6058 13998
rect 5916 13948 6058 13964
rect 6318 13998 6460 14014
rect 6318 13964 6338 13998
rect 6372 13964 6406 13998
rect 6440 13964 6460 13998
rect 6318 13948 6460 13964
rect 6836 13998 6978 14014
rect 6836 13964 6856 13998
rect 6890 13964 6924 13998
rect 6958 13964 6978 13998
rect 6836 13948 6978 13964
rect 7238 13998 7380 14014
rect 7238 13964 7258 13998
rect 7292 13964 7326 13998
rect 7360 13964 7380 13998
rect 7238 13948 7380 13964
rect 7756 13998 7898 14014
rect 7756 13964 7776 13998
rect 7810 13964 7844 13998
rect 7878 13964 7898 13998
rect 7756 13948 7898 13964
rect 8158 13998 8300 14014
rect 8158 13964 8178 13998
rect 8212 13964 8246 13998
rect 8280 13964 8300 13998
rect 8158 13948 8300 13964
rect 8676 13998 8818 14014
rect 8676 13964 8696 13998
rect 8730 13964 8764 13998
rect 8798 13964 8818 13998
rect 8676 13948 8818 13964
rect 9078 13998 9220 14014
rect 9078 13964 9098 13998
rect 9132 13964 9166 13998
rect 9200 13964 9220 13998
rect 9078 13948 9220 13964
rect 9596 13998 9738 14014
rect 9596 13964 9616 13998
rect 9650 13964 9684 13998
rect 9718 13964 9738 13998
rect 9596 13948 9738 13964
rect 9998 13998 10140 14014
rect 9998 13964 10018 13998
rect 10052 13964 10086 13998
rect 10120 13964 10140 13998
rect 9998 13948 10140 13964
rect 10516 13998 10658 14014
rect 10516 13964 10536 13998
rect 10570 13964 10604 13998
rect 10638 13964 10658 13998
rect 10516 13948 10658 13964
rect 10918 13998 11060 14014
rect 10918 13964 10938 13998
rect 10972 13964 11006 13998
rect 11040 13964 11060 13998
rect 10918 13948 11060 13964
rect 11436 13998 11578 14014
rect 11436 13964 11456 13998
rect 11490 13964 11524 13998
rect 11558 13964 11578 13998
rect 11436 13948 11578 13964
rect 11838 13998 11980 14014
rect 11838 13964 11858 13998
rect 11892 13964 11926 13998
rect 11960 13964 11980 13998
rect 11838 13948 11980 13964
rect 12356 13998 12498 14014
rect 12356 13964 12376 13998
rect 12410 13964 12444 13998
rect 12478 13964 12498 13998
rect 12356 13948 12498 13964
rect 12758 13998 12900 14014
rect 12758 13964 12778 13998
rect 12812 13964 12846 13998
rect 12880 13964 12900 13998
rect 12758 13948 12900 13964
rect 3156 13508 3298 13524
rect 3156 13474 3176 13508
rect 3210 13474 3244 13508
rect 3278 13474 3298 13508
rect 3156 13458 3298 13474
rect 3558 13508 3700 13524
rect 3558 13474 3578 13508
rect 3612 13474 3646 13508
rect 3680 13474 3700 13508
rect 3558 13458 3700 13474
rect 4076 13508 4218 13524
rect 4076 13474 4096 13508
rect 4130 13474 4164 13508
rect 4198 13474 4218 13508
rect 4076 13458 4218 13474
rect 4478 13508 4620 13524
rect 4478 13474 4498 13508
rect 4532 13474 4566 13508
rect 4600 13474 4620 13508
rect 4478 13458 4620 13474
rect 4996 13508 5138 13524
rect 4996 13474 5016 13508
rect 5050 13474 5084 13508
rect 5118 13474 5138 13508
rect 4996 13458 5138 13474
rect 5398 13508 5540 13524
rect 5398 13474 5418 13508
rect 5452 13474 5486 13508
rect 5520 13474 5540 13508
rect 5398 13458 5540 13474
rect 5916 13508 6058 13524
rect 5916 13474 5936 13508
rect 5970 13474 6004 13508
rect 6038 13474 6058 13508
rect 5916 13458 6058 13474
rect 6318 13508 6460 13524
rect 6318 13474 6338 13508
rect 6372 13474 6406 13508
rect 6440 13474 6460 13508
rect 6318 13458 6460 13474
rect 6836 13508 6978 13524
rect 6836 13474 6856 13508
rect 6890 13474 6924 13508
rect 6958 13474 6978 13508
rect 6836 13458 6978 13474
rect 7238 13508 7380 13524
rect 7238 13474 7258 13508
rect 7292 13474 7326 13508
rect 7360 13474 7380 13508
rect 7238 13458 7380 13474
rect 7756 13508 7898 13524
rect 7756 13474 7776 13508
rect 7810 13474 7844 13508
rect 7878 13474 7898 13508
rect 7756 13458 7898 13474
rect 8158 13508 8300 13524
rect 8158 13474 8178 13508
rect 8212 13474 8246 13508
rect 8280 13474 8300 13508
rect 8158 13458 8300 13474
rect 8676 13508 8818 13524
rect 8676 13474 8696 13508
rect 8730 13474 8764 13508
rect 8798 13474 8818 13508
rect 8676 13458 8818 13474
rect 9078 13508 9220 13524
rect 9078 13474 9098 13508
rect 9132 13474 9166 13508
rect 9200 13474 9220 13508
rect 9078 13458 9220 13474
rect 9596 13508 9738 13524
rect 9596 13474 9616 13508
rect 9650 13474 9684 13508
rect 9718 13474 9738 13508
rect 9596 13458 9738 13474
rect 9998 13508 10140 13524
rect 9998 13474 10018 13508
rect 10052 13474 10086 13508
rect 10120 13474 10140 13508
rect 9998 13458 10140 13474
rect 10516 13508 10658 13524
rect 10516 13474 10536 13508
rect 10570 13474 10604 13508
rect 10638 13474 10658 13508
rect 10516 13458 10658 13474
rect 10918 13508 11060 13524
rect 10918 13474 10938 13508
rect 10972 13474 11006 13508
rect 11040 13474 11060 13508
rect 10918 13458 11060 13474
rect 11436 13508 11578 13524
rect 11436 13474 11456 13508
rect 11490 13474 11524 13508
rect 11558 13474 11578 13508
rect 11436 13458 11578 13474
rect 11838 13508 11980 13524
rect 11838 13474 11858 13508
rect 11892 13474 11926 13508
rect 11960 13474 11980 13508
rect 11838 13458 11980 13474
rect 12356 13508 12498 13524
rect 12356 13474 12376 13508
rect 12410 13474 12444 13508
rect 12478 13474 12498 13508
rect 12356 13458 12498 13474
rect 12758 13508 12900 13524
rect 12758 13474 12778 13508
rect 12812 13474 12846 13508
rect 12880 13474 12900 13508
rect 12758 13458 12900 13474
rect 3156 9398 3298 9414
rect 3156 9364 3176 9398
rect 3210 9364 3244 9398
rect 3278 9364 3298 9398
rect 3156 9348 3298 9364
rect 3558 9398 3700 9414
rect 3558 9364 3578 9398
rect 3612 9364 3646 9398
rect 3680 9364 3700 9398
rect 3558 9348 3700 9364
rect 4076 9398 4218 9414
rect 4076 9364 4096 9398
rect 4130 9364 4164 9398
rect 4198 9364 4218 9398
rect 4076 9348 4218 9364
rect 4478 9398 4620 9414
rect 4478 9364 4498 9398
rect 4532 9364 4566 9398
rect 4600 9364 4620 9398
rect 4478 9348 4620 9364
rect 4996 9398 5138 9414
rect 4996 9364 5016 9398
rect 5050 9364 5084 9398
rect 5118 9364 5138 9398
rect 4996 9348 5138 9364
rect 5398 9398 5540 9414
rect 5398 9364 5418 9398
rect 5452 9364 5486 9398
rect 5520 9364 5540 9398
rect 5398 9348 5540 9364
rect 5916 9398 6058 9414
rect 5916 9364 5936 9398
rect 5970 9364 6004 9398
rect 6038 9364 6058 9398
rect 5916 9348 6058 9364
rect 6318 9398 6460 9414
rect 6318 9364 6338 9398
rect 6372 9364 6406 9398
rect 6440 9364 6460 9398
rect 6318 9348 6460 9364
rect 6836 9398 6978 9414
rect 6836 9364 6856 9398
rect 6890 9364 6924 9398
rect 6958 9364 6978 9398
rect 6836 9348 6978 9364
rect 7238 9398 7380 9414
rect 7238 9364 7258 9398
rect 7292 9364 7326 9398
rect 7360 9364 7380 9398
rect 7238 9348 7380 9364
rect 7756 9398 7898 9414
rect 7756 9364 7776 9398
rect 7810 9364 7844 9398
rect 7878 9364 7898 9398
rect 7756 9348 7898 9364
rect 8158 9398 8300 9414
rect 8158 9364 8178 9398
rect 8212 9364 8246 9398
rect 8280 9364 8300 9398
rect 8158 9348 8300 9364
rect 8676 9398 8818 9414
rect 8676 9364 8696 9398
rect 8730 9364 8764 9398
rect 8798 9364 8818 9398
rect 8676 9348 8818 9364
rect 9078 9398 9220 9414
rect 9078 9364 9098 9398
rect 9132 9364 9166 9398
rect 9200 9364 9220 9398
rect 9078 9348 9220 9364
rect 9596 9398 9738 9414
rect 9596 9364 9616 9398
rect 9650 9364 9684 9398
rect 9718 9364 9738 9398
rect 9596 9348 9738 9364
rect 9998 9398 10140 9414
rect 9998 9364 10018 9398
rect 10052 9364 10086 9398
rect 10120 9364 10140 9398
rect 9998 9348 10140 9364
rect 10516 9398 10658 9414
rect 10516 9364 10536 9398
rect 10570 9364 10604 9398
rect 10638 9364 10658 9398
rect 10516 9348 10658 9364
rect 10918 9398 11060 9414
rect 10918 9364 10938 9398
rect 10972 9364 11006 9398
rect 11040 9364 11060 9398
rect 10918 9348 11060 9364
rect 11436 9398 11578 9414
rect 11436 9364 11456 9398
rect 11490 9364 11524 9398
rect 11558 9364 11578 9398
rect 11436 9348 11578 9364
rect 11838 9398 11980 9414
rect 11838 9364 11858 9398
rect 11892 9364 11926 9398
rect 11960 9364 11980 9398
rect 11838 9348 11980 9364
rect 12356 9398 12498 9414
rect 12356 9364 12376 9398
rect 12410 9364 12444 9398
rect 12478 9364 12498 9398
rect 12356 9348 12498 9364
rect 12758 9398 12900 9414
rect 12758 9364 12778 9398
rect 12812 9364 12846 9398
rect 12880 9364 12900 9398
rect 12758 9348 12900 9364
rect 1268 7446 9012 7462
rect 1268 7412 1284 7446
rect 1318 7412 1353 7446
rect 1387 7412 1422 7446
rect 1456 7412 1491 7446
rect 1525 7412 1560 7446
rect 1594 7412 1629 7446
rect 1663 7412 1698 7446
rect 1732 7412 1767 7446
rect 1801 7412 1836 7446
rect 1870 7412 1905 7446
rect 1939 7412 1974 7446
rect 2008 7412 2043 7446
rect 2077 7412 2112 7446
rect 2146 7412 2181 7446
rect 2215 7412 2250 7446
rect 2284 7412 2319 7446
rect 2353 7412 2388 7446
rect 2422 7412 2457 7446
rect 2491 7412 2526 7446
rect 2560 7412 2595 7446
rect 2629 7412 2664 7446
rect 2698 7412 2733 7446
rect 2767 7412 2802 7446
rect 2836 7412 2871 7446
rect 2905 7412 2940 7446
rect 2974 7412 3009 7446
rect 3043 7412 3078 7446
rect 3112 7412 3147 7446
rect 3181 7412 3216 7446
rect 3250 7412 3285 7446
rect 3319 7412 3354 7446
rect 3388 7412 3423 7446
rect 3457 7412 3492 7446
rect 3526 7412 3561 7446
rect 3595 7412 3630 7446
rect 3664 7412 3699 7446
rect 3733 7412 3768 7446
rect 3802 7412 3837 7446
rect 3871 7412 3906 7446
rect 3940 7412 3975 7446
rect 4009 7412 4044 7446
rect 4078 7412 4113 7446
rect 4147 7412 4182 7446
rect 4216 7412 4251 7446
rect 4285 7412 4320 7446
rect 4354 7412 4389 7446
rect 4423 7412 4458 7446
rect 4492 7412 4527 7446
rect 4561 7412 4596 7446
rect 4630 7412 4665 7446
rect 4699 7412 4734 7446
rect 4768 7412 4803 7446
rect 4837 7412 4872 7446
rect 4906 7412 4941 7446
rect 4975 7412 5010 7446
rect 5044 7412 5079 7446
rect 5113 7412 5148 7446
rect 5182 7412 5217 7446
rect 5251 7412 5286 7446
rect 5320 7412 5355 7446
rect 5389 7412 5424 7446
rect 5458 7412 5493 7446
rect 5527 7412 5562 7446
rect 5596 7412 5630 7446
rect 5664 7412 5698 7446
rect 5732 7412 5766 7446
rect 5800 7412 5834 7446
rect 5868 7412 5902 7446
rect 5936 7412 5970 7446
rect 6004 7412 6038 7446
rect 6072 7412 6106 7446
rect 6140 7412 6174 7446
rect 6208 7412 6242 7446
rect 6276 7412 6310 7446
rect 6344 7412 6378 7446
rect 6412 7412 6446 7446
rect 6480 7412 6514 7446
rect 6548 7412 6582 7446
rect 6616 7412 6650 7446
rect 6684 7412 6718 7446
rect 6752 7412 6786 7446
rect 6820 7412 6854 7446
rect 6888 7412 6922 7446
rect 6956 7412 6990 7446
rect 7024 7412 7058 7446
rect 7092 7412 7126 7446
rect 7160 7412 7194 7446
rect 7228 7412 7262 7446
rect 7296 7412 7330 7446
rect 7364 7412 7398 7446
rect 7432 7412 7466 7446
rect 7500 7412 7534 7446
rect 7568 7412 7602 7446
rect 7636 7412 7670 7446
rect 7704 7412 7738 7446
rect 7772 7412 7806 7446
rect 7840 7412 7874 7446
rect 7908 7412 7942 7446
rect 7976 7412 8010 7446
rect 8044 7412 8078 7446
rect 8112 7412 8146 7446
rect 8180 7412 8214 7446
rect 8248 7412 8282 7446
rect 8316 7412 8350 7446
rect 8384 7412 8418 7446
rect 8452 7412 8486 7446
rect 8520 7412 8554 7446
rect 8588 7412 8622 7446
rect 8656 7412 8690 7446
rect 8724 7412 8758 7446
rect 8792 7412 8826 7446
rect 8860 7412 8894 7446
rect 8928 7412 8962 7446
rect 8996 7412 9012 7446
rect 1268 7386 9012 7412
rect 10988 7988 13267 8004
rect 10988 7954 11004 7988
rect 11038 7954 11074 7988
rect 11108 7954 11144 7988
rect 11178 7954 11214 7988
rect 11248 7954 11284 7988
rect 11318 7954 11354 7988
rect 11388 7954 11423 7988
rect 11457 7954 11492 7988
rect 11526 7954 11561 7988
rect 11595 7954 11630 7988
rect 11664 7954 11699 7988
rect 11733 7954 11768 7988
rect 11802 7954 11837 7988
rect 11871 7954 11906 7988
rect 11940 7954 11975 7988
rect 12009 7954 12044 7988
rect 12078 7954 12113 7988
rect 12147 7954 12182 7988
rect 12216 7954 12251 7988
rect 12285 7954 12320 7988
rect 12354 7954 12389 7988
rect 12423 7954 12458 7988
rect 12492 7954 12527 7988
rect 12561 7954 12596 7988
rect 12630 7954 12665 7988
rect 12699 7954 12734 7988
rect 12768 7954 12803 7988
rect 12837 7954 12872 7988
rect 12906 7954 12941 7988
rect 12975 7954 13010 7988
rect 13044 7954 13079 7988
rect 13113 7954 13148 7988
rect 13182 7954 13217 7988
rect 13251 7954 13267 7988
rect 10988 7938 13267 7954
rect 11563 4387 12363 4403
rect 11563 4353 11629 4387
rect 11663 4353 11697 4387
rect 11731 4353 11765 4387
rect 11799 4353 11833 4387
rect 11867 4353 11901 4387
rect 11935 4353 11969 4387
rect 12003 4353 12037 4387
rect 12071 4353 12105 4387
rect 12139 4353 12173 4387
rect 12207 4353 12241 4387
rect 12275 4353 12309 4387
rect 12343 4353 12363 4387
rect 11563 4337 12363 4353
<< polycont >>
rect 3176 39074 3210 39108
rect 3244 39074 3278 39108
rect 3578 39074 3612 39108
rect 3646 39074 3680 39108
rect 4096 39074 4130 39108
rect 4164 39074 4198 39108
rect 4498 39074 4532 39108
rect 4566 39074 4600 39108
rect 5016 39074 5050 39108
rect 5084 39074 5118 39108
rect 5418 39074 5452 39108
rect 5486 39074 5520 39108
rect 5936 39074 5970 39108
rect 6004 39074 6038 39108
rect 6338 39074 6372 39108
rect 6406 39074 6440 39108
rect 6856 39074 6890 39108
rect 6924 39074 6958 39108
rect 7258 39074 7292 39108
rect 7326 39074 7360 39108
rect 7776 39074 7810 39108
rect 7844 39074 7878 39108
rect 8178 39074 8212 39108
rect 8246 39074 8280 39108
rect 8696 39074 8730 39108
rect 8764 39074 8798 39108
rect 9098 39074 9132 39108
rect 9166 39074 9200 39108
rect 9616 39074 9650 39108
rect 9684 39074 9718 39108
rect 10018 39074 10052 39108
rect 10086 39074 10120 39108
rect 10536 39074 10570 39108
rect 10604 39074 10638 39108
rect 10938 39074 10972 39108
rect 11006 39074 11040 39108
rect 11456 39074 11490 39108
rect 11524 39074 11558 39108
rect 11858 39074 11892 39108
rect 11926 39074 11960 39108
rect 12376 39074 12410 39108
rect 12444 39074 12478 39108
rect 12778 39074 12812 39108
rect 12846 39074 12880 39108
rect 3176 36964 3210 36998
rect 3244 36964 3278 36998
rect 3578 36964 3612 36998
rect 3646 36964 3680 36998
rect 4096 36964 4130 36998
rect 4164 36964 4198 36998
rect 4498 36964 4532 36998
rect 4566 36964 4600 36998
rect 5016 36964 5050 36998
rect 5084 36964 5118 36998
rect 5418 36964 5452 36998
rect 5486 36964 5520 36998
rect 5936 36964 5970 36998
rect 6004 36964 6038 36998
rect 6338 36964 6372 36998
rect 6406 36964 6440 36998
rect 6856 36964 6890 36998
rect 6924 36964 6958 36998
rect 7258 36964 7292 36998
rect 7326 36964 7360 36998
rect 7776 36964 7810 36998
rect 7844 36964 7878 36998
rect 8178 36964 8212 36998
rect 8246 36964 8280 36998
rect 8696 36964 8730 36998
rect 8764 36964 8798 36998
rect 9098 36964 9132 36998
rect 9166 36964 9200 36998
rect 9616 36964 9650 36998
rect 9684 36964 9718 36998
rect 10018 36964 10052 36998
rect 10086 36964 10120 36998
rect 10536 36964 10570 36998
rect 10604 36964 10638 36998
rect 10938 36964 10972 36998
rect 11006 36964 11040 36998
rect 11456 36964 11490 36998
rect 11524 36964 11558 36998
rect 11858 36964 11892 36998
rect 11926 36964 11960 36998
rect 12376 36964 12410 36998
rect 12444 36964 12478 36998
rect 12778 36964 12812 36998
rect 12846 36964 12880 36998
rect 3176 36474 3210 36508
rect 3244 36474 3278 36508
rect 3578 36474 3612 36508
rect 3646 36474 3680 36508
rect 4096 36474 4130 36508
rect 4164 36474 4198 36508
rect 4498 36474 4532 36508
rect 4566 36474 4600 36508
rect 5016 36474 5050 36508
rect 5084 36474 5118 36508
rect 5418 36474 5452 36508
rect 5486 36474 5520 36508
rect 5936 36474 5970 36508
rect 6004 36474 6038 36508
rect 6338 36474 6372 36508
rect 6406 36474 6440 36508
rect 6856 36474 6890 36508
rect 6924 36474 6958 36508
rect 7258 36474 7292 36508
rect 7326 36474 7360 36508
rect 7776 36474 7810 36508
rect 7844 36474 7878 36508
rect 8178 36474 8212 36508
rect 8246 36474 8280 36508
rect 8696 36474 8730 36508
rect 8764 36474 8798 36508
rect 9098 36474 9132 36508
rect 9166 36474 9200 36508
rect 9616 36474 9650 36508
rect 9684 36474 9718 36508
rect 10018 36474 10052 36508
rect 10086 36474 10120 36508
rect 10536 36474 10570 36508
rect 10604 36474 10638 36508
rect 10938 36474 10972 36508
rect 11006 36474 11040 36508
rect 11456 36474 11490 36508
rect 11524 36474 11558 36508
rect 11858 36474 11892 36508
rect 11926 36474 11960 36508
rect 12376 36474 12410 36508
rect 12444 36474 12478 36508
rect 12778 36474 12812 36508
rect 12846 36474 12880 36508
rect 3176 32364 3210 32398
rect 3244 32364 3278 32398
rect 3578 32364 3612 32398
rect 3646 32364 3680 32398
rect 4096 32364 4130 32398
rect 4164 32364 4198 32398
rect 4498 32364 4532 32398
rect 4566 32364 4600 32398
rect 5016 32364 5050 32398
rect 5084 32364 5118 32398
rect 5418 32364 5452 32398
rect 5486 32364 5520 32398
rect 5936 32364 5970 32398
rect 6004 32364 6038 32398
rect 6338 32364 6372 32398
rect 6406 32364 6440 32398
rect 6856 32364 6890 32398
rect 6924 32364 6958 32398
rect 7258 32364 7292 32398
rect 7326 32364 7360 32398
rect 7776 32364 7810 32398
rect 7844 32364 7878 32398
rect 8178 32364 8212 32398
rect 8246 32364 8280 32398
rect 8696 32364 8730 32398
rect 8764 32364 8798 32398
rect 9098 32364 9132 32398
rect 9166 32364 9200 32398
rect 9616 32364 9650 32398
rect 9684 32364 9718 32398
rect 10018 32364 10052 32398
rect 10086 32364 10120 32398
rect 10536 32364 10570 32398
rect 10604 32364 10638 32398
rect 10938 32364 10972 32398
rect 11006 32364 11040 32398
rect 11456 32364 11490 32398
rect 11524 32364 11558 32398
rect 11858 32364 11892 32398
rect 11926 32364 11960 32398
rect 12376 32364 12410 32398
rect 12444 32364 12478 32398
rect 12778 32364 12812 32398
rect 12846 32364 12880 32398
rect 3176 31874 3210 31908
rect 3244 31874 3278 31908
rect 3578 31874 3612 31908
rect 3646 31874 3680 31908
rect 4096 31874 4130 31908
rect 4164 31874 4198 31908
rect 4498 31874 4532 31908
rect 4566 31874 4600 31908
rect 5016 31874 5050 31908
rect 5084 31874 5118 31908
rect 5418 31874 5452 31908
rect 5486 31874 5520 31908
rect 5936 31874 5970 31908
rect 6004 31874 6038 31908
rect 6338 31874 6372 31908
rect 6406 31874 6440 31908
rect 6856 31874 6890 31908
rect 6924 31874 6958 31908
rect 7258 31874 7292 31908
rect 7326 31874 7360 31908
rect 7776 31874 7810 31908
rect 7844 31874 7878 31908
rect 8178 31874 8212 31908
rect 8246 31874 8280 31908
rect 8696 31874 8730 31908
rect 8764 31874 8798 31908
rect 9098 31874 9132 31908
rect 9166 31874 9200 31908
rect 9616 31874 9650 31908
rect 9684 31874 9718 31908
rect 10018 31874 10052 31908
rect 10086 31874 10120 31908
rect 10536 31874 10570 31908
rect 10604 31874 10638 31908
rect 10938 31874 10972 31908
rect 11006 31874 11040 31908
rect 11456 31874 11490 31908
rect 11524 31874 11558 31908
rect 11858 31874 11892 31908
rect 11926 31874 11960 31908
rect 12376 31874 12410 31908
rect 12444 31874 12478 31908
rect 12778 31874 12812 31908
rect 12846 31874 12880 31908
rect 3176 27764 3210 27798
rect 3244 27764 3278 27798
rect 3578 27764 3612 27798
rect 3646 27764 3680 27798
rect 4096 27764 4130 27798
rect 4164 27764 4198 27798
rect 4498 27764 4532 27798
rect 4566 27764 4600 27798
rect 5016 27764 5050 27798
rect 5084 27764 5118 27798
rect 5418 27764 5452 27798
rect 5486 27764 5520 27798
rect 5936 27764 5970 27798
rect 6004 27764 6038 27798
rect 6338 27764 6372 27798
rect 6406 27764 6440 27798
rect 6856 27764 6890 27798
rect 6924 27764 6958 27798
rect 7258 27764 7292 27798
rect 7326 27764 7360 27798
rect 7776 27764 7810 27798
rect 7844 27764 7878 27798
rect 8178 27764 8212 27798
rect 8246 27764 8280 27798
rect 8696 27764 8730 27798
rect 8764 27764 8798 27798
rect 9098 27764 9132 27798
rect 9166 27764 9200 27798
rect 9616 27764 9650 27798
rect 9684 27764 9718 27798
rect 10018 27764 10052 27798
rect 10086 27764 10120 27798
rect 10536 27764 10570 27798
rect 10604 27764 10638 27798
rect 10938 27764 10972 27798
rect 11006 27764 11040 27798
rect 11456 27764 11490 27798
rect 11524 27764 11558 27798
rect 11858 27764 11892 27798
rect 11926 27764 11960 27798
rect 12376 27764 12410 27798
rect 12444 27764 12478 27798
rect 12778 27764 12812 27798
rect 12846 27764 12880 27798
rect 5016 27274 5050 27308
rect 5084 27274 5118 27308
rect 5418 27274 5452 27308
rect 5486 27274 5520 27308
rect 5936 27274 5970 27308
rect 6004 27274 6038 27308
rect 6338 27274 6372 27308
rect 6406 27274 6440 27308
rect 6856 27274 6890 27308
rect 6924 27274 6958 27308
rect 7258 27274 7292 27308
rect 7326 27274 7360 27308
rect 7776 27274 7810 27308
rect 7844 27274 7878 27308
rect 8178 27274 8212 27308
rect 8246 27274 8280 27308
rect 8696 27274 8730 27308
rect 8764 27274 8798 27308
rect 9098 27274 9132 27308
rect 9166 27274 9200 27308
rect 9616 27274 9650 27308
rect 9684 27274 9718 27308
rect 10018 27274 10052 27308
rect 10086 27274 10120 27308
rect 10536 27274 10570 27308
rect 10604 27274 10638 27308
rect 10938 27274 10972 27308
rect 11006 27274 11040 27308
rect 11456 27274 11490 27308
rect 11524 27274 11558 27308
rect 11858 27274 11892 27308
rect 11926 27274 11960 27308
rect 12376 27274 12410 27308
rect 12444 27274 12478 27308
rect 12778 27274 12812 27308
rect 12846 27274 12880 27308
rect 5016 23164 5050 23198
rect 5084 23164 5118 23198
rect 5418 23164 5452 23198
rect 5486 23164 5520 23198
rect 5936 23164 5970 23198
rect 6004 23164 6038 23198
rect 6338 23164 6372 23198
rect 6406 23164 6440 23198
rect 6856 23164 6890 23198
rect 6924 23164 6958 23198
rect 7258 23164 7292 23198
rect 7326 23164 7360 23198
rect 7776 23164 7810 23198
rect 7844 23164 7878 23198
rect 8178 23164 8212 23198
rect 8246 23164 8280 23198
rect 8696 23164 8730 23198
rect 8764 23164 8798 23198
rect 9098 23164 9132 23198
rect 9166 23164 9200 23198
rect 9616 23164 9650 23198
rect 9684 23164 9718 23198
rect 10018 23164 10052 23198
rect 10086 23164 10120 23198
rect 10536 23164 10570 23198
rect 10604 23164 10638 23198
rect 10938 23164 10972 23198
rect 11006 23164 11040 23198
rect 11456 23164 11490 23198
rect 11524 23164 11558 23198
rect 11858 23164 11892 23198
rect 11926 23164 11960 23198
rect 12376 23164 12410 23198
rect 12444 23164 12478 23198
rect 12778 23164 12812 23198
rect 12846 23164 12880 23198
rect 5016 22674 5050 22708
rect 5084 22674 5118 22708
rect 5418 22674 5452 22708
rect 5486 22674 5520 22708
rect 5936 22674 5970 22708
rect 6004 22674 6038 22708
rect 6338 22674 6372 22708
rect 6406 22674 6440 22708
rect 6856 22674 6890 22708
rect 6924 22674 6958 22708
rect 7258 22674 7292 22708
rect 7326 22674 7360 22708
rect 7776 22674 7810 22708
rect 7844 22674 7878 22708
rect 8178 22674 8212 22708
rect 8246 22674 8280 22708
rect 8696 22674 8730 22708
rect 8764 22674 8798 22708
rect 9098 22674 9132 22708
rect 9166 22674 9200 22708
rect 9616 22674 9650 22708
rect 9684 22674 9718 22708
rect 10018 22674 10052 22708
rect 10086 22674 10120 22708
rect 10536 22674 10570 22708
rect 10604 22674 10638 22708
rect 10938 22674 10972 22708
rect 11006 22674 11040 22708
rect 11456 22674 11490 22708
rect 11524 22674 11558 22708
rect 11858 22674 11892 22708
rect 11926 22674 11960 22708
rect 12376 22674 12410 22708
rect 12444 22674 12478 22708
rect 12778 22674 12812 22708
rect 12846 22674 12880 22708
rect 5016 18564 5050 18598
rect 5084 18564 5118 18598
rect 5418 18564 5452 18598
rect 5486 18564 5520 18598
rect 5936 18564 5970 18598
rect 6004 18564 6038 18598
rect 6338 18564 6372 18598
rect 6406 18564 6440 18598
rect 6856 18564 6890 18598
rect 6924 18564 6958 18598
rect 7258 18564 7292 18598
rect 7326 18564 7360 18598
rect 7776 18564 7810 18598
rect 7844 18564 7878 18598
rect 8178 18564 8212 18598
rect 8246 18564 8280 18598
rect 8696 18564 8730 18598
rect 8764 18564 8798 18598
rect 9098 18564 9132 18598
rect 9166 18564 9200 18598
rect 9616 18564 9650 18598
rect 9684 18564 9718 18598
rect 10018 18564 10052 18598
rect 10086 18564 10120 18598
rect 10536 18564 10570 18598
rect 10604 18564 10638 18598
rect 10938 18564 10972 18598
rect 11006 18564 11040 18598
rect 11456 18564 11490 18598
rect 11524 18564 11558 18598
rect 11858 18564 11892 18598
rect 11926 18564 11960 18598
rect 12376 18564 12410 18598
rect 12444 18564 12478 18598
rect 12778 18564 12812 18598
rect 12846 18564 12880 18598
rect 5016 18074 5050 18108
rect 5084 18074 5118 18108
rect 5418 18074 5452 18108
rect 5486 18074 5520 18108
rect 5936 18074 5970 18108
rect 6004 18074 6038 18108
rect 6338 18074 6372 18108
rect 6406 18074 6440 18108
rect 6856 18074 6890 18108
rect 6924 18074 6958 18108
rect 7258 18074 7292 18108
rect 7326 18074 7360 18108
rect 7776 18074 7810 18108
rect 7844 18074 7878 18108
rect 8178 18074 8212 18108
rect 8246 18074 8280 18108
rect 8696 18074 8730 18108
rect 8764 18074 8798 18108
rect 9098 18074 9132 18108
rect 9166 18074 9200 18108
rect 9616 18074 9650 18108
rect 9684 18074 9718 18108
rect 10018 18074 10052 18108
rect 10086 18074 10120 18108
rect 10536 18074 10570 18108
rect 10604 18074 10638 18108
rect 10938 18074 10972 18108
rect 11006 18074 11040 18108
rect 11456 18074 11490 18108
rect 11524 18074 11558 18108
rect 11858 18074 11892 18108
rect 11926 18074 11960 18108
rect 12376 18074 12410 18108
rect 12444 18074 12478 18108
rect 12778 18074 12812 18108
rect 12846 18074 12880 18108
rect 5016 13964 5050 13998
rect 5084 13964 5118 13998
rect 5418 13964 5452 13998
rect 5486 13964 5520 13998
rect 5936 13964 5970 13998
rect 6004 13964 6038 13998
rect 6338 13964 6372 13998
rect 6406 13964 6440 13998
rect 6856 13964 6890 13998
rect 6924 13964 6958 13998
rect 7258 13964 7292 13998
rect 7326 13964 7360 13998
rect 7776 13964 7810 13998
rect 7844 13964 7878 13998
rect 8178 13964 8212 13998
rect 8246 13964 8280 13998
rect 8696 13964 8730 13998
rect 8764 13964 8798 13998
rect 9098 13964 9132 13998
rect 9166 13964 9200 13998
rect 9616 13964 9650 13998
rect 9684 13964 9718 13998
rect 10018 13964 10052 13998
rect 10086 13964 10120 13998
rect 10536 13964 10570 13998
rect 10604 13964 10638 13998
rect 10938 13964 10972 13998
rect 11006 13964 11040 13998
rect 11456 13964 11490 13998
rect 11524 13964 11558 13998
rect 11858 13964 11892 13998
rect 11926 13964 11960 13998
rect 12376 13964 12410 13998
rect 12444 13964 12478 13998
rect 12778 13964 12812 13998
rect 12846 13964 12880 13998
rect 3176 13474 3210 13508
rect 3244 13474 3278 13508
rect 3578 13474 3612 13508
rect 3646 13474 3680 13508
rect 4096 13474 4130 13508
rect 4164 13474 4198 13508
rect 4498 13474 4532 13508
rect 4566 13474 4600 13508
rect 5016 13474 5050 13508
rect 5084 13474 5118 13508
rect 5418 13474 5452 13508
rect 5486 13474 5520 13508
rect 5936 13474 5970 13508
rect 6004 13474 6038 13508
rect 6338 13474 6372 13508
rect 6406 13474 6440 13508
rect 6856 13474 6890 13508
rect 6924 13474 6958 13508
rect 7258 13474 7292 13508
rect 7326 13474 7360 13508
rect 7776 13474 7810 13508
rect 7844 13474 7878 13508
rect 8178 13474 8212 13508
rect 8246 13474 8280 13508
rect 8696 13474 8730 13508
rect 8764 13474 8798 13508
rect 9098 13474 9132 13508
rect 9166 13474 9200 13508
rect 9616 13474 9650 13508
rect 9684 13474 9718 13508
rect 10018 13474 10052 13508
rect 10086 13474 10120 13508
rect 10536 13474 10570 13508
rect 10604 13474 10638 13508
rect 10938 13474 10972 13508
rect 11006 13474 11040 13508
rect 11456 13474 11490 13508
rect 11524 13474 11558 13508
rect 11858 13474 11892 13508
rect 11926 13474 11960 13508
rect 12376 13474 12410 13508
rect 12444 13474 12478 13508
rect 12778 13474 12812 13508
rect 12846 13474 12880 13508
rect 3176 9364 3210 9398
rect 3244 9364 3278 9398
rect 3578 9364 3612 9398
rect 3646 9364 3680 9398
rect 4096 9364 4130 9398
rect 4164 9364 4198 9398
rect 4498 9364 4532 9398
rect 4566 9364 4600 9398
rect 5016 9364 5050 9398
rect 5084 9364 5118 9398
rect 5418 9364 5452 9398
rect 5486 9364 5520 9398
rect 5936 9364 5970 9398
rect 6004 9364 6038 9398
rect 6338 9364 6372 9398
rect 6406 9364 6440 9398
rect 6856 9364 6890 9398
rect 6924 9364 6958 9398
rect 7258 9364 7292 9398
rect 7326 9364 7360 9398
rect 7776 9364 7810 9398
rect 7844 9364 7878 9398
rect 8178 9364 8212 9398
rect 8246 9364 8280 9398
rect 8696 9364 8730 9398
rect 8764 9364 8798 9398
rect 9098 9364 9132 9398
rect 9166 9364 9200 9398
rect 9616 9364 9650 9398
rect 9684 9364 9718 9398
rect 10018 9364 10052 9398
rect 10086 9364 10120 9398
rect 10536 9364 10570 9398
rect 10604 9364 10638 9398
rect 10938 9364 10972 9398
rect 11006 9364 11040 9398
rect 11456 9364 11490 9398
rect 11524 9364 11558 9398
rect 11858 9364 11892 9398
rect 11926 9364 11960 9398
rect 12376 9364 12410 9398
rect 12444 9364 12478 9398
rect 12778 9364 12812 9398
rect 12846 9364 12880 9398
rect 1284 7412 1318 7446
rect 1353 7412 1387 7446
rect 1422 7412 1456 7446
rect 1491 7412 1525 7446
rect 1560 7412 1594 7446
rect 1629 7412 1663 7446
rect 1698 7412 1732 7446
rect 1767 7412 1801 7446
rect 1836 7412 1870 7446
rect 1905 7412 1939 7446
rect 1974 7412 2008 7446
rect 2043 7412 2077 7446
rect 2112 7412 2146 7446
rect 2181 7412 2215 7446
rect 2250 7412 2284 7446
rect 2319 7412 2353 7446
rect 2388 7412 2422 7446
rect 2457 7412 2491 7446
rect 2526 7412 2560 7446
rect 2595 7412 2629 7446
rect 2664 7412 2698 7446
rect 2733 7412 2767 7446
rect 2802 7412 2836 7446
rect 2871 7412 2905 7446
rect 2940 7412 2974 7446
rect 3009 7412 3043 7446
rect 3078 7412 3112 7446
rect 3147 7412 3181 7446
rect 3216 7412 3250 7446
rect 3285 7412 3319 7446
rect 3354 7412 3388 7446
rect 3423 7412 3457 7446
rect 3492 7412 3526 7446
rect 3561 7412 3595 7446
rect 3630 7412 3664 7446
rect 3699 7412 3733 7446
rect 3768 7412 3802 7446
rect 3837 7412 3871 7446
rect 3906 7412 3940 7446
rect 3975 7412 4009 7446
rect 4044 7412 4078 7446
rect 4113 7412 4147 7446
rect 4182 7412 4216 7446
rect 4251 7412 4285 7446
rect 4320 7412 4354 7446
rect 4389 7412 4423 7446
rect 4458 7412 4492 7446
rect 4527 7412 4561 7446
rect 4596 7412 4630 7446
rect 4665 7412 4699 7446
rect 4734 7412 4768 7446
rect 4803 7412 4837 7446
rect 4872 7412 4906 7446
rect 4941 7412 4975 7446
rect 5010 7412 5044 7446
rect 5079 7412 5113 7446
rect 5148 7412 5182 7446
rect 5217 7412 5251 7446
rect 5286 7412 5320 7446
rect 5355 7412 5389 7446
rect 5424 7412 5458 7446
rect 5493 7412 5527 7446
rect 5562 7412 5596 7446
rect 5630 7412 5664 7446
rect 5698 7412 5732 7446
rect 5766 7412 5800 7446
rect 5834 7412 5868 7446
rect 5902 7412 5936 7446
rect 5970 7412 6004 7446
rect 6038 7412 6072 7446
rect 6106 7412 6140 7446
rect 6174 7412 6208 7446
rect 6242 7412 6276 7446
rect 6310 7412 6344 7446
rect 6378 7412 6412 7446
rect 6446 7412 6480 7446
rect 6514 7412 6548 7446
rect 6582 7412 6616 7446
rect 6650 7412 6684 7446
rect 6718 7412 6752 7446
rect 6786 7412 6820 7446
rect 6854 7412 6888 7446
rect 6922 7412 6956 7446
rect 6990 7412 7024 7446
rect 7058 7412 7092 7446
rect 7126 7412 7160 7446
rect 7194 7412 7228 7446
rect 7262 7412 7296 7446
rect 7330 7412 7364 7446
rect 7398 7412 7432 7446
rect 7466 7412 7500 7446
rect 7534 7412 7568 7446
rect 7602 7412 7636 7446
rect 7670 7412 7704 7446
rect 7738 7412 7772 7446
rect 7806 7412 7840 7446
rect 7874 7412 7908 7446
rect 7942 7412 7976 7446
rect 8010 7412 8044 7446
rect 8078 7412 8112 7446
rect 8146 7412 8180 7446
rect 8214 7412 8248 7446
rect 8282 7412 8316 7446
rect 8350 7412 8384 7446
rect 8418 7412 8452 7446
rect 8486 7412 8520 7446
rect 8554 7412 8588 7446
rect 8622 7412 8656 7446
rect 8690 7412 8724 7446
rect 8758 7412 8792 7446
rect 8826 7412 8860 7446
rect 8894 7412 8928 7446
rect 8962 7412 8996 7446
rect 11004 7954 11038 7988
rect 11074 7954 11108 7988
rect 11144 7954 11178 7988
rect 11214 7954 11248 7988
rect 11284 7954 11318 7988
rect 11354 7954 11388 7988
rect 11423 7954 11457 7988
rect 11492 7954 11526 7988
rect 11561 7954 11595 7988
rect 11630 7954 11664 7988
rect 11699 7954 11733 7988
rect 11768 7954 11802 7988
rect 11837 7954 11871 7988
rect 11906 7954 11940 7988
rect 11975 7954 12009 7988
rect 12044 7954 12078 7988
rect 12113 7954 12147 7988
rect 12182 7954 12216 7988
rect 12251 7954 12285 7988
rect 12320 7954 12354 7988
rect 12389 7954 12423 7988
rect 12458 7954 12492 7988
rect 12527 7954 12561 7988
rect 12596 7954 12630 7988
rect 12665 7954 12699 7988
rect 12734 7954 12768 7988
rect 12803 7954 12837 7988
rect 12872 7954 12906 7988
rect 12941 7954 12975 7988
rect 13010 7954 13044 7988
rect 13079 7954 13113 7988
rect 13148 7954 13182 7988
rect 13217 7954 13251 7988
rect 11629 4353 11663 4387
rect 11697 4353 11731 4387
rect 11765 4353 11799 4387
rect 11833 4353 11867 4387
rect 11901 4353 11935 4387
rect 11969 4353 12003 4387
rect 12037 4353 12071 4387
rect 12105 4353 12139 4387
rect 12173 4353 12207 4387
rect 12241 4353 12275 4387
rect 12309 4353 12343 4387
<< locali >>
rect 1830 39905 1902 39939
rect 1936 39933 1975 39939
rect 2009 39933 2048 39939
rect 2082 39933 2121 39939
rect 2155 39933 2194 39939
rect 2228 39933 2267 39939
rect 2301 39933 2340 39939
rect 2374 39933 2413 39939
rect 2447 39933 2486 39939
rect 2520 39933 2559 39939
rect 2593 39933 2632 39939
rect 2666 39933 2705 39939
rect 2739 39933 2778 39939
rect 2812 39933 2851 39939
rect 2885 39933 2924 39939
rect 2958 39933 2997 39939
rect 3031 39933 3070 39939
rect 3104 39933 3143 39939
rect 3177 39933 3216 39939
rect 3250 39933 3289 39939
rect 3323 39933 3362 39939
rect 3396 39933 3435 39939
rect 3469 39933 3508 39939
rect 3542 39933 3581 39939
rect 3615 39933 3654 39939
rect 3688 39933 3727 39939
rect 3761 39933 3800 39939
rect 3834 39933 3873 39939
rect 3907 39933 3946 39939
rect 3980 39933 4019 39939
rect 4053 39933 4092 39939
rect 4126 39933 4165 39939
rect 4199 39933 4238 39939
rect 4272 39933 4311 39939
rect 4345 39933 4384 39939
rect 4418 39933 4457 39939
rect 4491 39933 4530 39939
rect 4564 39933 4603 39939
rect 4637 39933 4676 39939
rect 4710 39933 4749 39939
rect 4783 39933 4822 39939
rect 4856 39933 4895 39939
rect 4929 39933 4968 39939
rect 5002 39933 5041 39939
rect 5075 39933 5114 39939
rect 5148 39933 5187 39939
rect 5221 39933 5260 39939
rect 5294 39933 5333 39939
rect 5367 39933 5406 39939
rect 5440 39933 5479 39939
rect 5513 39933 5552 39939
rect 5586 39933 5625 39939
rect 5659 39933 5698 39939
rect 5732 39933 5771 39939
rect 5805 39933 5844 39939
rect 5878 39933 5917 39939
rect 5951 39933 5990 39939
rect 6024 39933 6063 39939
rect 6097 39933 6136 39939
rect 6170 39933 6209 39939
rect 6243 39933 6282 39939
rect 6316 39933 6355 39939
rect 6389 39933 6428 39939
rect 6462 39933 6501 39939
rect 6535 39933 6574 39939
rect 6608 39933 6647 39939
rect 1936 39905 1949 39933
rect 2009 39905 2017 39933
rect 1830 39899 1949 39905
rect 1983 39899 2017 39905
rect 1830 39867 2017 39899
rect 1936 39833 1975 39867
rect 2009 39833 2017 39867
rect 13953 39867 14025 39939
rect 13953 39833 13991 39867
rect 14483 39842 14521 39876
rect 1936 39831 2017 39833
rect 1936 39797 2085 39831
rect 2004 39795 2085 39797
rect 2008 39761 2047 39795
rect 2081 39763 2085 39795
rect 2081 39761 2120 39763
rect 13951 39831 14025 39833
rect 13883 39812 14025 39831
rect 13883 39794 13985 39812
rect 14019 39794 14025 39812
rect 13883 39763 13919 39794
rect 13881 39761 13919 39763
rect 2008 39729 2153 39761
rect 2072 39723 2153 39729
rect 2080 39689 2119 39723
rect 13815 39760 13919 39761
rect 13953 39778 13985 39794
rect 13953 39760 13991 39778
rect 13815 39744 14025 39760
rect 13815 39722 13917 39744
rect 13815 39695 13847 39722
rect 2153 39689 2192 39695
rect 2226 39689 2265 39695
rect 2299 39689 2338 39695
rect 2372 39689 2411 39695
rect 2445 39689 2484 39695
rect 2518 39689 2557 39695
rect 2591 39689 2630 39695
rect 2664 39689 2703 39695
rect 2737 39689 2776 39695
rect 2810 39689 2849 39695
rect 2883 39689 2922 39695
rect 2956 39689 2995 39695
rect 3029 39689 3068 39695
rect 3102 39689 3141 39695
rect 3175 39689 3214 39695
rect 3248 39689 3287 39695
rect 3321 39689 3360 39695
rect 3394 39689 3433 39695
rect 3467 39689 3506 39695
rect 3540 39689 3579 39695
rect 3613 39689 3652 39695
rect 3686 39689 3725 39695
rect 3759 39689 3798 39695
rect 3832 39689 3871 39695
rect 3905 39689 3944 39695
rect 3978 39689 4017 39695
rect 4051 39689 4090 39695
rect 4124 39689 4163 39695
rect 4197 39689 4236 39695
rect 4270 39689 4309 39695
rect 4343 39689 4382 39695
rect 4416 39689 4455 39695
rect 4489 39689 4528 39695
rect 4562 39689 4601 39695
rect 4635 39689 4674 39695
rect 4708 39689 4747 39695
rect 4781 39689 4820 39695
rect 4854 39689 4893 39695
rect 4927 39689 4966 39695
rect 5000 39689 5039 39695
rect 5073 39689 5112 39695
rect 5146 39689 5185 39695
rect 5219 39689 5258 39695
rect 5292 39689 5331 39695
rect 5365 39689 5404 39695
rect 5438 39689 5477 39695
rect 5511 39689 5550 39695
rect 5584 39689 5623 39695
rect 5657 39689 5696 39695
rect 5730 39689 5769 39695
rect 5803 39689 5842 39695
rect 5876 39689 5915 39695
rect 5949 39689 5988 39695
rect 6022 39689 6061 39695
rect 6095 39689 6134 39695
rect 6168 39689 6207 39695
rect 6241 39689 6280 39695
rect 6314 39689 6353 39695
rect 6387 39689 6426 39695
rect 6460 39689 6499 39695
rect 6533 39689 6572 39695
rect 6606 39689 6645 39695
rect 6679 39689 6718 39695
rect 6752 39689 6791 39695
rect 13809 39689 13847 39695
rect 13775 39688 13847 39689
rect 13881 39688 13917 39722
rect 14019 39721 14025 39744
rect 13775 39676 13917 39688
rect 13775 39650 13849 39676
rect 13809 39649 13849 39650
rect 13809 39616 13847 39649
rect 13775 39615 13847 39616
rect 14019 39648 14025 39687
rect 13775 39608 13849 39615
rect 13775 39577 13781 39608
rect 1830 35834 1834 35873
rect 2072 35834 2080 35873
rect 1830 35761 1834 35800
rect 2072 35761 2080 35800
rect 1830 35688 1834 35727
rect 2072 35688 2080 35727
rect 1830 35615 1834 35654
rect 2072 35615 2080 35654
rect 1830 35542 1834 35581
rect 2072 35542 2080 35581
rect 1830 35469 1834 35508
rect 2072 35469 2080 35508
rect 1830 35396 1834 35435
rect 2072 35396 2080 35435
rect 1830 35323 1834 35362
rect 2072 35323 2080 35362
rect 1830 35250 1834 35289
rect 2072 35250 2080 35289
rect 1830 35177 1834 35216
rect 2072 35177 2080 35216
rect 1830 35104 1834 35143
rect 2072 35104 2080 35143
rect 1830 35031 1834 35070
rect 2072 35031 2080 35070
rect 1830 34958 1834 34997
rect 2072 34958 2080 34997
rect 1830 34885 1834 34924
rect 2072 34885 2080 34924
rect 1830 34812 1834 34851
rect 2072 34812 2080 34851
rect 1830 34739 1834 34778
rect 2072 34739 2080 34778
rect 1830 34666 1834 34705
rect 2072 34666 2080 34705
rect 1830 34593 1834 34632
rect 2072 34593 2080 34632
rect 1830 34520 1834 34559
rect 2072 34520 2080 34559
rect 1830 34447 1834 34486
rect 2072 34447 2080 34486
rect 1830 34374 1834 34413
rect 2072 34374 2080 34413
rect 1830 34301 1834 34340
rect 2072 34301 2080 34340
rect 1830 34228 1834 34267
rect 2072 34228 2080 34267
rect 2220 39511 2292 39545
rect 2326 39542 2365 39545
rect 13559 39542 13631 39545
rect 2220 39508 2306 39511
rect 2340 39508 2365 39542
rect 2220 39474 2365 39508
rect 2220 39473 2225 39474
rect 2327 39439 2365 39474
rect 13560 39473 13631 39542
rect 13560 39458 13597 39473
rect 13560 39440 13594 39458
rect 13559 39439 13594 39440
rect 2327 39406 2437 39439
rect 2395 39401 2437 39406
rect 2398 39367 2437 39401
rect 13492 39424 13594 39439
rect 13628 39424 13631 39439
rect 13492 39400 13631 39424
rect 13492 39372 13525 39400
rect 13559 39390 13597 39400
rect 13487 39367 13525 39372
rect 13453 39366 13525 39367
rect 13453 39328 13526 39366
rect 13487 39327 13526 39328
rect 13628 39327 13631 39366
rect 13487 39322 13525 39327
rect 13453 39255 13458 39294
rect 13628 39254 13631 39293
rect 13453 39182 13458 39221
rect 13628 39181 13631 39220
rect 13453 39109 13458 39148
rect 3156 39074 3176 39108
rect 3210 39074 3244 39108
rect 3282 39074 3298 39108
rect 3558 39074 3578 39108
rect 3612 39074 3646 39108
rect 3684 39074 3700 39108
rect 4076 39074 4096 39108
rect 4130 39074 4164 39108
rect 4202 39074 4218 39108
rect 4478 39074 4498 39108
rect 4532 39074 4566 39108
rect 4604 39074 4620 39108
rect 4996 39074 5016 39108
rect 5050 39074 5084 39108
rect 5122 39074 5138 39108
rect 5398 39074 5418 39108
rect 5452 39074 5486 39108
rect 5524 39074 5540 39108
rect 5916 39074 5936 39108
rect 5970 39074 6004 39108
rect 6042 39074 6058 39108
rect 6318 39074 6338 39108
rect 6372 39074 6406 39108
rect 6444 39074 6460 39108
rect 6836 39074 6856 39108
rect 6890 39074 6924 39108
rect 6962 39074 6978 39108
rect 7238 39074 7258 39108
rect 7292 39074 7326 39108
rect 7364 39074 7380 39108
rect 7756 39074 7776 39108
rect 7810 39074 7844 39108
rect 7882 39074 7898 39108
rect 8158 39074 8178 39108
rect 8212 39074 8246 39108
rect 8284 39074 8300 39108
rect 8676 39074 8696 39108
rect 8730 39074 8764 39108
rect 8802 39074 8818 39108
rect 9078 39074 9098 39108
rect 9132 39074 9166 39108
rect 9204 39074 9220 39108
rect 9596 39074 9616 39108
rect 9650 39074 9684 39108
rect 9722 39074 9738 39108
rect 9998 39074 10018 39108
rect 10052 39074 10086 39108
rect 10124 39074 10140 39108
rect 10516 39074 10536 39108
rect 10570 39074 10604 39108
rect 10642 39074 10658 39108
rect 10918 39074 10938 39108
rect 10972 39074 11006 39108
rect 11044 39074 11060 39108
rect 11436 39074 11456 39108
rect 11490 39074 11524 39108
rect 11562 39074 11578 39108
rect 11838 39074 11858 39108
rect 11892 39074 11926 39108
rect 11964 39074 11980 39108
rect 12356 39074 12376 39108
rect 12410 39074 12444 39108
rect 12482 39074 12498 39108
rect 12758 39074 12778 39108
rect 12812 39074 12846 39108
rect 12884 39074 12900 39108
rect 13628 39108 13631 39147
rect 2220 37816 2225 37855
rect 2395 37816 2398 37855
rect 2220 37743 2225 37782
rect 2395 37743 2398 37782
rect 2220 37670 2225 37709
rect 2395 37670 2398 37709
rect 2220 37597 2225 37636
rect 2395 37597 2398 37636
rect 2220 37524 2225 37563
rect 2395 37524 2398 37563
rect 2220 37451 2225 37490
rect 2395 37451 2398 37490
rect 2220 37378 2225 37417
rect 2395 37378 2398 37417
rect 2220 37305 2225 37344
rect 2395 37305 2398 37344
rect 2220 37232 2225 37271
rect 2395 37232 2398 37271
rect 2220 37159 2225 37198
rect 2395 37159 2398 37198
rect 2220 37086 2225 37125
rect 2395 37086 2398 37125
rect 2220 37013 2225 37052
rect 2395 37013 2398 37052
rect 2877 39015 3087 39037
rect 13453 39036 13458 39075
rect 12969 39028 13175 39036
rect 3055 37541 3087 39015
rect 2877 37502 3087 37541
rect 2911 37468 2949 37502
rect 2983 37468 3021 37502
rect 3055 37468 3087 37502
rect 2877 37429 3087 37468
rect 2911 37395 2949 37429
rect 2983 37395 3021 37429
rect 3055 37395 3087 37429
rect 2877 37356 3087 37395
rect 2911 37322 2949 37356
rect 2983 37322 3021 37356
rect 3055 37322 3087 37356
rect 2877 37283 3087 37322
rect 2911 37249 2949 37283
rect 2983 37249 3021 37283
rect 3055 37249 3087 37283
rect 2877 37210 3087 37249
rect 2911 37176 2949 37210
rect 2983 37176 3021 37210
rect 3055 37176 3087 37210
rect 2877 37137 3087 37176
rect 2911 37103 2949 37137
rect 2983 37103 3021 37137
rect 3055 37103 3087 37137
rect 3797 37502 3975 37541
rect 3831 37468 3869 37502
rect 3903 37468 3941 37502
rect 3797 37429 3975 37468
rect 3831 37395 3869 37429
rect 3903 37395 3941 37429
rect 3797 37356 3975 37395
rect 3831 37322 3869 37356
rect 3903 37322 3941 37356
rect 3797 37283 3975 37322
rect 3831 37249 3869 37283
rect 3903 37249 3941 37283
rect 3797 37210 3975 37249
rect 3831 37176 3869 37210
rect 3903 37176 3941 37210
rect 3797 37137 3975 37176
rect 3831 37103 3869 37137
rect 3903 37103 3941 37137
rect 4751 38972 4789 39006
rect 4823 38972 4861 39006
rect 4717 38932 4895 38972
rect 4751 38898 4789 38932
rect 4823 38898 4861 38932
rect 4717 38858 4895 38898
rect 4751 38824 4789 38858
rect 4823 38824 4861 38858
rect 4717 38784 4895 38824
rect 4751 38750 4789 38784
rect 4823 38750 4861 38784
rect 4717 38710 4895 38750
rect 4751 38676 4789 38710
rect 4823 38676 4861 38710
rect 4717 38636 4895 38676
rect 4751 38602 4789 38636
rect 4823 38602 4861 38636
rect 4717 38562 4895 38602
rect 4751 38528 4789 38562
rect 4823 38528 4861 38562
rect 4717 38487 4895 38528
rect 4751 38453 4789 38487
rect 4823 38453 4861 38487
rect 4717 38412 4895 38453
rect 4751 38378 4789 38412
rect 4823 38378 4861 38412
rect 4717 38337 4895 38378
rect 4751 38303 4789 38337
rect 4823 38303 4861 38337
rect 4717 38262 4895 38303
rect 4751 38228 4789 38262
rect 4823 38228 4861 38262
rect 4717 38187 4895 38228
rect 4751 38153 4789 38187
rect 4823 38153 4861 38187
rect 4717 38112 4895 38153
rect 4751 38078 4789 38112
rect 4823 38078 4861 38112
rect 4717 38037 4895 38078
rect 4751 38003 4789 38037
rect 4823 38003 4861 38037
rect 4717 37962 4895 38003
rect 4751 37928 4789 37962
rect 4823 37928 4861 37962
rect 4717 37887 4895 37928
rect 4751 37853 4789 37887
rect 4823 37853 4861 37887
rect 4717 37812 4895 37853
rect 4751 37778 4789 37812
rect 4823 37778 4861 37812
rect 4717 37737 4895 37778
rect 4751 37703 4789 37737
rect 4823 37703 4861 37737
rect 4717 37662 4895 37703
rect 4751 37628 4789 37662
rect 4823 37628 4861 37662
rect 4717 37587 4895 37628
rect 4751 37553 4789 37587
rect 4823 37553 4861 37587
rect 4717 37512 4895 37553
rect 4751 37478 4789 37512
rect 4823 37478 4861 37512
rect 4717 37437 4895 37478
rect 4751 37403 4789 37437
rect 4823 37403 4861 37437
rect 4717 37362 4895 37403
rect 4751 37328 4789 37362
rect 4823 37328 4861 37362
rect 4717 37287 4895 37328
rect 4751 37253 4789 37287
rect 4823 37253 4861 37287
rect 4717 37212 4895 37253
rect 4751 37178 4789 37212
rect 4823 37178 4861 37212
rect 4717 37137 4895 37178
rect 4751 37103 4789 37137
rect 4823 37103 4861 37137
rect 5671 38972 5709 39006
rect 5743 38972 5781 39006
rect 5637 38932 5815 38972
rect 5671 38898 5709 38932
rect 5743 38898 5781 38932
rect 5637 38858 5815 38898
rect 5671 38824 5709 38858
rect 5743 38824 5781 38858
rect 5637 38784 5815 38824
rect 5671 38750 5709 38784
rect 5743 38750 5781 38784
rect 5637 38710 5815 38750
rect 5671 38676 5709 38710
rect 5743 38676 5781 38710
rect 5637 38636 5815 38676
rect 5671 38602 5709 38636
rect 5743 38602 5781 38636
rect 5637 38562 5815 38602
rect 5671 38528 5709 38562
rect 5743 38528 5781 38562
rect 5637 38487 5815 38528
rect 5671 38453 5709 38487
rect 5743 38453 5781 38487
rect 5637 38412 5815 38453
rect 5671 38378 5709 38412
rect 5743 38378 5781 38412
rect 5637 38337 5815 38378
rect 5671 38303 5709 38337
rect 5743 38303 5781 38337
rect 5637 38262 5815 38303
rect 5671 38228 5709 38262
rect 5743 38228 5781 38262
rect 5637 38187 5815 38228
rect 5671 38153 5709 38187
rect 5743 38153 5781 38187
rect 5637 38112 5815 38153
rect 5671 38078 5709 38112
rect 5743 38078 5781 38112
rect 5637 38037 5815 38078
rect 5671 38003 5709 38037
rect 5743 38003 5781 38037
rect 5637 37962 5815 38003
rect 5671 37928 5709 37962
rect 5743 37928 5781 37962
rect 5637 37887 5815 37928
rect 5671 37853 5709 37887
rect 5743 37853 5781 37887
rect 5637 37812 5815 37853
rect 5671 37778 5709 37812
rect 5743 37778 5781 37812
rect 5637 37737 5815 37778
rect 5671 37703 5709 37737
rect 5743 37703 5781 37737
rect 5637 37662 5815 37703
rect 5671 37628 5709 37662
rect 5743 37628 5781 37662
rect 5637 37587 5815 37628
rect 5671 37553 5709 37587
rect 5743 37553 5781 37587
rect 5637 37512 5815 37553
rect 5671 37478 5709 37512
rect 5743 37478 5781 37512
rect 5637 37437 5815 37478
rect 5671 37403 5709 37437
rect 5743 37403 5781 37437
rect 5637 37362 5815 37403
rect 5671 37328 5709 37362
rect 5743 37328 5781 37362
rect 5637 37287 5815 37328
rect 5671 37253 5709 37287
rect 5743 37253 5781 37287
rect 5637 37212 5815 37253
rect 5671 37178 5709 37212
rect 5743 37178 5781 37212
rect 5637 37137 5815 37178
rect 5671 37103 5709 37137
rect 5743 37103 5781 37137
rect 6591 38972 6629 39006
rect 6663 38972 6701 39006
rect 6557 38932 6735 38972
rect 6591 38898 6629 38932
rect 6663 38898 6701 38932
rect 6557 38858 6735 38898
rect 6591 38824 6629 38858
rect 6663 38824 6701 38858
rect 6557 38784 6735 38824
rect 6591 38750 6629 38784
rect 6663 38750 6701 38784
rect 6557 38710 6735 38750
rect 6591 38676 6629 38710
rect 6663 38676 6701 38710
rect 6557 38636 6735 38676
rect 6591 38602 6629 38636
rect 6663 38602 6701 38636
rect 6557 38562 6735 38602
rect 6591 38528 6629 38562
rect 6663 38528 6701 38562
rect 6557 38487 6735 38528
rect 6591 38453 6629 38487
rect 6663 38453 6701 38487
rect 6557 38412 6735 38453
rect 6591 38378 6629 38412
rect 6663 38378 6701 38412
rect 6557 38337 6735 38378
rect 6591 38303 6629 38337
rect 6663 38303 6701 38337
rect 6557 38262 6735 38303
rect 6591 38228 6629 38262
rect 6663 38228 6701 38262
rect 6557 38187 6735 38228
rect 6591 38153 6629 38187
rect 6663 38153 6701 38187
rect 6557 38112 6735 38153
rect 6591 38078 6629 38112
rect 6663 38078 6701 38112
rect 6557 38037 6735 38078
rect 6591 38003 6629 38037
rect 6663 38003 6701 38037
rect 6557 37962 6735 38003
rect 6591 37928 6629 37962
rect 6663 37928 6701 37962
rect 6557 37887 6735 37928
rect 6591 37853 6629 37887
rect 6663 37853 6701 37887
rect 6557 37812 6735 37853
rect 6591 37778 6629 37812
rect 6663 37778 6701 37812
rect 6557 37737 6735 37778
rect 6591 37703 6629 37737
rect 6663 37703 6701 37737
rect 6557 37662 6735 37703
rect 6591 37628 6629 37662
rect 6663 37628 6701 37662
rect 6557 37587 6735 37628
rect 6591 37553 6629 37587
rect 6663 37553 6701 37587
rect 6557 37512 6735 37553
rect 6591 37478 6629 37512
rect 6663 37478 6701 37512
rect 6557 37437 6735 37478
rect 6591 37403 6629 37437
rect 6663 37403 6701 37437
rect 6557 37362 6735 37403
rect 6591 37328 6629 37362
rect 6663 37328 6701 37362
rect 6557 37287 6735 37328
rect 6591 37253 6629 37287
rect 6663 37253 6701 37287
rect 6557 37212 6735 37253
rect 6591 37178 6629 37212
rect 6663 37178 6701 37212
rect 6557 37137 6735 37178
rect 6591 37103 6629 37137
rect 6663 37103 6701 37137
rect 7511 38972 7549 39006
rect 7583 38972 7621 39006
rect 7477 38932 7655 38972
rect 7511 38898 7549 38932
rect 7583 38898 7621 38932
rect 7477 38858 7655 38898
rect 7511 38824 7549 38858
rect 7583 38824 7621 38858
rect 7477 38784 7655 38824
rect 7511 38750 7549 38784
rect 7583 38750 7621 38784
rect 7477 38710 7655 38750
rect 7511 38676 7549 38710
rect 7583 38676 7621 38710
rect 7477 38636 7655 38676
rect 7511 38602 7549 38636
rect 7583 38602 7621 38636
rect 7477 38562 7655 38602
rect 7511 38528 7549 38562
rect 7583 38528 7621 38562
rect 7477 38487 7655 38528
rect 7511 38453 7549 38487
rect 7583 38453 7621 38487
rect 7477 38412 7655 38453
rect 7511 38378 7549 38412
rect 7583 38378 7621 38412
rect 7477 38337 7655 38378
rect 7511 38303 7549 38337
rect 7583 38303 7621 38337
rect 7477 38262 7655 38303
rect 7511 38228 7549 38262
rect 7583 38228 7621 38262
rect 7477 38187 7655 38228
rect 7511 38153 7549 38187
rect 7583 38153 7621 38187
rect 7477 38112 7655 38153
rect 7511 38078 7549 38112
rect 7583 38078 7621 38112
rect 7477 38037 7655 38078
rect 7511 38003 7549 38037
rect 7583 38003 7621 38037
rect 7477 37962 7655 38003
rect 7511 37928 7549 37962
rect 7583 37928 7621 37962
rect 7477 37887 7655 37928
rect 7511 37853 7549 37887
rect 7583 37853 7621 37887
rect 7477 37812 7655 37853
rect 7511 37778 7549 37812
rect 7583 37778 7621 37812
rect 7477 37737 7655 37778
rect 7511 37703 7549 37737
rect 7583 37703 7621 37737
rect 7477 37662 7655 37703
rect 7511 37628 7549 37662
rect 7583 37628 7621 37662
rect 7477 37587 7655 37628
rect 7511 37553 7549 37587
rect 7583 37553 7621 37587
rect 7477 37512 7655 37553
rect 7511 37478 7549 37512
rect 7583 37478 7621 37512
rect 7477 37437 7655 37478
rect 7511 37403 7549 37437
rect 7583 37403 7621 37437
rect 7477 37362 7655 37403
rect 7511 37328 7549 37362
rect 7583 37328 7621 37362
rect 7477 37287 7655 37328
rect 7511 37253 7549 37287
rect 7583 37253 7621 37287
rect 7477 37212 7655 37253
rect 7511 37178 7549 37212
rect 7583 37178 7621 37212
rect 7477 37137 7655 37178
rect 7511 37103 7549 37137
rect 7583 37103 7621 37137
rect 8431 38972 8469 39006
rect 8503 38972 8541 39006
rect 8397 38932 8575 38972
rect 8431 38898 8469 38932
rect 8503 38898 8541 38932
rect 8397 38858 8575 38898
rect 8431 38824 8469 38858
rect 8503 38824 8541 38858
rect 8397 38784 8575 38824
rect 8431 38750 8469 38784
rect 8503 38750 8541 38784
rect 8397 38710 8575 38750
rect 8431 38676 8469 38710
rect 8503 38676 8541 38710
rect 8397 38636 8575 38676
rect 8431 38602 8469 38636
rect 8503 38602 8541 38636
rect 8397 38562 8575 38602
rect 8431 38528 8469 38562
rect 8503 38528 8541 38562
rect 8397 38487 8575 38528
rect 8431 38453 8469 38487
rect 8503 38453 8541 38487
rect 8397 38412 8575 38453
rect 8431 38378 8469 38412
rect 8503 38378 8541 38412
rect 8397 38337 8575 38378
rect 8431 38303 8469 38337
rect 8503 38303 8541 38337
rect 8397 38262 8575 38303
rect 8431 38228 8469 38262
rect 8503 38228 8541 38262
rect 8397 38187 8575 38228
rect 8431 38153 8469 38187
rect 8503 38153 8541 38187
rect 8397 38112 8575 38153
rect 8431 38078 8469 38112
rect 8503 38078 8541 38112
rect 8397 38037 8575 38078
rect 8431 38003 8469 38037
rect 8503 38003 8541 38037
rect 8397 37962 8575 38003
rect 8431 37928 8469 37962
rect 8503 37928 8541 37962
rect 8397 37887 8575 37928
rect 8431 37853 8469 37887
rect 8503 37853 8541 37887
rect 8397 37812 8575 37853
rect 8431 37778 8469 37812
rect 8503 37778 8541 37812
rect 8397 37737 8575 37778
rect 8431 37703 8469 37737
rect 8503 37703 8541 37737
rect 8397 37662 8575 37703
rect 8431 37628 8469 37662
rect 8503 37628 8541 37662
rect 8397 37587 8575 37628
rect 8431 37553 8469 37587
rect 8503 37553 8541 37587
rect 8397 37512 8575 37553
rect 8431 37478 8469 37512
rect 8503 37478 8541 37512
rect 8397 37437 8575 37478
rect 8431 37403 8469 37437
rect 8503 37403 8541 37437
rect 8397 37362 8575 37403
rect 8431 37328 8469 37362
rect 8503 37328 8541 37362
rect 8397 37287 8575 37328
rect 8431 37253 8469 37287
rect 8503 37253 8541 37287
rect 8397 37212 8575 37253
rect 8431 37178 8469 37212
rect 8503 37178 8541 37212
rect 8397 37137 8575 37178
rect 8431 37103 8469 37137
rect 8503 37103 8541 37137
rect 9351 38972 9389 39006
rect 9423 38972 9461 39006
rect 9317 38932 9495 38972
rect 9351 38898 9389 38932
rect 9423 38898 9461 38932
rect 9317 38858 9495 38898
rect 9351 38824 9389 38858
rect 9423 38824 9461 38858
rect 9317 38784 9495 38824
rect 9351 38750 9389 38784
rect 9423 38750 9461 38784
rect 9317 38710 9495 38750
rect 9351 38676 9389 38710
rect 9423 38676 9461 38710
rect 9317 38636 9495 38676
rect 9351 38602 9389 38636
rect 9423 38602 9461 38636
rect 9317 38562 9495 38602
rect 9351 38528 9389 38562
rect 9423 38528 9461 38562
rect 9317 38487 9495 38528
rect 9351 38453 9389 38487
rect 9423 38453 9461 38487
rect 9317 38412 9495 38453
rect 9351 38378 9389 38412
rect 9423 38378 9461 38412
rect 9317 38337 9495 38378
rect 9351 38303 9389 38337
rect 9423 38303 9461 38337
rect 9317 38262 9495 38303
rect 9351 38228 9389 38262
rect 9423 38228 9461 38262
rect 9317 38187 9495 38228
rect 9351 38153 9389 38187
rect 9423 38153 9461 38187
rect 9317 38112 9495 38153
rect 9351 38078 9389 38112
rect 9423 38078 9461 38112
rect 9317 38037 9495 38078
rect 9351 38003 9389 38037
rect 9423 38003 9461 38037
rect 9317 37962 9495 38003
rect 9351 37928 9389 37962
rect 9423 37928 9461 37962
rect 9317 37887 9495 37928
rect 9351 37853 9389 37887
rect 9423 37853 9461 37887
rect 9317 37812 9495 37853
rect 9351 37778 9389 37812
rect 9423 37778 9461 37812
rect 9317 37737 9495 37778
rect 9351 37703 9389 37737
rect 9423 37703 9461 37737
rect 9317 37662 9495 37703
rect 9351 37628 9389 37662
rect 9423 37628 9461 37662
rect 9317 37587 9495 37628
rect 9351 37553 9389 37587
rect 9423 37553 9461 37587
rect 9317 37512 9495 37553
rect 9351 37478 9389 37512
rect 9423 37478 9461 37512
rect 9317 37437 9495 37478
rect 9351 37403 9389 37437
rect 9423 37403 9461 37437
rect 9317 37362 9495 37403
rect 9351 37328 9389 37362
rect 9423 37328 9461 37362
rect 9317 37287 9495 37328
rect 9351 37253 9389 37287
rect 9423 37253 9461 37287
rect 9317 37212 9495 37253
rect 9351 37178 9389 37212
rect 9423 37178 9461 37212
rect 9317 37137 9495 37178
rect 9351 37103 9389 37137
rect 9423 37103 9461 37137
rect 10271 38972 10309 39006
rect 10343 38972 10381 39006
rect 10237 38932 10415 38972
rect 10271 38898 10309 38932
rect 10343 38898 10381 38932
rect 10237 38858 10415 38898
rect 10271 38824 10309 38858
rect 10343 38824 10381 38858
rect 10237 38784 10415 38824
rect 10271 38750 10309 38784
rect 10343 38750 10381 38784
rect 10237 38710 10415 38750
rect 10271 38676 10309 38710
rect 10343 38676 10381 38710
rect 10237 38636 10415 38676
rect 10271 38602 10309 38636
rect 10343 38602 10381 38636
rect 10237 38562 10415 38602
rect 10271 38528 10309 38562
rect 10343 38528 10381 38562
rect 10237 38487 10415 38528
rect 10271 38453 10309 38487
rect 10343 38453 10381 38487
rect 10237 38412 10415 38453
rect 10271 38378 10309 38412
rect 10343 38378 10381 38412
rect 10237 38337 10415 38378
rect 10271 38303 10309 38337
rect 10343 38303 10381 38337
rect 10237 38262 10415 38303
rect 10271 38228 10309 38262
rect 10343 38228 10381 38262
rect 10237 38187 10415 38228
rect 10271 38153 10309 38187
rect 10343 38153 10381 38187
rect 10237 38112 10415 38153
rect 10271 38078 10309 38112
rect 10343 38078 10381 38112
rect 10237 38037 10415 38078
rect 10271 38003 10309 38037
rect 10343 38003 10381 38037
rect 10237 37962 10415 38003
rect 10271 37928 10309 37962
rect 10343 37928 10381 37962
rect 10237 37887 10415 37928
rect 10271 37853 10309 37887
rect 10343 37853 10381 37887
rect 10237 37812 10415 37853
rect 10271 37778 10309 37812
rect 10343 37778 10381 37812
rect 10237 37737 10415 37778
rect 10271 37703 10309 37737
rect 10343 37703 10381 37737
rect 10237 37662 10415 37703
rect 10271 37628 10309 37662
rect 10343 37628 10381 37662
rect 10237 37587 10415 37628
rect 10271 37553 10309 37587
rect 10343 37553 10381 37587
rect 10237 37512 10415 37553
rect 10271 37478 10309 37512
rect 10343 37478 10381 37512
rect 10237 37437 10415 37478
rect 10271 37403 10309 37437
rect 10343 37403 10381 37437
rect 10237 37362 10415 37403
rect 10271 37328 10309 37362
rect 10343 37328 10381 37362
rect 10237 37287 10415 37328
rect 10271 37253 10309 37287
rect 10343 37253 10381 37287
rect 10237 37212 10415 37253
rect 10271 37178 10309 37212
rect 10343 37178 10381 37212
rect 10237 37137 10415 37178
rect 10271 37103 10309 37137
rect 10343 37103 10381 37137
rect 11157 38451 11335 38490
rect 11191 38417 11229 38451
rect 11263 38417 11301 38451
rect 11157 38378 11335 38417
rect 11191 38344 11229 38378
rect 11263 38344 11301 38378
rect 11157 38305 11335 38344
rect 11191 38271 11229 38305
rect 11263 38271 11301 38305
rect 11157 38232 11335 38271
rect 11191 38198 11229 38232
rect 11263 38198 11301 38232
rect 11157 38159 11335 38198
rect 11191 38125 11229 38159
rect 11263 38125 11301 38159
rect 11157 38086 11335 38125
rect 11191 38052 11229 38086
rect 11263 38052 11301 38086
rect 11157 38013 11335 38052
rect 11191 37979 11229 38013
rect 11263 37979 11301 38013
rect 11157 37940 11335 37979
rect 11191 37906 11229 37940
rect 11263 37906 11301 37940
rect 11157 37867 11335 37906
rect 11191 37833 11229 37867
rect 11263 37833 11301 37867
rect 11157 37794 11335 37833
rect 11191 37760 11229 37794
rect 11263 37760 11301 37794
rect 11157 37721 11335 37760
rect 11191 37687 11229 37721
rect 11263 37687 11301 37721
rect 11157 37648 11335 37687
rect 11191 37614 11229 37648
rect 11263 37614 11301 37648
rect 11157 37575 11335 37614
rect 11191 37541 11229 37575
rect 11263 37541 11301 37575
rect 11157 37502 11335 37541
rect 11191 37468 11229 37502
rect 11263 37468 11301 37502
rect 11157 37429 11335 37468
rect 11191 37395 11229 37429
rect 11263 37395 11301 37429
rect 11157 37356 11335 37395
rect 11191 37322 11229 37356
rect 11263 37322 11301 37356
rect 11157 37283 11335 37322
rect 11191 37249 11229 37283
rect 11263 37249 11301 37283
rect 11157 37210 11335 37249
rect 11191 37176 11229 37210
rect 11263 37176 11301 37210
rect 11157 37137 11335 37176
rect 11191 37103 11229 37137
rect 11263 37103 11301 37137
rect 12077 38451 12255 38490
rect 12111 38417 12149 38451
rect 12183 38417 12221 38451
rect 12077 38378 12255 38417
rect 12111 38344 12149 38378
rect 12183 38344 12221 38378
rect 12077 38305 12255 38344
rect 12111 38271 12149 38305
rect 12183 38271 12221 38305
rect 12077 38232 12255 38271
rect 12111 38198 12149 38232
rect 12183 38198 12221 38232
rect 12077 38159 12255 38198
rect 12111 38125 12149 38159
rect 12183 38125 12221 38159
rect 12077 38086 12255 38125
rect 12111 38052 12149 38086
rect 12183 38052 12221 38086
rect 12077 38013 12255 38052
rect 12111 37979 12149 38013
rect 12183 37979 12221 38013
rect 12077 37940 12255 37979
rect 12111 37906 12149 37940
rect 12183 37906 12221 37940
rect 12077 37867 12255 37906
rect 12111 37833 12149 37867
rect 12183 37833 12221 37867
rect 12077 37794 12255 37833
rect 12111 37760 12149 37794
rect 12183 37760 12221 37794
rect 12077 37721 12255 37760
rect 12111 37687 12149 37721
rect 12183 37687 12221 37721
rect 12077 37648 12255 37687
rect 12111 37614 12149 37648
rect 12183 37614 12221 37648
rect 12077 37575 12255 37614
rect 12111 37541 12149 37575
rect 12183 37541 12221 37575
rect 12077 37502 12255 37541
rect 12111 37468 12149 37502
rect 12183 37468 12221 37502
rect 12077 37429 12255 37468
rect 12111 37395 12149 37429
rect 12183 37395 12221 37429
rect 12077 37356 12255 37395
rect 12111 37322 12149 37356
rect 12183 37322 12221 37356
rect 12077 37283 12255 37322
rect 12111 37249 12149 37283
rect 12183 37249 12221 37283
rect 12077 37210 12255 37249
rect 12111 37176 12149 37210
rect 12183 37176 12221 37210
rect 12077 37137 12255 37176
rect 12111 37103 12149 37137
rect 12183 37103 12221 37137
rect 12969 38490 12997 39028
rect 12969 38451 13175 38490
rect 12969 38417 12997 38451
rect 13031 38417 13069 38451
rect 13103 38417 13141 38451
rect 12969 38378 13175 38417
rect 12969 38344 12997 38378
rect 13031 38344 13069 38378
rect 13103 38344 13141 38378
rect 12969 38305 13175 38344
rect 12969 38271 12997 38305
rect 13031 38271 13069 38305
rect 13103 38271 13141 38305
rect 12969 38232 13175 38271
rect 12969 38198 12997 38232
rect 13031 38198 13069 38232
rect 13103 38198 13141 38232
rect 12969 38159 13175 38198
rect 12969 38125 12997 38159
rect 13031 38125 13069 38159
rect 13103 38125 13141 38159
rect 12969 38086 13175 38125
rect 12969 38052 12997 38086
rect 13031 38052 13069 38086
rect 13103 38052 13141 38086
rect 12969 38013 13175 38052
rect 12969 37979 12997 38013
rect 13031 37979 13069 38013
rect 13103 37979 13141 38013
rect 12969 37940 13175 37979
rect 12969 37906 12997 37940
rect 13031 37906 13069 37940
rect 13103 37906 13141 37940
rect 12969 37867 13175 37906
rect 12969 37833 12997 37867
rect 13031 37833 13069 37867
rect 13103 37833 13141 37867
rect 12969 37794 13175 37833
rect 12969 37760 12997 37794
rect 13031 37760 13069 37794
rect 13103 37760 13141 37794
rect 12969 37721 13175 37760
rect 12969 37687 12997 37721
rect 13031 37687 13069 37721
rect 13103 37687 13141 37721
rect 12969 37648 13175 37687
rect 12969 37614 12997 37648
rect 13031 37614 13069 37648
rect 13103 37614 13141 37648
rect 12969 37575 13175 37614
rect 12969 37541 12997 37575
rect 13031 37541 13069 37575
rect 13103 37541 13141 37575
rect 12969 37502 13175 37541
rect 12969 37468 12997 37502
rect 13031 37468 13069 37502
rect 13103 37468 13141 37502
rect 12969 37429 13175 37468
rect 12969 37395 12997 37429
rect 13031 37395 13069 37429
rect 13103 37395 13141 37429
rect 12969 37356 13175 37395
rect 12969 37322 12997 37356
rect 13031 37322 13069 37356
rect 13103 37322 13141 37356
rect 12969 37283 13175 37322
rect 12969 37249 12997 37283
rect 13031 37249 13069 37283
rect 13103 37249 13141 37283
rect 12969 37210 13175 37249
rect 12969 37176 12997 37210
rect 13031 37176 13069 37210
rect 13103 37176 13141 37210
rect 12969 37137 13175 37176
rect 12969 37103 12997 37137
rect 13031 37103 13069 37137
rect 13103 37103 13141 37137
rect 2877 37032 3087 37103
rect 12969 37032 13175 37103
rect 13628 39035 13631 39074
rect 13453 38963 13458 39002
rect 13628 38962 13631 39001
rect 13453 38890 13458 38929
rect 13628 38889 13631 38928
rect 13453 38817 13458 38856
rect 13628 38816 13631 38855
rect 13453 38744 13458 38783
rect 13628 38743 13631 38782
rect 13453 38671 13458 38710
rect 13628 38670 13631 38709
rect 13453 38598 13458 38637
rect 13628 38597 13631 38636
rect 13453 38525 13458 38564
rect 13628 38524 13631 38563
rect 13453 38452 13458 38491
rect 13628 38451 13631 38490
rect 13453 38379 13458 38418
rect 13628 38378 13631 38417
rect 13453 38306 13458 38345
rect 13628 38305 13631 38344
rect 13453 38233 13458 38272
rect 13628 38232 13631 38271
rect 13453 38160 13458 38199
rect 13628 38159 13631 38198
rect 13453 38087 13458 38126
rect 13628 38086 13631 38125
rect 13453 38014 13458 38053
rect 13628 38013 13631 38052
rect 13453 37941 13458 37980
rect 13628 37940 13631 37979
rect 13453 37868 13458 37907
rect 13628 37867 13631 37906
rect 13453 37795 13458 37834
rect 13628 37794 13631 37833
rect 13453 37722 13458 37761
rect 13628 37721 13631 37760
rect 13453 37649 13458 37688
rect 13628 37648 13631 37687
rect 13453 37576 13458 37615
rect 13628 37575 13631 37614
rect 13453 37503 13458 37542
rect 13628 37502 13631 37541
rect 13453 37430 13458 37469
rect 13628 37429 13631 37468
rect 13453 37357 13458 37396
rect 13628 37356 13631 37395
rect 13453 37284 13458 37323
rect 13628 37283 13631 37322
rect 13453 37211 13458 37250
rect 13628 37210 13631 37249
rect 13453 37138 13458 37177
rect 13628 37137 13631 37176
rect 13453 37065 13458 37104
rect 13628 37064 13631 37103
rect 2220 36940 2225 36979
rect 2395 36940 2398 36979
rect 2220 36867 2225 36906
rect 2395 36867 2398 36906
rect 2220 36794 2225 36833
rect 2395 36794 2398 36833
rect 2220 36721 2225 36760
rect 2395 36721 2398 36760
rect 2220 36648 2225 36687
rect 2395 36648 2398 36687
rect 2220 36575 2225 36614
rect 2395 36575 2398 36614
rect 2220 36502 2225 36541
rect 2395 36502 2398 36541
rect 2566 36986 3176 36998
rect 2566 36952 2583 36986
rect 2617 36964 3176 36986
rect 3210 36964 3244 36998
rect 3278 36964 3578 36998
rect 3612 36964 3646 36998
rect 3680 36964 4096 36998
rect 4130 36964 4164 36998
rect 4198 36964 4498 36998
rect 4532 36964 4566 36998
rect 4600 36964 5016 36998
rect 5050 36964 5084 36998
rect 5118 36964 5418 36998
rect 5452 36964 5486 36998
rect 5520 36964 5936 36998
rect 5970 36964 6004 36998
rect 6038 36964 6338 36998
rect 6372 36964 6406 36998
rect 6440 36964 6856 36998
rect 6890 36964 6924 36998
rect 6958 36964 7258 36998
rect 7292 36964 7326 36998
rect 7360 36964 7776 36998
rect 7810 36964 7844 36998
rect 7878 36964 8178 36998
rect 8212 36964 8246 36998
rect 8280 36964 8696 36998
rect 8730 36964 8764 36998
rect 8798 36964 9098 36998
rect 9132 36964 9166 36998
rect 9200 36964 9616 36998
rect 9650 36964 9684 36998
rect 9718 36964 10018 36998
rect 10052 36964 10086 36998
rect 10120 36964 10536 36998
rect 10570 36964 10604 36998
rect 10638 36964 10938 36998
rect 10972 36964 11006 36998
rect 11040 36964 11456 36998
rect 11490 36964 11524 36998
rect 11558 36964 11858 36998
rect 11892 36964 11926 36998
rect 11960 36964 12376 36998
rect 12410 36964 12444 36998
rect 12478 36964 12778 36998
rect 12812 36964 12846 36998
rect 12880 36964 13337 36998
rect 2617 36952 13337 36964
rect 2566 36901 13337 36952
rect 2566 36867 2583 36901
rect 2617 36867 13337 36901
rect 2566 36816 13337 36867
rect 2566 36782 2583 36816
rect 2617 36782 13337 36816
rect 2566 36731 13337 36782
rect 2566 36697 2583 36731
rect 2617 36697 13337 36731
rect 2566 36646 13337 36697
rect 2566 36612 2583 36646
rect 2617 36612 13337 36646
rect 2566 36560 13337 36612
rect 2566 36526 2583 36560
rect 2617 36526 13337 36560
rect 2566 36514 13337 36526
rect 3156 36508 13337 36514
rect 3156 36474 3176 36508
rect 3210 36474 3244 36508
rect 3278 36474 3578 36508
rect 3612 36474 3646 36508
rect 3680 36474 4096 36508
rect 4130 36474 4164 36508
rect 4198 36474 4498 36508
rect 4532 36474 4566 36508
rect 4600 36474 5016 36508
rect 5050 36474 5084 36508
rect 5118 36474 5418 36508
rect 5452 36474 5486 36508
rect 5520 36474 5936 36508
rect 5970 36474 6004 36508
rect 6038 36474 6338 36508
rect 6372 36474 6406 36508
rect 6440 36474 6856 36508
rect 6890 36474 6924 36508
rect 6958 36474 7258 36508
rect 7292 36474 7326 36508
rect 7360 36474 7776 36508
rect 7810 36474 7844 36508
rect 7878 36474 8178 36508
rect 8212 36474 8246 36508
rect 8280 36474 8696 36508
rect 8730 36474 8764 36508
rect 8798 36474 9098 36508
rect 9132 36474 9166 36508
rect 9200 36474 9616 36508
rect 9650 36474 9684 36508
rect 9718 36474 10018 36508
rect 10052 36474 10086 36508
rect 10120 36474 10536 36508
rect 10570 36474 10604 36508
rect 10638 36474 10938 36508
rect 10972 36474 11006 36508
rect 11040 36474 11456 36508
rect 11490 36474 11524 36508
rect 11558 36474 11858 36508
rect 11892 36474 11926 36508
rect 11960 36474 12376 36508
rect 12410 36474 12444 36508
rect 12478 36474 12778 36508
rect 12812 36474 12846 36508
rect 12880 36474 13337 36508
rect 3156 36468 13337 36474
rect 13453 36992 13458 37031
rect 13628 36991 13631 37030
rect 13453 36919 13458 36958
rect 13628 36918 13631 36957
rect 13453 36846 13458 36885
rect 13628 36845 13631 36884
rect 13453 36773 13458 36812
rect 13628 36772 13631 36811
rect 13453 36700 13458 36739
rect 13628 36699 13631 36738
rect 13453 36627 13458 36666
rect 13628 36626 13631 36665
rect 13453 36554 13458 36593
rect 13628 36553 13631 36592
rect 13453 36481 13458 36520
rect 2220 36429 2225 36468
rect 2395 36429 2398 36468
rect 2220 36356 2225 36395
rect 2395 36356 2398 36395
rect 13628 36480 13631 36519
rect 13453 36408 13458 36447
rect 2220 36283 2225 36322
rect 2395 36283 2398 36322
rect 2220 36210 2225 36249
rect 2395 36210 2398 36249
rect 2220 36137 2225 36176
rect 2395 36137 2398 36176
rect 2220 36064 2225 36103
rect 2395 36064 2398 36103
rect 2220 35991 2225 36030
rect 2395 35991 2398 36030
rect 2220 35918 2225 35957
rect 2395 35918 2398 35957
rect 2220 35845 2225 35884
rect 2395 35845 2398 35884
rect 2220 35772 2225 35811
rect 2395 35772 2398 35811
rect 2220 35699 2225 35738
rect 2395 35699 2398 35738
rect 2220 35626 2225 35665
rect 2395 35626 2398 35665
rect 2220 35553 2225 35592
rect 2395 35553 2398 35592
rect 2220 35480 2225 35519
rect 2395 35480 2398 35519
rect 2220 35407 2225 35446
rect 2395 35407 2398 35446
rect 2220 35334 2225 35373
rect 2395 35334 2398 35373
rect 2220 35261 2225 35300
rect 2395 35261 2398 35300
rect 2220 35188 2225 35227
rect 2395 35188 2398 35227
rect 2220 35115 2225 35154
rect 2395 35115 2398 35154
rect 2220 35042 2225 35081
rect 2395 35042 2398 35081
rect 2220 34969 2225 35008
rect 2395 34969 2398 35008
rect 2220 34896 2225 34935
rect 2395 34896 2398 34935
rect 2220 34823 2225 34862
rect 2395 34823 2398 34862
rect 2220 34750 2225 34789
rect 2395 34750 2398 34789
rect 2220 34677 2225 34716
rect 2395 34677 2398 34716
rect 2220 34604 2225 34643
rect 2395 34604 2398 34643
rect 2220 34531 2225 34570
rect 2395 34531 2398 34570
rect 2220 34458 2225 34497
rect 2395 34458 2398 34497
rect 2220 34385 2225 34424
rect 2395 34385 2398 34424
rect 2220 34312 2225 34351
rect 2395 34312 2398 34351
rect 2220 34239 2225 34278
rect 2395 34239 2398 34278
rect 2877 36362 3083 36386
rect 2877 36328 2943 36362
rect 2977 36328 3021 36362
rect 3055 36328 3083 36362
rect 2877 36290 3083 36328
rect 2877 36256 2943 36290
rect 2977 36256 3021 36290
rect 3055 36256 3083 36290
rect 2877 36218 3083 36256
rect 2877 36184 2943 36218
rect 2977 36184 3021 36218
rect 3055 36184 3083 36218
rect 2877 36146 3083 36184
rect 2877 36112 2943 36146
rect 2977 36112 3021 36146
rect 3055 36112 3083 36146
rect 2877 36074 3083 36112
rect 2877 36040 2943 36074
rect 2977 36040 3021 36074
rect 3055 36040 3083 36074
rect 2877 36002 3083 36040
rect 2877 35968 2943 36002
rect 2977 35968 3021 36002
rect 3055 35968 3083 36002
rect 2877 35930 3083 35968
rect 2877 35896 2943 35930
rect 2977 35896 3021 35930
rect 3055 35896 3083 35930
rect 2877 35858 3083 35896
rect 2877 35824 2943 35858
rect 2977 35824 3021 35858
rect 3055 35824 3083 35858
rect 2877 35786 3083 35824
rect 2877 35752 2943 35786
rect 2977 35752 3021 35786
rect 3055 35752 3083 35786
rect 2877 35714 3083 35752
rect 2877 35680 2943 35714
rect 2977 35680 3021 35714
rect 3055 35680 3083 35714
rect 2877 35642 3083 35680
rect 2877 35608 2943 35642
rect 2977 35608 3021 35642
rect 3055 35608 3083 35642
rect 2877 35570 3083 35608
rect 2877 35536 2943 35570
rect 2977 35536 3021 35570
rect 3055 35536 3083 35570
rect 2877 35498 3083 35536
rect 2877 35464 2943 35498
rect 2977 35464 3021 35498
rect 3055 35464 3083 35498
rect 2877 35426 3083 35464
rect 2877 35392 2943 35426
rect 2977 35392 3021 35426
rect 3055 35392 3083 35426
rect 2877 35354 3083 35392
rect 2877 35320 2943 35354
rect 2977 35320 3021 35354
rect 3055 35320 3083 35354
rect 2877 35282 3083 35320
rect 2877 35248 2943 35282
rect 2977 35248 3021 35282
rect 3055 35248 3083 35282
rect 2877 35210 3083 35248
rect 2877 35176 2943 35210
rect 2977 35176 3021 35210
rect 3055 35176 3083 35210
rect 2877 35138 3083 35176
rect 2877 35104 2943 35138
rect 2977 35104 3021 35138
rect 3055 35104 3083 35138
rect 2877 35066 3083 35104
rect 2877 35032 2943 35066
rect 2977 35032 3021 35066
rect 3055 35032 3083 35066
rect 2877 34994 3083 35032
rect 2877 34960 2943 34994
rect 2977 34960 3021 34994
rect 3055 34960 3083 34994
rect 2877 34922 3083 34960
rect 2877 34888 2943 34922
rect 2977 34888 3021 34922
rect 3055 34888 3083 34922
rect 2877 34850 3083 34888
rect 2877 34816 2943 34850
rect 2977 34816 3021 34850
rect 3055 34816 3083 34850
rect 2877 34778 3083 34816
rect 2877 34744 2943 34778
rect 2977 34744 3021 34778
rect 3055 34744 3083 34778
rect 2877 34706 3083 34744
rect 2877 34672 2943 34706
rect 2977 34672 3021 34706
rect 3055 34672 3083 34706
rect 2877 34634 3083 34672
rect 2877 34600 2943 34634
rect 2977 34600 3021 34634
rect 3055 34600 3083 34634
rect 2877 34562 3083 34600
rect 2877 34528 2943 34562
rect 2977 34528 3021 34562
rect 3055 34528 3083 34562
rect 2877 34490 3083 34528
rect 2877 34456 2943 34490
rect 2977 34456 3021 34490
rect 3055 34456 3083 34490
rect 2877 34418 3083 34456
rect 2877 34384 2943 34418
rect 2977 34384 3021 34418
rect 3055 34384 3083 34418
rect 2877 34346 3083 34384
rect 2877 34312 2943 34346
rect 2977 34312 3021 34346
rect 3055 34312 3083 34346
rect 2877 34274 3083 34312
rect 2877 34240 2943 34274
rect 2977 34240 3021 34274
rect 3055 34240 3083 34274
rect 1736 34110 1808 34144
rect 1702 34069 1834 34110
rect 1736 34035 1808 34069
rect 1702 33994 1834 34035
rect 1736 33960 1808 33994
rect 1702 33919 1834 33960
rect 1736 33885 1808 33919
rect 1702 33844 1834 33885
rect 1736 33810 1808 33844
rect 1702 33769 1834 33810
rect 1736 33735 1808 33769
rect 1702 33694 1834 33735
rect 1736 33660 1808 33694
rect 1702 33619 1834 33660
rect 1736 33585 1808 33619
rect 1702 33544 1834 33585
rect 1736 33510 1808 33544
rect 1702 33469 1834 33510
rect 1736 33435 1808 33469
rect 1702 33394 1834 33435
rect 1736 33360 1808 33394
rect 1702 33319 1834 33360
rect 1736 33285 1808 33319
rect 1702 33244 1834 33285
rect 1736 33210 1808 33244
rect 1702 33169 1834 33210
rect 1736 33135 1808 33169
rect 1702 33094 1834 33135
rect 1736 33060 1808 33094
rect 1702 33019 1834 33060
rect 1736 32985 1808 33019
rect 1702 32944 1834 32985
rect 1736 32910 1808 32944
rect 1702 32869 1834 32910
rect 1736 32835 1808 32869
rect 1702 32793 1834 32835
rect 1736 32759 1808 32793
rect 1702 32717 1834 32759
rect 1736 32683 1808 32717
rect 1702 32641 1834 32683
rect 1736 32607 1808 32641
rect 1702 32565 1834 32607
rect 1736 32531 1808 32565
rect 2188 34069 2225 34103
rect 2154 34030 2225 34069
rect 2188 33996 2225 34030
rect 2154 33957 2225 33996
rect 2188 33923 2225 33957
rect 2154 33884 2225 33923
rect 2188 33850 2225 33884
rect 2154 33811 2225 33850
rect 2188 33777 2225 33811
rect 2154 33738 2225 33777
rect 2188 33704 2225 33738
rect 2154 33665 2225 33704
rect 2188 33631 2225 33665
rect 2154 33592 2225 33631
rect 2188 33558 2225 33592
rect 2154 33519 2225 33558
rect 2188 33485 2225 33519
rect 2154 33446 2225 33485
rect 2188 33412 2225 33446
rect 2154 33373 2225 33412
rect 2188 33339 2225 33373
rect 2154 33300 2225 33339
rect 2188 33266 2225 33300
rect 2154 33227 2225 33266
rect 2188 33193 2225 33227
rect 2154 33154 2225 33193
rect 2188 33120 2225 33154
rect 2154 33081 2225 33120
rect 2188 33047 2225 33081
rect 2154 33008 2225 33047
rect 2188 32974 2225 33008
rect 2154 32935 2225 32974
rect 2188 32901 2225 32935
rect 2154 32861 2225 32901
rect 2188 32827 2225 32861
rect 2154 32787 2225 32827
rect 2188 32753 2225 32787
rect 2154 32713 2225 32753
rect 2188 32679 2225 32713
rect 2154 32639 2225 32679
rect 2188 32605 2225 32639
rect 2154 32565 2225 32605
rect 2188 32531 2225 32565
rect 2877 34202 3083 34240
rect 2877 34168 2943 34202
rect 2977 34168 3021 34202
rect 3055 34168 3083 34202
rect 2877 34130 3083 34168
rect 2877 34096 2943 34130
rect 2977 34096 3021 34130
rect 3055 34096 3083 34130
rect 2877 34058 3083 34096
rect 2877 34024 2943 34058
rect 2977 34024 3021 34058
rect 3055 34024 3083 34058
rect 2877 33986 3083 34024
rect 2877 33952 2943 33986
rect 2977 33952 3021 33986
rect 3055 33952 3083 33986
rect 2877 33914 3083 33952
rect 2877 33880 2943 33914
rect 2977 33880 3021 33914
rect 3055 33880 3083 33914
rect 2877 33842 3083 33880
rect 2877 33808 2943 33842
rect 2977 33808 3021 33842
rect 3055 33808 3083 33842
rect 2877 33770 3083 33808
rect 2877 33736 2943 33770
rect 2977 33736 3021 33770
rect 3055 33736 3083 33770
rect 2877 33698 3083 33736
rect 2877 33664 2943 33698
rect 2977 33664 3021 33698
rect 3055 33664 3083 33698
rect 2877 33626 3083 33664
rect 2877 33592 2943 33626
rect 2977 33592 3021 33626
rect 3055 33592 3083 33626
rect 2877 33554 3083 33592
rect 2877 33520 2943 33554
rect 2977 33520 3021 33554
rect 3055 33520 3083 33554
rect 2877 33482 3083 33520
rect 2877 33448 2943 33482
rect 2977 33448 3021 33482
rect 3055 33448 3083 33482
rect 2877 33410 3083 33448
rect 2877 33376 2943 33410
rect 2977 33376 3021 33410
rect 3055 33376 3083 33410
rect 2877 33338 3083 33376
rect 2877 33304 2943 33338
rect 2977 33304 3021 33338
rect 3055 33304 3083 33338
rect 2877 33266 3083 33304
rect 2877 33232 2943 33266
rect 2977 33232 3021 33266
rect 3055 33232 3083 33266
rect 2877 33194 3083 33232
rect 2877 33160 2943 33194
rect 2977 33160 3021 33194
rect 3055 33160 3083 33194
rect 2877 33121 3083 33160
rect 2877 33087 2943 33121
rect 2977 33087 3021 33121
rect 3055 33087 3083 33121
rect 2877 33048 3083 33087
rect 2877 33014 2943 33048
rect 2977 33014 3021 33048
rect 3055 33014 3083 33048
rect 2877 32975 3083 33014
rect 2877 32941 2943 32975
rect 2977 32941 3021 32975
rect 3055 32941 3083 32975
rect 2877 32902 3083 32941
rect 2877 32868 2943 32902
rect 2977 32868 3021 32902
rect 3055 32868 3083 32902
rect 2877 32829 3083 32868
rect 2877 32795 2943 32829
rect 2977 32795 3021 32829
rect 3055 32795 3083 32829
rect 2877 32756 3083 32795
rect 2877 32722 2943 32756
rect 2977 32722 3021 32756
rect 3055 32722 3083 32756
rect 2877 32683 3083 32722
rect 2877 32649 2943 32683
rect 2977 32649 3021 32683
rect 3055 32649 3083 32683
rect 2877 32610 3083 32649
rect 2877 32576 2943 32610
rect 2977 32576 3021 32610
rect 3055 32576 3083 32610
rect 2877 32537 3083 32576
rect 2877 32503 2943 32537
rect 2977 32503 3021 32537
rect 3055 32503 3083 32537
rect 12969 36353 13175 36386
rect 3797 33121 3975 33160
rect 3831 33087 3869 33121
rect 3903 33087 3941 33121
rect 3797 33048 3975 33087
rect 3831 33014 3869 33048
rect 3903 33014 3941 33048
rect 3797 32975 3975 33014
rect 3831 32941 3869 32975
rect 3903 32941 3941 32975
rect 3797 32902 3975 32941
rect 3831 32868 3869 32902
rect 3903 32868 3941 32902
rect 3797 32829 3975 32868
rect 3831 32795 3869 32829
rect 3903 32795 3941 32829
rect 3797 32756 3975 32795
rect 3831 32722 3869 32756
rect 3903 32722 3941 32756
rect 3797 32683 3975 32722
rect 3831 32649 3869 32683
rect 3903 32649 3941 32683
rect 3797 32610 3975 32649
rect 3831 32576 3869 32610
rect 3903 32576 3941 32610
rect 3797 32537 3975 32576
rect 3831 32503 3869 32537
rect 3903 32503 3941 32537
rect 12969 32503 12997 36353
rect 13628 36407 13631 36446
rect 13453 36335 13458 36374
rect 13628 36334 13631 36373
rect 13453 36262 13458 36301
rect 13628 36261 13631 36300
rect 13453 36189 13458 36228
rect 13628 36188 13631 36227
rect 13453 36116 13458 36155
rect 13628 36115 13631 36154
rect 13453 36043 13458 36082
rect 13628 36042 13631 36081
rect 13453 35970 13458 36009
rect 13628 35969 13631 36008
rect 13453 35897 13458 35936
rect 13628 35896 13631 35935
rect 13453 35824 13458 35863
rect 13775 39504 13781 39543
rect 14019 39575 14025 39614
rect 13775 39431 13781 39470
rect 14019 39502 14025 39541
rect 13775 39358 13781 39397
rect 14019 39429 14025 39468
rect 13775 39285 13781 39324
rect 14019 39356 14025 39395
rect 13775 39212 13781 39251
rect 14019 39283 14025 39322
rect 13775 39139 13781 39178
rect 14019 39210 14025 39249
rect 13775 39066 13781 39105
rect 14019 39137 14025 39176
rect 13775 38993 13781 39032
rect 14019 39064 14025 39103
rect 13775 38920 13781 38959
rect 14019 38991 14025 39030
rect 13775 38847 13781 38886
rect 14019 38918 14025 38957
rect 13775 38774 13781 38813
rect 14019 38845 14025 38884
rect 13775 38701 13781 38740
rect 14019 38772 14025 38811
rect 13775 38628 13781 38667
rect 14019 38699 14025 38738
rect 13775 38555 13781 38594
rect 14019 38626 14025 38665
rect 13775 38482 13781 38521
rect 14019 38553 14025 38592
rect 13775 38409 13781 38448
rect 14019 38480 14025 38519
rect 13775 38336 13781 38375
rect 14019 38407 14025 38446
rect 13775 38263 13781 38302
rect 14019 38334 14025 38373
rect 13775 38190 13781 38229
rect 14019 38261 14025 38300
rect 13775 38117 13781 38156
rect 14019 38188 14025 38227
rect 13775 38044 13781 38083
rect 14019 38115 14025 38154
rect 13775 37971 13781 38010
rect 14019 38042 14025 38081
rect 13775 37898 13781 37937
rect 14019 37969 14025 38008
rect 13775 37825 13781 37864
rect 14019 37896 14025 37935
rect 13775 37752 13781 37791
rect 14019 37823 14025 37862
rect 13775 37679 13781 37718
rect 14019 37750 14025 37789
rect 13775 37606 13781 37645
rect 14019 37677 14025 37716
rect 13775 37533 13781 37572
rect 14019 37604 14025 37643
rect 13775 37460 13781 37499
rect 14019 37531 14025 37570
rect 13775 37387 13781 37426
rect 14019 37458 14025 37497
rect 13775 37314 13781 37353
rect 14019 37385 14025 37424
rect 13775 37241 13781 37280
rect 14019 37312 14025 37351
rect 13775 37168 13781 37207
rect 14019 37239 14025 37278
rect 13775 37095 13781 37134
rect 14019 37166 14025 37205
rect 13775 37022 13781 37061
rect 14019 37093 14025 37132
rect 13775 36949 13781 36988
rect 14019 37020 14025 37059
rect 13775 36876 13781 36915
rect 14019 36947 14025 36986
rect 13775 36803 13781 36842
rect 14019 36874 14025 36913
rect 13775 36730 13781 36769
rect 14019 36801 14025 36840
rect 13775 36657 13781 36696
rect 14019 36728 14025 36767
rect 13775 36584 13781 36623
rect 14019 36655 14025 36694
rect 13775 36511 13781 36550
rect 14019 36582 14025 36621
rect 13775 36438 13781 36477
rect 14019 36509 14025 36548
rect 13775 36365 13781 36404
rect 14019 36436 14025 36475
rect 13775 36292 13781 36331
rect 14019 36363 14025 36402
rect 13775 36219 13781 36258
rect 14019 36290 14025 36329
rect 13775 36146 13781 36185
rect 14019 36217 14025 36256
rect 13775 36073 13781 36112
rect 14019 36144 14025 36183
rect 13775 36000 13781 36039
rect 14019 36071 14025 36110
rect 13775 35927 13781 35966
rect 14019 35998 14025 36037
rect 13775 35854 13781 35893
rect 14019 35925 14025 35964
rect 13775 35781 13781 35820
rect 14019 35852 14025 35891
rect 13775 35708 13781 35747
rect 14019 35779 14025 35818
rect 13775 35635 13781 35674
rect 14019 35706 14025 35745
rect 13775 35562 13781 35601
rect 14019 35633 14025 35672
rect 13775 35489 13781 35528
rect 14019 35560 14025 35599
rect 13775 35416 13781 35455
rect 14019 35487 14025 35526
rect 13775 35343 13781 35382
rect 14019 35414 14025 35453
rect 13775 35270 13781 35309
rect 14019 35341 14025 35380
rect 13775 35197 13781 35236
rect 14019 35268 14025 35307
rect 13775 35124 13781 35163
rect 14019 35195 14025 35234
rect 13775 35051 13781 35090
rect 14019 35122 14025 35161
rect 13775 34978 13781 35017
rect 2877 32432 3083 32503
rect 12969 32432 13175 32503
rect 13628 33046 13631 33084
rect 13628 32974 13631 33012
rect 13628 32902 13631 32940
rect 13628 32830 13631 32868
rect 13628 32758 13631 32796
rect 13628 32686 13631 32724
rect 13628 32614 13631 32652
rect 13628 32542 13631 32580
rect 13628 32470 13631 32508
rect 13628 32398 13631 32436
rect 2480 32364 3176 32398
rect 3210 32364 3244 32398
rect 3278 32364 3578 32398
rect 3612 32364 3646 32398
rect 3680 32364 4096 32398
rect 4130 32364 4164 32398
rect 4198 32364 4498 32398
rect 4532 32364 4566 32398
rect 4600 32364 5016 32398
rect 5050 32364 5084 32398
rect 5118 32364 5418 32398
rect 5452 32364 5486 32398
rect 5520 32364 5936 32398
rect 5970 32364 6004 32398
rect 6038 32364 6338 32398
rect 6372 32364 6406 32398
rect 6440 32364 6856 32398
rect 6890 32364 6924 32398
rect 6958 32364 7258 32398
rect 7292 32364 7326 32398
rect 7360 32364 7776 32398
rect 7810 32364 7844 32398
rect 7878 32364 8178 32398
rect 8212 32364 8246 32398
rect 8280 32364 8696 32398
rect 8730 32364 8764 32398
rect 8798 32364 9098 32398
rect 9132 32364 9166 32398
rect 9200 32364 9616 32398
rect 9650 32364 9684 32398
rect 9718 32364 10018 32398
rect 10052 32364 10086 32398
rect 10120 32364 10536 32398
rect 10570 32364 10604 32398
rect 10638 32364 10938 32398
rect 10972 32364 11006 32398
rect 11040 32364 11456 32398
rect 11490 32364 11524 32398
rect 11558 32364 11858 32398
rect 11892 32364 11926 32398
rect 11960 32364 12376 32398
rect 12410 32364 12444 32398
rect 12478 32364 12778 32398
rect 12812 32364 12846 32398
rect 12880 32364 12900 32398
rect 2480 32210 12900 32364
rect 2480 32176 2494 32210
rect 2528 32176 2579 32210
rect 2613 32176 2664 32210
rect 2698 32176 12900 32210
rect 2480 32138 12900 32176
rect 2480 32104 2494 32138
rect 2528 32104 2579 32138
rect 2613 32104 2664 32138
rect 2698 32104 12900 32138
rect 2480 31911 12900 32104
rect 3156 31908 12900 31911
rect 3156 31874 3176 31908
rect 3210 31874 3244 31908
rect 3278 31874 3578 31908
rect 3612 31874 3646 31908
rect 3680 31874 4096 31908
rect 4130 31874 4164 31908
rect 4198 31874 4498 31908
rect 4532 31874 4566 31908
rect 4600 31874 5016 31908
rect 5050 31874 5084 31908
rect 5118 31874 5418 31908
rect 5452 31874 5486 31908
rect 5520 31874 5936 31908
rect 5970 31874 6004 31908
rect 6038 31874 6338 31908
rect 6372 31874 6406 31908
rect 6440 31874 6856 31908
rect 6890 31874 6924 31908
rect 6958 31874 7258 31908
rect 7292 31874 7326 31908
rect 7360 31874 7776 31908
rect 7810 31874 7844 31908
rect 7878 31874 8178 31908
rect 8212 31874 8246 31908
rect 8280 31874 8696 31908
rect 8730 31874 8764 31908
rect 8798 31874 9098 31908
rect 9132 31874 9166 31908
rect 9200 31874 9616 31908
rect 9650 31874 9684 31908
rect 9718 31874 10018 31908
rect 10052 31874 10086 31908
rect 10120 31874 10536 31908
rect 10570 31874 10604 31908
rect 10638 31874 10938 31908
rect 10972 31874 11006 31908
rect 11040 31874 11456 31908
rect 11490 31874 11524 31908
rect 11558 31874 11858 31908
rect 11892 31874 11926 31908
rect 11960 31874 12376 31908
rect 12410 31874 12444 31908
rect 12478 31874 12778 31908
rect 12812 31874 12846 31908
rect 12880 31874 12900 31908
rect 3156 31868 12900 31874
rect 13628 32326 13631 32364
rect 13628 32254 13631 32292
rect 13628 32182 13631 32220
rect 13628 32110 13631 32148
rect 13628 32038 13631 32076
rect 13628 31966 13631 32004
rect 13628 31894 13631 31932
rect 13628 31822 13631 31860
rect 2395 30342 2420 30381
rect 2395 30269 2420 30308
rect 2395 30196 2420 30235
rect 2395 30123 2420 30162
rect 2395 30050 2420 30089
rect 2395 29977 2420 30016
rect 2395 29904 2420 29943
rect 2395 29831 2420 29870
rect 2395 29758 2420 29797
rect 2395 29685 2420 29724
rect 2395 29612 2420 29651
rect 2395 29539 2420 29578
rect 2395 29466 2420 29505
rect 2395 29393 2420 29432
rect 2395 29320 2420 29359
rect 2395 29247 2420 29286
rect 2395 29174 2420 29213
rect 2395 29101 2420 29140
rect 2395 29028 2420 29067
rect 2395 28955 2420 28994
rect 2395 28882 2420 28921
rect 2395 28809 2420 28848
rect 2395 28736 2420 28775
rect 2395 28663 2420 28702
rect 2395 28590 2420 28629
rect 2395 28517 2420 28556
rect 2395 28444 2420 28483
rect 2395 28371 2420 28410
rect 2395 28298 2420 28337
rect 2395 28225 2420 28264
rect 2395 28152 2420 28191
rect 2395 28079 2420 28118
rect 2395 28006 2420 28045
rect 2395 27933 2420 27972
rect 2395 27860 2420 27899
rect 2877 31762 3083 31786
rect 3055 28560 3083 31762
rect 2877 28521 3083 28560
rect 2911 28487 2949 28521
rect 2983 28487 3021 28521
rect 3055 28487 3083 28521
rect 2877 28448 3083 28487
rect 2911 28414 2949 28448
rect 2983 28414 3021 28448
rect 3055 28414 3083 28448
rect 2877 28375 3083 28414
rect 2911 28341 2949 28375
rect 2983 28341 3021 28375
rect 3055 28341 3083 28375
rect 2877 28302 3083 28341
rect 2911 28268 2949 28302
rect 2983 28268 3021 28302
rect 3055 28268 3083 28302
rect 2877 28229 3083 28268
rect 2911 28195 2949 28229
rect 2983 28195 3021 28229
rect 3055 28195 3083 28229
rect 2877 28156 3083 28195
rect 2911 28122 2949 28156
rect 2983 28122 3021 28156
rect 3055 28122 3083 28156
rect 2877 28083 3083 28122
rect 2911 28049 2949 28083
rect 2983 28049 3021 28083
rect 3055 28049 3083 28083
rect 2877 28010 3083 28049
rect 2911 27976 2949 28010
rect 2983 27976 3021 28010
rect 3055 27976 3083 28010
rect 2877 27937 3083 27976
rect 2911 27903 2949 27937
rect 2983 27903 3021 27937
rect 3055 27903 3083 27937
rect 12969 31753 13175 31786
rect 3797 28521 3975 28560
rect 3831 28487 3869 28521
rect 3903 28487 3941 28521
rect 3797 28448 3975 28487
rect 3831 28414 3869 28448
rect 3903 28414 3941 28448
rect 3797 28375 3975 28414
rect 3831 28341 3869 28375
rect 3903 28341 3941 28375
rect 3797 28302 3975 28341
rect 3831 28268 3869 28302
rect 3903 28268 3941 28302
rect 3797 28229 3975 28268
rect 3831 28195 3869 28229
rect 3903 28195 3941 28229
rect 3797 28156 3975 28195
rect 3831 28122 3869 28156
rect 3903 28122 3941 28156
rect 3797 28083 3975 28122
rect 3831 28049 3869 28083
rect 3903 28049 3941 28083
rect 3797 28010 3975 28049
rect 3831 27976 3869 28010
rect 3903 27976 3941 28010
rect 3797 27937 3975 27976
rect 3831 27903 3869 27937
rect 3903 27903 3941 27937
rect 12969 27903 12997 31753
rect 2877 27832 3083 27903
rect 12969 27832 13175 27903
rect 13628 31750 13631 31788
rect 13628 31678 13631 31716
rect 13628 31606 13631 31644
rect 13628 31534 13631 31572
rect 13628 31462 13631 31500
rect 13628 31390 13631 31428
rect 13628 31318 13631 31356
rect 13628 31246 13631 31284
rect 13628 31174 13631 31212
rect 13628 31102 13631 31140
rect 13628 31030 13631 31068
rect 13628 30958 13631 30996
rect 13628 30886 13631 30924
rect 13628 30814 13631 30852
rect 13628 30742 13631 30780
rect 13628 30670 13631 30708
rect 13628 30598 13631 30636
rect 13628 30526 13631 30564
rect 13628 30454 13631 30492
rect 13628 30382 13631 30420
rect 13628 30310 13631 30348
rect 13628 30238 13631 30276
rect 13628 30166 13631 30204
rect 13628 30094 13631 30132
rect 13628 30022 13631 30060
rect 13628 29950 13631 29988
rect 13628 29878 13631 29916
rect 13628 29806 13631 29844
rect 13628 29734 13631 29772
rect 13628 29662 13631 29700
rect 13628 29590 13631 29628
rect 13628 29518 13631 29556
rect 13628 29446 13631 29484
rect 13628 29374 13631 29412
rect 13628 29302 13631 29340
rect 13628 29230 13631 29268
rect 13628 29158 13631 29196
rect 13628 29086 13631 29124
rect 13628 29014 13631 29052
rect 13628 28942 13631 28980
rect 13628 28870 13631 28908
rect 13628 28798 13631 28836
rect 13628 28726 13631 28764
rect 13628 28654 13631 28692
rect 13628 28582 13631 28620
rect 13628 28510 13631 28548
rect 13628 28438 13631 28476
rect 13628 28366 13631 28404
rect 13628 28294 13631 28332
rect 13628 28222 13631 28260
rect 13628 28150 13631 28188
rect 13628 28078 13631 28116
rect 13628 28006 13631 28044
rect 13628 27934 13631 27972
rect 13628 27862 13631 27900
rect 2395 27787 2420 27826
rect 2395 27714 2420 27753
rect 2395 27641 2420 27680
rect 2395 27568 2420 27607
rect 2395 27495 2420 27534
rect 2395 27422 2420 27461
rect 2395 27349 2420 27388
rect 2395 27276 2420 27315
rect 3156 27764 3176 27798
rect 3210 27764 3244 27798
rect 3278 27764 3578 27798
rect 3612 27764 3646 27798
rect 3680 27764 4096 27798
rect 4130 27764 4164 27798
rect 4198 27764 4498 27798
rect 4532 27764 4566 27798
rect 4600 27764 5016 27798
rect 5050 27764 5084 27798
rect 5118 27764 5418 27798
rect 5452 27764 5486 27798
rect 5520 27764 5936 27798
rect 5970 27764 6004 27798
rect 6038 27764 6338 27798
rect 6372 27764 6406 27798
rect 6440 27764 6856 27798
rect 6890 27764 6924 27798
rect 6958 27764 7258 27798
rect 7292 27764 7326 27798
rect 7360 27764 7776 27798
rect 7810 27764 7844 27798
rect 7878 27764 8178 27798
rect 8212 27764 8246 27798
rect 8280 27764 8696 27798
rect 8730 27764 8764 27798
rect 8798 27764 9098 27798
rect 9132 27764 9166 27798
rect 9200 27764 9616 27798
rect 9650 27764 9684 27798
rect 9718 27764 10018 27798
rect 10052 27764 10086 27798
rect 10120 27764 10536 27798
rect 10570 27764 10604 27798
rect 10638 27764 10938 27798
rect 10972 27764 11006 27798
rect 11040 27764 11456 27798
rect 11490 27764 11524 27798
rect 11558 27764 11858 27798
rect 11892 27764 11926 27798
rect 11960 27764 12376 27798
rect 12410 27764 12444 27798
rect 12478 27764 12778 27798
rect 12812 27764 12846 27798
rect 12880 27764 12900 27798
rect 3156 27574 12900 27764
rect 3156 27540 3170 27574
rect 3204 27540 3245 27574
rect 3279 27540 3320 27574
rect 3354 27540 12900 27574
rect 3156 27308 12900 27540
rect 4996 27274 5016 27308
rect 5050 27274 5084 27308
rect 5118 27274 5418 27308
rect 5452 27274 5486 27308
rect 5520 27274 5936 27308
rect 5970 27274 6004 27308
rect 6038 27274 6338 27308
rect 6372 27274 6406 27308
rect 6440 27274 6856 27308
rect 6890 27274 6924 27308
rect 6958 27274 7258 27308
rect 7292 27274 7326 27308
rect 7360 27274 7776 27308
rect 7810 27274 7844 27308
rect 7878 27274 8178 27308
rect 8212 27274 8246 27308
rect 8280 27274 8696 27308
rect 8730 27274 8764 27308
rect 8798 27274 9098 27308
rect 9132 27274 9166 27308
rect 9200 27274 9616 27308
rect 9650 27274 9684 27308
rect 9718 27274 10018 27308
rect 10052 27274 10086 27308
rect 10120 27274 10536 27308
rect 10570 27274 10604 27308
rect 10638 27274 10938 27308
rect 10972 27274 11006 27308
rect 11040 27274 11456 27308
rect 11490 27274 11524 27308
rect 11558 27274 11858 27308
rect 11892 27274 11926 27308
rect 11960 27274 12376 27308
rect 12410 27274 12444 27308
rect 12478 27274 12778 27308
rect 12812 27274 12846 27308
rect 12880 27274 12900 27308
rect 5134 27268 12900 27274
rect 13628 27790 13631 27828
rect 13628 27718 13631 27756
rect 13628 27646 13631 27684
rect 13628 27574 13631 27612
rect 13628 27502 13631 27540
rect 13628 27430 13631 27468
rect 13628 27358 13631 27396
rect 13628 27286 13631 27324
rect 2348 27242 2386 27268
rect 2327 27233 2420 27242
rect 2327 27203 2361 27233
rect 4367 27231 4401 27233
rect 2225 27169 2314 27200
rect 2348 27169 2361 27203
rect 4397 27199 4401 27231
rect 4435 27199 4532 27233
rect 4397 27197 4532 27199
rect 2225 27166 2361 27169
rect 2259 27165 2361 27166
rect 4367 27165 4532 27197
rect 13628 27214 13631 27252
rect 2259 27132 2293 27165
rect 2225 27063 2293 27132
rect 4367 27131 4430 27165
rect 4299 27123 4430 27131
rect 4320 27097 4363 27123
rect 4397 27097 4430 27123
rect 4320 27089 4362 27097
rect 4299 27063 4362 27089
rect 2004 26911 2072 26979
rect 1936 26893 1946 26911
rect 1980 26908 2072 26911
rect 1980 26893 2038 26908
rect 1936 26854 2038 26893
rect 1936 26843 1946 26854
rect 1834 26820 1946 26843
rect 1980 26840 2038 26854
rect 4044 26874 4078 26908
rect 4112 26874 4198 26908
rect 4044 26840 4198 26874
rect 1834 26809 1840 26820
rect 1874 26786 1970 26820
rect 4044 26806 4096 26840
rect 1868 26781 1970 26786
rect 1868 26775 1946 26781
rect 1834 26772 1946 26775
rect 1834 26747 1902 26772
rect 3976 26772 4096 26806
rect 3976 26769 4028 26772
rect 1834 26713 1840 26747
rect 1874 26713 1902 26747
rect 3908 26735 3947 26738
rect 3981 26735 4028 26769
rect 1834 26670 1902 26713
rect 3908 26704 4028 26735
rect 3908 26670 3960 26704
rect 1840 26641 1914 26670
rect 1948 26641 1988 26670
rect 2022 26641 2062 26670
rect 2096 26641 2136 26670
rect 2170 26641 2210 26670
rect 2244 26641 2284 26670
rect 2318 26641 2358 26670
rect 2392 26641 2432 26670
rect 2466 26641 2506 26670
rect 2540 26641 2580 26670
rect 2614 26641 2654 26670
rect 2688 26641 2729 26670
rect 2763 26641 2804 26670
rect 3567 26663 3960 26670
rect 3601 26629 3653 26663
rect 3687 26629 3739 26663
rect 3773 26629 3826 26663
rect 3860 26629 3913 26663
rect 3947 26629 3960 26663
rect 3913 26591 3960 26629
rect 3947 26557 3960 26591
rect 3913 26519 3960 26557
rect 3947 26485 3960 26519
rect 3913 26447 3960 26485
rect 3947 26413 3960 26447
rect 3913 26375 3960 26413
rect 3947 26341 3960 26375
rect 3913 26303 3960 26341
rect 3947 26269 3960 26303
rect 3913 26231 3960 26269
rect 3947 26197 3960 26231
rect 3913 26159 3960 26197
rect 3947 26125 3960 26159
rect 3913 26087 3960 26125
rect 3947 26053 3960 26087
rect 3913 26015 3960 26053
rect 3947 25981 3960 26015
rect 3913 25943 3960 25981
rect 3947 25909 3960 25943
rect 3913 25871 3960 25909
rect 3947 25837 3960 25871
rect 3913 25799 3960 25837
rect 3947 25765 3960 25799
rect 3913 25727 3960 25765
rect 3947 25693 3960 25727
rect 3913 25655 3960 25693
rect 3947 25621 3960 25655
rect 3913 25583 3960 25621
rect 3947 25549 3960 25583
rect 3913 25511 3960 25549
rect 3947 25477 3960 25511
rect 3913 25439 3960 25477
rect 3947 25405 3960 25439
rect 3913 25367 3960 25405
rect 3947 25333 3960 25367
rect 3913 25295 3960 25333
rect 3947 25261 3960 25295
rect 3913 25223 3960 25261
rect 3947 25189 3960 25223
rect 3913 25151 3960 25189
rect 3947 25117 3960 25151
rect 3913 25079 3960 25117
rect 3947 25045 3960 25079
rect 3913 25007 3960 25045
rect 3947 24973 3960 25007
rect 3913 24935 3960 24973
rect 3947 24901 3960 24935
rect 3913 24863 3960 24901
rect 3947 24829 3960 24863
rect 3913 24791 3960 24829
rect 3947 24757 3960 24791
rect 3913 24719 3960 24757
rect 3947 24685 3960 24719
rect 3913 24647 3960 24685
rect 3947 24613 3960 24647
rect 3913 24575 3960 24613
rect 3947 24541 3960 24575
rect 3913 24503 3960 24541
rect 3947 24469 3960 24503
rect 3913 24431 3960 24469
rect 3947 24397 3960 24431
rect 3913 24359 3960 24397
rect 3947 24325 3960 24359
rect 3913 24287 3960 24325
rect 3947 24253 3960 24287
rect 3913 24215 3960 24253
rect 3947 24181 3960 24215
rect 3913 24143 3960 24181
rect 3947 24109 3960 24143
rect 3913 24071 3960 24109
rect 3947 24037 3960 24071
rect 3913 23999 3960 24037
rect 3947 23965 3960 23999
rect 3913 23927 3960 23965
rect 3947 23893 3960 23927
rect 3913 23855 3960 23893
rect 3947 23821 3960 23855
rect 3913 23783 3960 23821
rect 3947 23749 3960 23783
rect 3913 23711 3960 23749
rect 3947 23677 3960 23711
rect 3913 23639 3960 23677
rect 3947 23605 3960 23639
rect 3913 23567 3960 23605
rect 3947 23533 3960 23567
rect 3913 23495 3960 23533
rect 3947 23461 3960 23495
rect 3913 23423 3960 23461
rect 3947 23389 3960 23423
rect 3913 23351 3960 23389
rect 3947 23317 3960 23351
rect 3913 23279 3960 23317
rect 3947 23245 3960 23279
rect 3913 23207 3960 23245
rect 3947 23173 3960 23207
rect 3913 23135 3960 23173
rect 3947 23101 3960 23135
rect 3913 23063 3960 23101
rect 3947 23029 3960 23063
rect 3913 22991 3960 23029
rect 3947 22957 3960 22991
rect 3913 22919 3960 22957
rect 3947 22885 3960 22919
rect 3913 22847 3960 22885
rect 3947 22813 3960 22847
rect 3913 22775 3960 22813
rect 3947 22741 3960 22775
rect 3913 22703 3960 22741
rect 3947 22669 3960 22703
rect 3913 22631 3960 22669
rect 3947 22597 3960 22631
rect 3913 22559 3960 22597
rect 3947 22525 3960 22559
rect 3913 22487 3960 22525
rect 3947 22453 3960 22487
rect 3913 22415 3960 22453
rect 3947 22381 3960 22415
rect 3913 22343 3960 22381
rect 3947 22309 3960 22343
rect 3913 22271 3960 22309
rect 3947 22237 3960 22271
rect 3913 22199 3960 22237
rect 3947 22165 3960 22199
rect 3913 22127 3960 22165
rect 3947 22093 3960 22127
rect 3913 22055 3960 22093
rect 3947 22021 3960 22055
rect 3913 21983 3960 22021
rect 3947 21949 3960 21983
rect 3913 21911 3960 21949
rect 3947 21877 3960 21911
rect 3913 21839 3960 21877
rect 3947 21805 3960 21839
rect 3913 21767 3960 21805
rect 3947 21733 3960 21767
rect 3913 21695 3960 21733
rect 3947 21661 3960 21695
rect 3913 21623 3960 21661
rect 3947 21589 3960 21623
rect 3913 21551 3960 21589
rect 3947 21517 3960 21551
rect 3913 21479 3960 21517
rect 3947 21445 3960 21479
rect 3913 21407 3960 21445
rect 3947 21373 3960 21407
rect 3913 21335 3960 21373
rect 3947 21301 3960 21335
rect 3913 21263 3960 21301
rect 3947 21229 3960 21263
rect 3913 21191 3960 21229
rect 3947 21157 3960 21191
rect 3913 21119 3960 21157
rect 3947 21085 3960 21119
rect 3913 21047 3960 21085
rect 3947 21013 3960 21047
rect 3913 20975 3960 21013
rect 3947 20941 3960 20975
rect 3913 20903 3960 20941
rect 3947 20869 3960 20903
rect 3913 20831 3960 20869
rect 3947 20797 3960 20831
rect 3913 20759 3960 20797
rect 3947 20725 3960 20759
rect 3913 20687 3960 20725
rect 3947 20653 3960 20687
rect 3913 20615 3960 20653
rect 3947 20581 3960 20615
rect 3913 20543 3960 20581
rect 3947 20509 3960 20543
rect 3913 20471 3960 20509
rect 3947 20437 3960 20471
rect 3913 20399 3960 20437
rect 3947 20365 3960 20399
rect 3913 20327 3960 20365
rect 3947 20293 3960 20327
rect 3913 20255 3960 20293
rect 3947 20221 3960 20255
rect 3913 20183 3960 20221
rect 3947 20149 3960 20183
rect 3913 20111 3960 20149
rect 3947 20077 3960 20111
rect 3913 20039 3960 20077
rect 3947 20005 3960 20039
rect 3913 19967 3960 20005
rect 3947 19933 3960 19967
rect 3913 19895 3960 19933
rect 3947 19861 3960 19895
rect 3913 19823 3960 19861
rect 3947 19789 3960 19823
rect 3913 19751 3960 19789
rect 3947 19717 3960 19751
rect 3913 19679 3960 19717
rect 3947 19645 3960 19679
rect 3913 19607 3960 19645
rect 3947 19573 3960 19607
rect 3913 19534 3960 19573
rect 3947 19500 3960 19534
rect 4717 27162 4923 27186
rect 4717 27128 4783 27162
rect 4817 27128 4861 27162
rect 4895 27128 4923 27162
rect 4717 27089 4923 27128
rect 4717 27055 4783 27089
rect 4817 27055 4861 27089
rect 4895 27055 4923 27089
rect 4717 27016 4923 27055
rect 4717 26982 4783 27016
rect 4817 26982 4861 27016
rect 4895 26982 4923 27016
rect 4717 26943 4923 26982
rect 4717 26909 4783 26943
rect 4817 26909 4861 26943
rect 4895 26909 4923 26943
rect 4717 26870 4923 26909
rect 4717 26836 4783 26870
rect 4817 26836 4861 26870
rect 4895 26836 4923 26870
rect 4717 26797 4923 26836
rect 4717 26763 4783 26797
rect 4817 26763 4861 26797
rect 4895 26763 4923 26797
rect 4717 26724 4923 26763
rect 4717 26690 4783 26724
rect 4817 26690 4861 26724
rect 4895 26690 4923 26724
rect 4717 26651 4923 26690
rect 4717 26617 4783 26651
rect 4817 26617 4861 26651
rect 4895 26617 4923 26651
rect 4717 26578 4923 26617
rect 4717 26544 4783 26578
rect 4817 26544 4861 26578
rect 4895 26544 4923 26578
rect 4717 26505 4923 26544
rect 4717 26471 4783 26505
rect 4817 26471 4861 26505
rect 4895 26471 4923 26505
rect 4717 26432 4923 26471
rect 4717 26398 4783 26432
rect 4817 26398 4861 26432
rect 4895 26398 4923 26432
rect 4717 26359 4923 26398
rect 4717 26325 4783 26359
rect 4817 26325 4861 26359
rect 4895 26325 4923 26359
rect 4717 26286 4923 26325
rect 4717 26252 4783 26286
rect 4817 26252 4861 26286
rect 4895 26252 4923 26286
rect 4717 26213 4923 26252
rect 4717 26179 4783 26213
rect 4817 26179 4861 26213
rect 4895 26179 4923 26213
rect 4717 26140 4923 26179
rect 4717 26106 4783 26140
rect 4817 26106 4861 26140
rect 4895 26106 4923 26140
rect 4717 26067 4923 26106
rect 4717 26033 4783 26067
rect 4817 26033 4861 26067
rect 4895 26033 4923 26067
rect 4717 25994 4923 26033
rect 4717 25960 4783 25994
rect 4817 25960 4861 25994
rect 4895 25960 4923 25994
rect 4717 25921 4923 25960
rect 4717 25887 4783 25921
rect 4817 25887 4861 25921
rect 4895 25887 4923 25921
rect 4717 25848 4923 25887
rect 4717 25814 4783 25848
rect 4817 25814 4861 25848
rect 4895 25814 4923 25848
rect 4717 25775 4923 25814
rect 4717 25741 4783 25775
rect 4817 25741 4861 25775
rect 4895 25741 4923 25775
rect 4717 25702 4923 25741
rect 4717 25668 4783 25702
rect 4817 25668 4861 25702
rect 4895 25668 4923 25702
rect 4717 25629 4923 25668
rect 4717 25595 4783 25629
rect 4817 25595 4861 25629
rect 4895 25595 4923 25629
rect 4717 25556 4923 25595
rect 4717 25522 4783 25556
rect 4817 25522 4861 25556
rect 4895 25522 4923 25556
rect 4717 25483 4923 25522
rect 4717 25449 4783 25483
rect 4817 25449 4861 25483
rect 4895 25449 4923 25483
rect 4717 25410 4923 25449
rect 4717 25376 4783 25410
rect 4817 25376 4861 25410
rect 4895 25376 4923 25410
rect 4717 25337 4923 25376
rect 4717 25303 4783 25337
rect 4817 25303 4861 25337
rect 4895 25303 4923 25337
rect 4717 25264 4923 25303
rect 4717 25230 4783 25264
rect 4817 25230 4861 25264
rect 4895 25230 4923 25264
rect 4717 25191 4923 25230
rect 4717 25157 4783 25191
rect 4817 25157 4861 25191
rect 4895 25157 4923 25191
rect 4717 25118 4923 25157
rect 4717 25084 4783 25118
rect 4817 25084 4861 25118
rect 4895 25084 4923 25118
rect 4717 25045 4923 25084
rect 4717 25011 4783 25045
rect 4817 25011 4861 25045
rect 4895 25011 4923 25045
rect 4717 24972 4923 25011
rect 4717 24938 4783 24972
rect 4817 24938 4861 24972
rect 4895 24938 4923 24972
rect 4717 24899 4923 24938
rect 4717 24865 4783 24899
rect 4817 24865 4861 24899
rect 4895 24865 4923 24899
rect 4717 24826 4923 24865
rect 4717 24792 4783 24826
rect 4817 24792 4861 24826
rect 4895 24792 4923 24826
rect 4717 24753 4923 24792
rect 4717 24719 4783 24753
rect 4817 24719 4861 24753
rect 4895 24719 4923 24753
rect 4717 24680 4923 24719
rect 4717 24646 4783 24680
rect 4817 24646 4861 24680
rect 4895 24646 4923 24680
rect 4717 24606 4923 24646
rect 4717 24572 4783 24606
rect 4817 24572 4861 24606
rect 4895 24572 4923 24606
rect 4717 24532 4923 24572
rect 4717 24498 4783 24532
rect 4817 24498 4861 24532
rect 4895 24498 4923 24532
rect 4717 24458 4923 24498
rect 4717 24424 4783 24458
rect 4817 24424 4861 24458
rect 4895 24424 4923 24458
rect 4717 24384 4923 24424
rect 4717 24350 4783 24384
rect 4817 24350 4861 24384
rect 4895 24350 4923 24384
rect 4717 24310 4923 24350
rect 4717 24276 4783 24310
rect 4817 24276 4861 24310
rect 4895 24276 4923 24310
rect 4717 24236 4923 24276
rect 4717 24202 4783 24236
rect 4817 24202 4861 24236
rect 4895 24202 4923 24236
rect 4717 24162 4923 24202
rect 4717 24128 4783 24162
rect 4817 24128 4861 24162
rect 4895 24128 4923 24162
rect 4717 24088 4923 24128
rect 4717 24054 4783 24088
rect 4817 24054 4861 24088
rect 4895 24054 4923 24088
rect 4717 24014 4923 24054
rect 4717 23980 4783 24014
rect 4817 23980 4861 24014
rect 4895 23980 4923 24014
rect 4717 23940 4923 23980
rect 4717 23906 4783 23940
rect 4817 23906 4861 23940
rect 4895 23906 4923 23940
rect 4717 23866 4923 23906
rect 4717 23832 4783 23866
rect 4817 23832 4861 23866
rect 4895 23832 4923 23866
rect 4717 23792 4923 23832
rect 4717 23758 4783 23792
rect 4817 23758 4861 23792
rect 4895 23758 4923 23792
rect 4717 23718 4923 23758
rect 4717 23684 4783 23718
rect 4817 23684 4861 23718
rect 4895 23684 4923 23718
rect 4717 23644 4923 23684
rect 4717 23610 4783 23644
rect 4817 23610 4861 23644
rect 4895 23610 4923 23644
rect 4717 23570 4923 23610
rect 4717 23536 4783 23570
rect 4817 23536 4861 23570
rect 4895 23536 4923 23570
rect 4717 23496 4923 23536
rect 4717 23462 4783 23496
rect 4817 23462 4861 23496
rect 4895 23462 4923 23496
rect 4717 23422 4923 23462
rect 4717 23388 4783 23422
rect 4817 23388 4861 23422
rect 4895 23388 4923 23422
rect 4717 23348 4923 23388
rect 4717 23314 4783 23348
rect 4817 23314 4861 23348
rect 4895 23314 4923 23348
rect 4717 23232 4923 23314
rect 12969 27153 13175 27186
rect 5637 23921 5815 23960
rect 5671 23887 5709 23921
rect 5743 23887 5781 23921
rect 5637 23848 5815 23887
rect 5671 23814 5709 23848
rect 5743 23814 5781 23848
rect 5637 23775 5815 23814
rect 5671 23741 5709 23775
rect 5743 23741 5781 23775
rect 5637 23702 5815 23741
rect 5671 23668 5709 23702
rect 5743 23668 5781 23702
rect 5637 23629 5815 23668
rect 5671 23595 5709 23629
rect 5743 23595 5781 23629
rect 5637 23556 5815 23595
rect 5671 23522 5709 23556
rect 5743 23522 5781 23556
rect 5637 23483 5815 23522
rect 5671 23449 5709 23483
rect 5743 23449 5781 23483
rect 5637 23410 5815 23449
rect 5671 23376 5709 23410
rect 5743 23376 5781 23410
rect 5637 23337 5815 23376
rect 5671 23303 5709 23337
rect 5743 23303 5781 23337
rect 12969 26628 12997 27153
rect 12969 23303 12997 23790
rect 12969 23232 13175 23303
rect 13628 27142 13631 27180
rect 13628 27070 13631 27108
rect 13628 26998 13631 27036
rect 13628 26926 13631 26964
rect 13628 26854 13631 26892
rect 13628 26782 13631 26820
rect 13628 26710 13631 26748
rect 13628 26638 13631 26676
rect 13628 26566 13631 26604
rect 13628 26494 13631 26532
rect 13628 26422 13631 26460
rect 13628 26350 13631 26388
rect 13628 26278 13631 26316
rect 13628 26206 13631 26244
rect 13628 26134 13631 26172
rect 13628 26062 13631 26100
rect 13628 25990 13631 26028
rect 13628 25918 13631 25956
rect 13628 25846 13631 25884
rect 13628 25774 13631 25812
rect 13628 25702 13631 25740
rect 13628 25630 13631 25668
rect 13628 25558 13631 25596
rect 13628 25486 13631 25524
rect 13628 25413 13631 25452
rect 13628 25340 13631 25379
rect 13628 25267 13631 25306
rect 13628 25194 13631 25233
rect 13628 25121 13631 25160
rect 13628 25048 13631 25087
rect 13628 24975 13631 25014
rect 13628 24902 13631 24941
rect 13628 24829 13631 24868
rect 13628 24756 13631 24795
rect 13628 24683 13631 24722
rect 13628 24610 13631 24649
rect 13628 24537 13631 24576
rect 13628 24464 13631 24503
rect 13628 24391 13631 24430
rect 13628 24318 13631 24357
rect 13628 24245 13631 24284
rect 13628 24172 13631 24211
rect 13628 24099 13631 24138
rect 13628 24026 13631 24065
rect 13628 23953 13631 23992
rect 13628 23880 13631 23919
rect 13628 23807 13631 23846
rect 13628 23734 13631 23773
rect 13628 23661 13631 23700
rect 13628 23588 13631 23627
rect 13628 23515 13631 23554
rect 13628 23442 13631 23481
rect 13628 23369 13631 23408
rect 13628 23296 13631 23335
rect 13628 23223 13631 23262
rect 4611 23164 5016 23198
rect 5050 23164 5084 23198
rect 5118 23164 5418 23198
rect 5452 23164 5486 23198
rect 5520 23164 5936 23198
rect 5970 23164 6004 23198
rect 6038 23164 6338 23198
rect 6372 23164 6406 23198
rect 6440 23164 6856 23198
rect 6890 23164 6924 23198
rect 6958 23164 7258 23198
rect 7292 23164 7326 23198
rect 7360 23164 7776 23198
rect 7810 23164 7844 23198
rect 7878 23164 8178 23198
rect 8212 23164 8246 23198
rect 8280 23164 8696 23198
rect 8730 23164 8764 23198
rect 8798 23164 9098 23198
rect 9132 23164 9166 23198
rect 9200 23164 9616 23198
rect 9650 23164 9684 23198
rect 9718 23164 10018 23198
rect 10052 23164 10086 23198
rect 10120 23164 10536 23198
rect 10570 23164 10604 23198
rect 10638 23164 10938 23198
rect 10972 23164 11006 23198
rect 11040 23164 11456 23198
rect 11490 23164 11524 23198
rect 11558 23164 11858 23198
rect 11892 23164 11926 23198
rect 11960 23164 12376 23198
rect 12410 23164 12444 23198
rect 12478 23164 12778 23198
rect 12812 23164 12846 23198
rect 12880 23164 12900 23198
rect 4611 22993 12900 23164
rect 4611 22959 4789 22993
rect 4823 22959 12900 22993
rect 4611 22921 12900 22959
rect 4611 22887 4789 22921
rect 4823 22887 12900 22921
rect 4611 22708 12900 22887
rect 4611 22674 5016 22708
rect 5050 22674 5084 22708
rect 5118 22674 5418 22708
rect 5452 22674 5486 22708
rect 5520 22674 5936 22708
rect 5970 22674 6004 22708
rect 6038 22674 6338 22708
rect 6372 22674 6406 22708
rect 6440 22674 6856 22708
rect 6890 22674 6924 22708
rect 6958 22674 7258 22708
rect 7292 22674 7326 22708
rect 7360 22674 7776 22708
rect 7810 22674 7844 22708
rect 7878 22674 8178 22708
rect 8212 22674 8246 22708
rect 8280 22674 8696 22708
rect 8730 22674 8764 22708
rect 8798 22674 9098 22708
rect 9132 22674 9166 22708
rect 9200 22674 9616 22708
rect 9650 22674 9684 22708
rect 9718 22674 10018 22708
rect 10052 22674 10086 22708
rect 10120 22674 10536 22708
rect 10570 22674 10604 22708
rect 10638 22674 10938 22708
rect 10972 22674 11006 22708
rect 11040 22674 11456 22708
rect 11490 22674 11524 22708
rect 11558 22674 11858 22708
rect 11892 22674 11926 22708
rect 11960 22674 12376 22708
rect 12410 22674 12444 22708
rect 12478 22674 12778 22708
rect 12812 22674 12846 22708
rect 12880 22674 12900 22708
rect 4611 22668 12900 22674
rect 13628 23150 13631 23189
rect 13628 23077 13631 23116
rect 13628 23004 13631 23043
rect 13628 22931 13631 22970
rect 13628 22858 13631 22897
rect 13628 22785 13631 22824
rect 13628 22712 13631 22751
rect 13628 22639 13631 22678
rect 4717 22484 4923 22586
rect 4198 18946 4217 18985
rect 4198 18873 4217 18912
rect 4198 18800 4217 18839
rect 4198 18727 4217 18766
rect 4198 18654 4217 18693
rect 4198 18581 4217 18620
rect 4198 18508 4217 18547
rect 4198 18435 4217 18474
rect 4198 18362 4217 18401
rect 4198 18289 4217 18328
rect 4198 18216 4217 18255
rect 4198 18143 4217 18182
rect 4198 18070 4217 18109
rect 4198 17997 4217 18036
rect 4198 17924 4217 17963
rect 4198 17851 4217 17890
rect 4198 17778 4217 17817
rect 4198 17705 4217 17744
rect 4198 17632 4217 17671
rect 4198 17559 4217 17598
rect 4198 17486 4217 17525
rect 4198 17413 4217 17452
rect 4198 17340 4217 17379
rect 4198 17267 4217 17306
rect 4198 17194 4217 17233
rect 4198 17121 4217 17160
rect 4198 17048 4217 17087
rect 4198 16975 4217 17014
rect 4198 16902 4217 16941
rect 4198 16829 4217 16868
rect 4198 16756 4217 16795
rect 4198 16683 4217 16722
rect 4198 16610 4217 16649
rect 4198 16537 4217 16576
rect 4198 16464 4217 16503
rect 4198 16391 4217 16430
rect 4198 16318 4217 16357
rect 4198 16245 4217 16284
rect 4198 16172 4217 16211
rect 4198 16099 4217 16138
rect 4198 16026 4217 16065
rect 4198 15953 4217 15992
rect 4198 15880 4217 15919
rect 4198 15807 4217 15846
rect 4198 15734 4217 15773
rect 4198 15661 4217 15700
rect 4198 15588 4217 15627
rect 4198 15515 4217 15554
rect 4198 15442 4217 15481
rect 4198 15369 4217 15408
rect 4198 15296 4217 15335
rect 4198 15223 4217 15262
rect 4198 15150 4217 15189
rect 4198 15077 4217 15116
rect 4198 15004 4217 15043
rect 4198 14931 4217 14970
rect 1915 14836 1953 14870
rect 3728 14840 3766 14874
rect 4198 14858 4217 14897
rect 4198 14785 4217 14824
rect 4198 14712 4217 14751
rect 4198 14639 4217 14678
rect 3960 14603 3967 14634
rect 4001 14603 4028 14634
rect 3960 14566 4028 14603
rect 4198 14566 4217 14605
rect 3960 14565 4096 14566
rect 3960 14564 4039 14565
rect 1827 14530 1899 14564
rect 1933 14562 1973 14564
rect 2007 14562 2047 14564
rect 2081 14562 2121 14564
rect 2155 14562 2195 14564
rect 2229 14562 2269 14564
rect 2303 14562 2343 14564
rect 2377 14562 2417 14564
rect 2451 14562 2491 14564
rect 2525 14562 2565 14564
rect 2599 14562 2639 14564
rect 2673 14562 2713 14564
rect 2747 14562 2787 14564
rect 2821 14562 2861 14564
rect 2895 14562 2935 14564
rect 2969 14562 3009 14564
rect 3043 14562 3083 14564
rect 3117 14562 3157 14564
rect 3191 14562 3231 14564
rect 3265 14562 3305 14564
rect 3339 14562 3379 14564
rect 3413 14562 3453 14564
rect 3487 14562 3527 14564
rect 3561 14562 3601 14564
rect 3635 14562 3675 14564
rect 3709 14562 3748 14564
rect 3782 14562 3821 14564
rect 3855 14562 3894 14564
rect 3928 14562 3967 14564
rect 1954 14530 1973 14562
rect 4001 14531 4039 14564
rect 4073 14531 4096 14565
rect 4001 14530 4096 14531
rect 1827 14528 1920 14530
rect 1954 14528 1988 14530
rect 1827 14494 1988 14528
rect 3994 14498 4096 14530
rect 4198 14498 4217 14532
rect 3994 14494 4217 14498
rect 1827 14492 1834 14494
rect 1936 14492 1988 14494
rect 4062 14493 4217 14494
rect 4062 14492 4111 14493
rect 1936 14458 1973 14492
rect 2007 14458 2047 14460
rect 4073 14459 4111 14492
rect 4145 14464 4183 14493
rect 4145 14459 4164 14464
rect 4073 14458 4164 14459
rect 1936 14426 2056 14458
rect 4062 14430 4164 14458
rect 4198 14430 4217 14459
rect 4062 14426 4217 14430
rect 2004 14420 2056 14426
rect 4130 14420 4217 14426
rect 2005 14386 2045 14420
rect 2079 14386 2119 14392
rect 4145 14386 4183 14420
rect 2005 14358 2124 14386
rect 2072 14348 2124 14358
rect 4130 14348 4217 14386
rect 2077 14314 2117 14348
rect 2151 14314 2191 14324
rect 2225 14314 2265 14324
rect 2299 14314 2339 14324
rect 2373 14314 2413 14324
rect 2447 14314 2487 14324
rect 2521 14314 2561 14324
rect 2595 14314 2635 14324
rect 2669 14314 2709 14324
rect 2743 14314 2783 14324
rect 2817 14314 2857 14324
rect 2891 14314 2931 14324
rect 2965 14314 3005 14324
rect 3039 14314 3079 14324
rect 3113 14314 3153 14324
rect 3187 14314 3227 14324
rect 3261 14314 3301 14324
rect 3335 14314 3375 14324
rect 3409 14314 3449 14324
rect 3483 14314 3523 14324
rect 3557 14314 3597 14324
rect 3631 14314 3671 14324
rect 3705 14314 3745 14324
rect 3779 14314 3818 14324
rect 3852 14314 3891 14324
rect 3925 14314 3964 14324
rect 3998 14314 4037 14324
rect 4071 14314 4110 14324
rect 4144 14314 4217 14348
rect 4358 18553 4362 18592
rect 4717 18922 4784 22484
rect 4890 18922 4923 22484
rect 4717 18883 4923 18922
rect 4717 18849 4784 18883
rect 4818 18849 4856 18883
rect 4890 18849 4923 18883
rect 4717 18810 4923 18849
rect 4717 18776 4784 18810
rect 4818 18776 4856 18810
rect 4890 18776 4923 18810
rect 4717 18737 4923 18776
rect 4717 18703 4784 18737
rect 4818 18703 4856 18737
rect 4890 18703 4923 18737
rect 12969 22562 13175 22587
rect 5637 19978 5815 20017
rect 5671 19944 5709 19978
rect 5743 19944 5781 19978
rect 5637 19905 5815 19944
rect 5671 19871 5709 19905
rect 5743 19871 5781 19905
rect 5637 19832 5815 19871
rect 5671 19798 5709 19832
rect 5743 19798 5781 19832
rect 5637 19759 5815 19798
rect 5671 19725 5709 19759
rect 5743 19725 5781 19759
rect 5637 19686 5815 19725
rect 5671 19652 5709 19686
rect 5743 19652 5781 19686
rect 5637 19613 5815 19652
rect 5671 19579 5709 19613
rect 5743 19579 5781 19613
rect 5637 19540 5815 19579
rect 5671 19506 5709 19540
rect 5743 19506 5781 19540
rect 5637 19467 5815 19506
rect 5671 19433 5709 19467
rect 5743 19433 5781 19467
rect 5637 19394 5815 19433
rect 5671 19360 5709 19394
rect 5743 19360 5781 19394
rect 5637 19321 5815 19360
rect 5671 19287 5709 19321
rect 5743 19287 5781 19321
rect 5637 19248 5815 19287
rect 5671 19214 5709 19248
rect 5743 19214 5781 19248
rect 5637 19175 5815 19214
rect 5671 19141 5709 19175
rect 5743 19141 5781 19175
rect 5637 19102 5815 19141
rect 5671 19068 5709 19102
rect 5743 19068 5781 19102
rect 5637 19029 5815 19068
rect 5671 18995 5709 19029
rect 5743 18995 5781 19029
rect 5637 18956 5815 18995
rect 5671 18922 5709 18956
rect 5743 18922 5781 18956
rect 5637 18883 5815 18922
rect 5671 18849 5709 18883
rect 5743 18849 5781 18883
rect 5637 18810 5815 18849
rect 5671 18776 5709 18810
rect 5743 18776 5781 18810
rect 5637 18737 5815 18776
rect 5671 18703 5709 18737
rect 5743 18703 5781 18737
rect 6557 19321 6735 19360
rect 6591 19287 6629 19321
rect 6663 19287 6701 19321
rect 6557 19248 6735 19287
rect 6591 19214 6629 19248
rect 6663 19214 6701 19248
rect 6557 19175 6735 19214
rect 6591 19141 6629 19175
rect 6663 19141 6701 19175
rect 6557 19102 6735 19141
rect 6591 19068 6629 19102
rect 6663 19068 6701 19102
rect 6557 19029 6735 19068
rect 6591 18995 6629 19029
rect 6663 18995 6701 19029
rect 6557 18956 6735 18995
rect 6591 18922 6629 18956
rect 6663 18922 6701 18956
rect 6557 18883 6735 18922
rect 6591 18849 6629 18883
rect 6663 18849 6701 18883
rect 6557 18810 6735 18849
rect 6591 18776 6629 18810
rect 6663 18776 6701 18810
rect 6557 18737 6735 18776
rect 6591 18703 6629 18737
rect 6663 18703 6701 18737
rect 7477 19321 7655 19360
rect 7511 19287 7549 19321
rect 7583 19287 7621 19321
rect 7477 19248 7655 19287
rect 7511 19214 7549 19248
rect 7583 19214 7621 19248
rect 7477 19175 7655 19214
rect 7511 19141 7549 19175
rect 7583 19141 7621 19175
rect 7477 19102 7655 19141
rect 7511 19068 7549 19102
rect 7583 19068 7621 19102
rect 7477 19029 7655 19068
rect 7511 18995 7549 19029
rect 7583 18995 7621 19029
rect 7477 18956 7655 18995
rect 7511 18922 7549 18956
rect 7583 18922 7621 18956
rect 7477 18883 7655 18922
rect 7511 18849 7549 18883
rect 7583 18849 7621 18883
rect 7477 18810 7655 18849
rect 7511 18776 7549 18810
rect 7583 18776 7621 18810
rect 7477 18737 7655 18776
rect 7511 18703 7549 18737
rect 7583 18703 7621 18737
rect 8397 19321 8575 19360
rect 8431 19287 8469 19321
rect 8503 19287 8541 19321
rect 8397 19248 8575 19287
rect 8431 19214 8469 19248
rect 8503 19214 8541 19248
rect 8397 19175 8575 19214
rect 8431 19141 8469 19175
rect 8503 19141 8541 19175
rect 8397 19102 8575 19141
rect 8431 19068 8469 19102
rect 8503 19068 8541 19102
rect 8397 19029 8575 19068
rect 8431 18995 8469 19029
rect 8503 18995 8541 19029
rect 8397 18956 8575 18995
rect 8431 18922 8469 18956
rect 8503 18922 8541 18956
rect 8397 18883 8575 18922
rect 8431 18849 8469 18883
rect 8503 18849 8541 18883
rect 8397 18810 8575 18849
rect 8431 18776 8469 18810
rect 8503 18776 8541 18810
rect 8397 18737 8575 18776
rect 8431 18703 8469 18737
rect 8503 18703 8541 18737
rect 9317 19321 9495 19360
rect 9351 19287 9389 19321
rect 9423 19287 9461 19321
rect 9317 19248 9495 19287
rect 9351 19214 9389 19248
rect 9423 19214 9461 19248
rect 9317 19175 9495 19214
rect 9351 19141 9389 19175
rect 9423 19141 9461 19175
rect 9317 19102 9495 19141
rect 9351 19068 9389 19102
rect 9423 19068 9461 19102
rect 9317 19029 9495 19068
rect 9351 18995 9389 19029
rect 9423 18995 9461 19029
rect 9317 18956 9495 18995
rect 9351 18922 9389 18956
rect 9423 18922 9461 18956
rect 9317 18883 9495 18922
rect 9351 18849 9389 18883
rect 9423 18849 9461 18883
rect 9317 18810 9495 18849
rect 9351 18776 9389 18810
rect 9423 18776 9461 18810
rect 9317 18737 9495 18776
rect 9351 18703 9389 18737
rect 9423 18703 9461 18737
rect 10237 19321 10415 19360
rect 10271 19287 10309 19321
rect 10343 19287 10381 19321
rect 10237 19248 10415 19287
rect 10271 19214 10309 19248
rect 10343 19214 10381 19248
rect 10237 19175 10415 19214
rect 10271 19141 10309 19175
rect 10343 19141 10381 19175
rect 10237 19102 10415 19141
rect 10271 19068 10309 19102
rect 10343 19068 10381 19102
rect 10237 19029 10415 19068
rect 10271 18995 10309 19029
rect 10343 18995 10381 19029
rect 10237 18956 10415 18995
rect 10271 18922 10309 18956
rect 10343 18922 10381 18956
rect 10237 18883 10415 18922
rect 10271 18849 10309 18883
rect 10343 18849 10381 18883
rect 10237 18810 10415 18849
rect 10271 18776 10309 18810
rect 10343 18776 10381 18810
rect 10237 18737 10415 18776
rect 10271 18703 10309 18737
rect 10343 18703 10381 18737
rect 11157 19321 11335 19360
rect 11191 19287 11229 19321
rect 11263 19287 11301 19321
rect 11157 19248 11335 19287
rect 11191 19214 11229 19248
rect 11263 19214 11301 19248
rect 11157 19175 11335 19214
rect 11191 19141 11229 19175
rect 11263 19141 11301 19175
rect 11157 19102 11335 19141
rect 11191 19068 11229 19102
rect 11263 19068 11301 19102
rect 11157 19029 11335 19068
rect 11191 18995 11229 19029
rect 11263 18995 11301 19029
rect 11157 18956 11335 18995
rect 11191 18922 11229 18956
rect 11263 18922 11301 18956
rect 11157 18883 11335 18922
rect 11191 18849 11229 18883
rect 11263 18849 11301 18883
rect 11157 18810 11335 18849
rect 11191 18776 11229 18810
rect 11263 18776 11301 18810
rect 11157 18737 11335 18776
rect 11191 18703 11229 18737
rect 11263 18703 11301 18737
rect 12969 22029 12997 22562
rect 12077 19321 12255 19360
rect 12111 19287 12149 19321
rect 12183 19287 12221 19321
rect 12077 19248 12255 19287
rect 12111 19214 12149 19248
rect 12183 19214 12221 19248
rect 12077 19175 12255 19214
rect 13628 22566 13631 22605
rect 13628 22493 13631 22532
rect 13628 22420 13631 22459
rect 13628 22347 13631 22386
rect 13628 22274 13631 22313
rect 13628 22201 13631 22240
rect 13628 22128 13631 22167
rect 13628 22055 13631 22094
rect 13628 21982 13631 22021
rect 13628 21909 13631 21948
rect 13628 21836 13631 21875
rect 13628 21763 13631 21802
rect 13628 21690 13631 21729
rect 13628 21617 13631 21656
rect 13628 21544 13631 21583
rect 13628 21471 13631 21510
rect 13628 21398 13631 21437
rect 13628 21325 13631 21364
rect 13628 21252 13631 21291
rect 13628 21179 13631 21218
rect 13628 21106 13631 21145
rect 13628 21033 13631 21072
rect 13628 20960 13631 20999
rect 13628 20887 13631 20926
rect 13628 20814 13631 20853
rect 13628 20741 13631 20780
rect 13628 20668 13631 20707
rect 13628 20595 13631 20634
rect 13628 20522 13631 20561
rect 13628 20449 13631 20488
rect 13628 20376 13631 20415
rect 13775 32657 13781 32712
rect 14019 32657 14025 32712
rect 13775 32584 13781 32623
rect 14019 32584 14025 32623
rect 13775 32511 13781 32550
rect 14019 32511 14025 32550
rect 13775 32438 13781 32477
rect 14019 32438 14025 32477
rect 13775 32365 13781 32404
rect 14019 32365 14025 32404
rect 13775 32292 13781 32331
rect 14019 32292 14025 32331
rect 13775 32219 13781 32258
rect 14019 32219 14025 32258
rect 13775 32146 13781 32185
rect 14019 32146 14025 32185
rect 13775 32073 13781 32112
rect 14019 32073 14025 32112
rect 13775 32000 13781 32039
rect 14019 32000 14025 32039
rect 13775 31927 13781 31966
rect 14019 31927 14025 31966
rect 13775 31854 13781 31893
rect 14019 31854 14025 31893
rect 13775 31781 13781 31820
rect 14019 31781 14025 31820
rect 13775 31708 13781 31747
rect 14019 31708 14025 31747
rect 13775 31635 13781 31674
rect 14019 31635 14025 31674
rect 13775 31562 13781 31601
rect 14019 31562 14025 31601
rect 13775 31489 13781 31528
rect 14019 31489 14025 31528
rect 13775 31416 13781 31455
rect 14019 31416 14025 31455
rect 13775 31343 13781 31382
rect 14019 31343 14025 31382
rect 13775 31270 13781 31309
rect 14019 31270 14025 31309
rect 13775 31197 13781 31236
rect 14019 31197 14025 31236
rect 13775 31124 13781 31163
rect 14019 31124 14025 31163
rect 13775 31051 13781 31090
rect 14019 31051 14025 31090
rect 13775 30978 13781 31017
rect 14019 30978 14025 31017
rect 13775 30905 13781 30944
rect 14019 30905 14025 30944
rect 13775 30832 13781 30871
rect 14019 30832 14025 30871
rect 13775 30759 13781 30798
rect 14019 30759 14025 30798
rect 13775 30686 13781 30725
rect 14019 30686 14025 30725
rect 13775 30613 13781 30652
rect 14019 30613 14025 30652
rect 13775 30540 13781 30579
rect 14019 30540 14025 30579
rect 13775 30467 13781 30506
rect 14019 30467 14025 30506
rect 13775 30394 13781 30433
rect 14019 30394 14025 30433
rect 13775 30321 13781 30360
rect 14019 30321 14025 30360
rect 13775 30248 13781 30287
rect 14019 30248 14025 30287
rect 13775 30175 13781 30214
rect 14019 30175 14025 30214
rect 13775 30102 13781 30141
rect 14019 30102 14025 30141
rect 13775 30029 13781 30068
rect 14019 30029 14025 30068
rect 13775 29956 13781 29995
rect 14019 29956 14025 29995
rect 13775 29883 13781 29922
rect 14019 29883 14025 29922
rect 13775 29810 13781 29849
rect 14019 29810 14025 29849
rect 13775 29737 13781 29776
rect 14019 29737 14025 29776
rect 13775 29664 13781 29703
rect 14019 29664 14025 29703
rect 13775 29591 13781 29630
rect 14019 29591 14025 29630
rect 13775 29518 13781 29557
rect 14019 29518 14025 29557
rect 13775 29445 13781 29484
rect 14019 29445 14025 29484
rect 13775 29372 13781 29411
rect 14019 29372 14025 29411
rect 13775 29299 13781 29338
rect 14019 29299 14025 29338
rect 13775 29226 13781 29265
rect 14019 29226 14025 29265
rect 13775 29153 13781 29192
rect 14019 29153 14025 29192
rect 13775 29080 13781 29119
rect 14019 29080 14025 29119
rect 13775 29007 13781 29046
rect 14019 29007 14025 29046
rect 13775 28934 13781 28973
rect 14019 28934 14025 28973
rect 13775 28861 13781 28900
rect 14019 28861 14025 28900
rect 13775 28788 13781 28827
rect 14019 28788 14025 28827
rect 13775 28715 13781 28754
rect 14019 28715 14025 28754
rect 13775 28642 13781 28681
rect 14019 28642 14025 28681
rect 13775 28569 13781 28608
rect 14019 28569 14025 28608
rect 13775 28496 13781 28535
rect 14019 28496 14025 28535
rect 13775 28423 13781 28462
rect 14019 28423 14025 28462
rect 12997 19321 13175 19360
rect 13031 19287 13069 19321
rect 13103 19287 13141 19321
rect 12997 19248 13175 19287
rect 13031 19214 13069 19248
rect 13103 19214 13141 19248
rect 12997 19190 13175 19214
rect 12111 19141 12149 19175
rect 12183 19141 12221 19175
rect 12077 19102 12255 19141
rect 12111 19068 12149 19102
rect 12183 19068 12221 19102
rect 12077 19029 12255 19068
rect 12111 18995 12149 19029
rect 12183 18995 12221 19029
rect 12077 18956 12255 18995
rect 12111 18922 12149 18956
rect 12183 18922 12221 18956
rect 12077 18883 12255 18922
rect 12111 18849 12149 18883
rect 12183 18849 12221 18883
rect 12077 18810 12255 18849
rect 12111 18776 12149 18810
rect 12183 18776 12221 18810
rect 12077 18737 12255 18776
rect 12111 18703 12149 18737
rect 12183 18703 12221 18737
rect 12969 19175 13175 19190
rect 12969 19141 12997 19175
rect 13031 19141 13069 19175
rect 13103 19141 13141 19175
rect 12969 19102 13175 19141
rect 12969 19068 12997 19102
rect 13031 19068 13069 19102
rect 13103 19068 13141 19102
rect 12969 19029 13175 19068
rect 12969 18995 12997 19029
rect 13031 18995 13069 19029
rect 13103 18995 13141 19029
rect 12969 18956 13175 18995
rect 12969 18922 12997 18956
rect 13031 18922 13069 18956
rect 13103 18922 13141 18956
rect 12969 18883 13175 18922
rect 12969 18849 12997 18883
rect 13031 18849 13069 18883
rect 13103 18849 13141 18883
rect 12969 18810 13175 18849
rect 12969 18776 12997 18810
rect 13031 18776 13069 18810
rect 13103 18776 13141 18810
rect 12969 18737 13175 18776
rect 12969 18703 12997 18737
rect 13031 18703 13069 18737
rect 13103 18703 13141 18737
rect 4717 18632 4923 18703
rect 12969 18632 13175 18703
rect 13453 20190 13458 20229
rect 13628 20190 13631 20229
rect 13453 20117 13458 20156
rect 13628 20117 13631 20156
rect 13453 20044 13458 20083
rect 13628 20044 13631 20083
rect 13453 19971 13458 20010
rect 13628 19971 13631 20010
rect 13453 19898 13458 19937
rect 13628 19898 13631 19937
rect 13453 19825 13458 19864
rect 13628 19825 13631 19864
rect 13453 19752 13458 19791
rect 13628 19752 13631 19791
rect 13453 19679 13458 19718
rect 13628 19679 13631 19718
rect 13453 19606 13458 19645
rect 13628 19606 13631 19645
rect 13453 19533 13458 19572
rect 13628 19533 13631 19572
rect 13453 19460 13458 19499
rect 13628 19460 13631 19499
rect 13453 19387 13458 19426
rect 13628 19387 13631 19426
rect 13453 19314 13458 19353
rect 13628 19314 13631 19353
rect 13453 19241 13458 19280
rect 13628 19241 13631 19280
rect 13453 19168 13458 19207
rect 13628 19168 13631 19207
rect 13453 19095 13458 19134
rect 13628 19095 13631 19134
rect 13453 19022 13458 19061
rect 13628 19022 13631 19061
rect 13453 18949 13458 18988
rect 13628 18949 13631 18988
rect 13453 18876 13458 18915
rect 13628 18876 13631 18915
rect 13453 18803 13458 18842
rect 13628 18803 13631 18842
rect 13453 18730 13458 18769
rect 13628 18730 13631 18769
rect 13453 18657 13458 18696
rect 13628 18657 13631 18696
rect 4358 18480 4362 18519
rect 4532 18481 4536 18520
rect 4358 18407 4362 18446
rect 4532 18408 4536 18447
rect 4358 18334 4362 18373
rect 4532 18335 4536 18374
rect 4358 18261 4362 18300
rect 4532 18262 4536 18301
rect 4358 18188 4362 18227
rect 4532 18189 4536 18228
rect 4358 18115 4362 18154
rect 4532 18116 4536 18155
rect 4605 18586 5016 18598
rect 4605 18552 4611 18586
rect 4645 18564 5016 18586
rect 5050 18564 5084 18598
rect 5118 18564 5418 18598
rect 5452 18564 5486 18598
rect 5520 18564 5936 18598
rect 5970 18564 6004 18598
rect 6038 18564 6338 18598
rect 6372 18564 6406 18598
rect 6440 18564 6856 18598
rect 6890 18564 6924 18598
rect 6958 18564 7258 18598
rect 7292 18564 7326 18598
rect 7360 18564 7776 18598
rect 7810 18564 7844 18598
rect 7878 18564 8178 18598
rect 8212 18564 8246 18598
rect 8280 18564 8696 18598
rect 8730 18564 8764 18598
rect 8798 18564 9098 18598
rect 9132 18564 9166 18598
rect 9200 18564 9616 18598
rect 9650 18564 9684 18598
rect 9718 18564 10018 18598
rect 10052 18564 10086 18598
rect 10120 18564 10536 18598
rect 10570 18564 10604 18598
rect 10638 18564 10938 18598
rect 10972 18564 11006 18598
rect 11040 18564 11456 18598
rect 11490 18564 11524 18598
rect 11558 18564 11858 18598
rect 11892 18564 11926 18598
rect 11960 18564 12376 18598
rect 12410 18564 12444 18598
rect 12478 18564 12778 18598
rect 12812 18564 12846 18598
rect 12880 18564 12900 18598
rect 4645 18552 12900 18564
rect 4605 18513 12900 18552
rect 4605 18479 4611 18513
rect 4645 18479 12900 18513
rect 4605 18440 12900 18479
rect 4605 18406 4611 18440
rect 4645 18406 12900 18440
rect 4605 18367 12900 18406
rect 4605 18333 4611 18367
rect 4645 18333 12900 18367
rect 4605 18293 12900 18333
rect 4605 18259 4611 18293
rect 4645 18259 12900 18293
rect 4605 18219 12900 18259
rect 4605 18185 4611 18219
rect 4645 18185 12900 18219
rect 4605 18145 12900 18185
rect 4605 18111 4611 18145
rect 4645 18111 12900 18145
rect 4605 18108 12900 18111
rect 4605 18099 5016 18108
rect 4358 18042 4362 18081
rect 4532 18043 4536 18082
rect 4996 18074 5016 18099
rect 5050 18074 5084 18108
rect 5118 18074 5418 18108
rect 5452 18074 5486 18108
rect 5520 18074 5936 18108
rect 5970 18074 6004 18108
rect 6038 18074 6338 18108
rect 6372 18074 6406 18108
rect 6440 18074 6856 18108
rect 6890 18074 6924 18108
rect 6958 18074 7258 18108
rect 7292 18074 7326 18108
rect 7360 18074 7776 18108
rect 7810 18074 7844 18108
rect 7878 18074 8178 18108
rect 8212 18074 8246 18108
rect 8280 18074 8696 18108
rect 8730 18074 8764 18108
rect 8798 18074 9098 18108
rect 9132 18074 9166 18108
rect 9200 18074 9616 18108
rect 9650 18074 9684 18108
rect 9718 18074 10018 18108
rect 10052 18074 10086 18108
rect 10120 18074 10536 18108
rect 10570 18074 10604 18108
rect 10638 18074 10938 18108
rect 10972 18074 11006 18108
rect 11040 18074 11456 18108
rect 11490 18074 11524 18108
rect 11558 18074 11858 18108
rect 11892 18074 11926 18108
rect 11960 18074 12376 18108
rect 12410 18074 12444 18108
rect 12478 18074 12778 18108
rect 12812 18074 12846 18108
rect 12880 18074 12900 18108
rect 5134 18068 12900 18074
rect 13453 18584 13458 18623
rect 13628 18584 13631 18623
rect 13453 18511 13458 18550
rect 13628 18511 13631 18550
rect 13453 18438 13458 18477
rect 13628 18438 13631 18477
rect 13453 18365 13458 18404
rect 13628 18365 13631 18404
rect 13453 18292 13458 18331
rect 13628 18292 13631 18331
rect 13453 18219 13458 18258
rect 13628 18219 13631 18258
rect 13453 18146 13458 18185
rect 13628 18146 13631 18185
rect 13453 18073 13458 18112
rect 13628 18073 13631 18112
rect 4358 17969 4362 18008
rect 4532 17970 4536 18009
rect 13453 18000 13458 18039
rect 13628 18000 13631 18039
rect 4358 17896 4362 17935
rect 4532 17897 4536 17936
rect 4358 17823 4362 17862
rect 4532 17824 4536 17863
rect 4358 17750 4362 17789
rect 4532 17751 4536 17790
rect 4358 17677 4362 17716
rect 4532 17678 4536 17717
rect 4358 17604 4362 17643
rect 4532 17605 4536 17644
rect 4358 17531 4362 17570
rect 4532 17532 4536 17571
rect 4358 17458 4362 17497
rect 4532 17459 4536 17498
rect 4358 17385 4362 17424
rect 4532 17386 4536 17425
rect 4358 17312 4362 17351
rect 4532 17313 4536 17352
rect 4358 17239 4362 17278
rect 4532 17240 4536 17279
rect 4358 17166 4362 17205
rect 4532 17167 4536 17206
rect 4358 17093 4362 17132
rect 4532 17094 4536 17133
rect 4358 17020 4362 17059
rect 4532 17021 4536 17060
rect 4358 16947 4362 16986
rect 4532 16948 4536 16987
rect 4358 16874 4362 16913
rect 4532 16875 4536 16914
rect 4358 16801 4362 16840
rect 4532 16802 4536 16841
rect 4358 16728 4362 16767
rect 4532 16729 4536 16768
rect 4358 16655 4362 16694
rect 4532 16656 4536 16695
rect 4358 16582 4362 16621
rect 4532 16583 4536 16622
rect 4358 16509 4362 16548
rect 4532 16510 4536 16549
rect 4358 16436 4362 16475
rect 4532 16437 4536 16476
rect 4358 16363 4362 16402
rect 4532 16364 4536 16403
rect 4358 16290 4362 16329
rect 4532 16291 4536 16330
rect 4358 16217 4362 16256
rect 4532 16218 4536 16257
rect 4358 16144 4362 16183
rect 4532 16145 4536 16184
rect 4358 16071 4362 16110
rect 4532 16072 4536 16111
rect 4358 15998 4362 16037
rect 4532 15999 4536 16038
rect 4358 15925 4362 15964
rect 4532 15926 4536 15965
rect 4358 15852 4362 15891
rect 4532 15853 4536 15892
rect 4358 15779 4362 15818
rect 4532 15780 4536 15819
rect 4358 15706 4362 15745
rect 4532 15707 4536 15746
rect 4358 15633 4362 15672
rect 4532 15634 4536 15673
rect 4358 15560 4362 15599
rect 4532 15561 4536 15600
rect 4358 15487 4362 15526
rect 4532 15488 4536 15527
rect 4358 15414 4362 15453
rect 4532 15415 4536 15454
rect 4358 15341 4362 15380
rect 4532 15342 4536 15381
rect 4358 15268 4362 15307
rect 4532 15269 4536 15308
rect 4358 15195 4362 15234
rect 4532 15196 4536 15235
rect 4358 15122 4362 15161
rect 4532 15123 4536 15162
rect 4358 15049 4362 15088
rect 4532 15050 4536 15089
rect 4358 14976 4362 15015
rect 4532 14977 4536 15016
rect 4358 14903 4362 14942
rect 4532 14904 4536 14943
rect 4358 14830 4362 14869
rect 4532 14831 4536 14870
rect 4358 14757 4362 14796
rect 4532 14758 4536 14797
rect 4358 14684 4362 14723
rect 4532 14685 4536 14724
rect 4358 14611 4362 14650
rect 4532 14612 4536 14651
rect 4358 14538 4362 14577
rect 4532 14539 4536 14578
rect 4358 14465 4362 14504
rect 4532 14466 4536 14505
rect 4358 14392 4362 14431
rect 4532 14393 4536 14432
rect 4358 14319 4362 14358
rect 4532 14320 4536 14359
rect 4358 14246 4362 14285
rect 4532 14247 4536 14286
rect 4358 14211 4362 14212
rect 4358 14173 4430 14211
rect 4532 14174 4536 14213
rect 1827 13843 1834 13882
rect 2072 13843 2077 13882
rect 1827 13770 1834 13809
rect 2072 13770 2077 13809
rect 1827 13697 1834 13736
rect 2072 13697 2077 13736
rect 1827 13624 1834 13663
rect 2072 13624 2077 13663
rect 1827 13543 1834 13590
rect 2072 13543 2077 13590
rect 2072 12966 2077 13005
rect 1827 12822 1834 12861
rect 2072 12893 2077 12932
rect 1827 12749 1834 12788
rect 2072 12820 2077 12859
rect 1827 12676 1834 12715
rect 2072 12747 2077 12786
rect 1827 12603 1834 12642
rect 2072 12674 2077 12713
rect 1827 12530 1834 12569
rect 2072 12601 2077 12640
rect 1827 12457 1834 12496
rect 2072 12528 2077 12567
rect 1827 12384 1834 12423
rect 2072 12455 2077 12494
rect 1827 12311 1834 12350
rect 2072 12382 2077 12421
rect 1827 12238 1834 12277
rect 2072 12309 2077 12348
rect 1827 12165 1834 12204
rect 2072 12236 2077 12275
rect 1827 12092 1834 12131
rect 2072 12163 2077 12202
rect 1827 12019 1834 12058
rect 2072 12090 2077 12129
rect 1827 11946 1834 11985
rect 2072 12017 2077 12056
rect 1827 11873 1834 11912
rect 2072 11944 2077 11983
rect 1827 11800 1834 11839
rect 2072 11871 2077 11910
rect 1827 11727 1834 11766
rect 2072 11798 2077 11837
rect 1827 11654 1834 11693
rect 2072 11725 2077 11764
rect 1827 11581 1834 11620
rect 2072 11652 2077 11691
rect 1827 11508 1834 11547
rect 2072 11579 2077 11618
rect 1827 11435 1834 11474
rect 2072 11506 2077 11545
rect 1827 11362 1834 11401
rect 2072 11433 2077 11472
rect 1827 11289 1834 11328
rect 2072 11360 2077 11399
rect 1827 11216 1834 11255
rect 2072 11287 2077 11326
rect 1827 11143 1834 11182
rect 2072 11214 2077 11253
rect 1827 11070 1834 11109
rect 2072 11141 2077 11180
rect 1827 10997 1834 11036
rect 2072 11068 2077 11107
rect 1827 10924 1834 10963
rect 2072 10995 2077 11034
rect 1827 10856 1834 10890
rect 2072 10922 2077 10961
rect 2072 10856 2077 10888
rect 1827 10851 2077 10856
rect 1861 10817 1899 10851
rect 1933 10850 2077 10851
rect 1933 10817 1971 10850
rect 1827 10816 1971 10817
rect 2005 10849 2077 10850
rect 2005 10816 2043 10849
rect 1827 10815 2043 10816
rect 1827 10778 2077 10815
rect 1861 10746 1899 10778
rect 1933 10777 2077 10778
rect 1933 10746 1971 10777
rect 2005 10776 2077 10777
rect 2005 10746 2043 10776
rect 1827 10705 1834 10744
rect 1827 10632 1834 10671
rect 2072 10703 2077 10742
rect 1827 10559 1834 10598
rect 2072 10630 2077 10669
rect 1827 10486 1834 10525
rect 2072 10557 2077 10596
rect 1827 10413 1834 10452
rect 2072 10484 2077 10523
rect 1827 10340 1834 10379
rect 2072 10411 2077 10450
rect 1827 10267 1834 10306
rect 2072 10338 2077 10377
rect 1827 10194 1834 10233
rect 2072 10265 2077 10304
rect 1827 10121 1834 10160
rect 2072 10192 2077 10231
rect 1827 10048 1834 10087
rect 2072 10119 2077 10158
rect 1827 9975 1834 10014
rect 2072 10046 2077 10085
rect 1827 9902 1834 9941
rect 2072 9973 2077 10012
rect 1827 9829 1834 9868
rect 2072 9900 2077 9939
rect 1827 9756 1834 9795
rect 2072 9827 2077 9866
rect 1827 9683 1834 9722
rect 2072 9754 2077 9793
rect 1827 9610 1834 9649
rect 2072 9681 2077 9720
rect 1827 9537 1834 9576
rect 2072 9608 2077 9647
rect 1827 9464 1834 9503
rect 2072 9535 2077 9574
rect 1827 9391 1834 9430
rect 2072 9462 2077 9501
rect 1827 9318 1834 9357
rect 2072 9389 2077 9428
rect 1827 9245 1834 9284
rect 2072 9316 2077 9355
rect 1827 9172 1834 9211
rect 2072 9243 2077 9282
rect 1827 9099 1834 9138
rect 2072 9170 2077 9209
rect 1827 9026 1834 9065
rect 2072 9097 2077 9136
rect 2221 14139 2293 14173
rect 2327 14169 2367 14173
rect 2401 14169 2441 14173
rect 2475 14169 2515 14173
rect 2549 14169 2589 14173
rect 2623 14169 2663 14173
rect 2697 14169 2737 14173
rect 2771 14169 2811 14173
rect 2845 14169 2885 14173
rect 2919 14169 2959 14173
rect 2993 14169 3033 14173
rect 3067 14169 3107 14173
rect 3141 14169 3181 14173
rect 3215 14169 3255 14173
rect 3289 14169 3329 14173
rect 3363 14169 3403 14173
rect 3437 14169 3477 14173
rect 3511 14169 3551 14173
rect 3585 14169 3625 14173
rect 3659 14169 3699 14173
rect 3733 14169 3773 14173
rect 3807 14169 3847 14173
rect 3881 14169 3920 14173
rect 3954 14169 3993 14173
rect 4027 14169 4066 14173
rect 4100 14169 4139 14173
rect 4173 14169 4212 14173
rect 4246 14169 4285 14173
rect 4319 14169 4358 14173
rect 4392 14169 4430 14173
rect 2356 14139 2367 14169
rect 4396 14140 4430 14169
rect 4464 14140 4502 14143
rect 2221 14135 2322 14139
rect 2356 14135 2390 14139
rect 2221 14101 2390 14135
rect 4396 14109 4536 14140
rect 4396 14101 4498 14109
rect 4532 14101 4536 14109
rect 2221 14095 2225 14101
rect 2327 14067 2367 14101
rect 4464 14075 4498 14101
rect 4464 14067 4502 14075
rect 2221 14017 2225 14061
rect 2327 14033 2458 14067
rect 2395 14029 2458 14033
rect 2399 13995 2439 14029
rect 4464 13999 4536 14067
rect 4717 17962 4923 17986
rect 4895 14760 4923 17962
rect 4717 14721 4923 14760
rect 4751 14687 4789 14721
rect 4823 14687 4861 14721
rect 4895 14687 4923 14721
rect 4717 14648 4923 14687
rect 4751 14614 4789 14648
rect 4823 14614 4861 14648
rect 4895 14614 4923 14648
rect 4717 14575 4923 14614
rect 4751 14541 4789 14575
rect 4823 14541 4861 14575
rect 4895 14541 4923 14575
rect 4717 14502 4923 14541
rect 4751 14468 4789 14502
rect 4823 14468 4861 14502
rect 4895 14468 4923 14502
rect 4717 14429 4923 14468
rect 4751 14395 4789 14429
rect 4823 14395 4861 14429
rect 4895 14395 4923 14429
rect 4717 14356 4923 14395
rect 4751 14322 4789 14356
rect 4823 14322 4861 14356
rect 4895 14322 4923 14356
rect 4717 14283 4923 14322
rect 4751 14249 4789 14283
rect 4823 14249 4861 14283
rect 4895 14249 4923 14283
rect 4717 14210 4923 14249
rect 4751 14176 4789 14210
rect 4823 14176 4861 14210
rect 4895 14176 4923 14210
rect 4717 14137 4923 14176
rect 4751 14103 4789 14137
rect 4823 14103 4861 14137
rect 4895 14103 4923 14137
rect 12969 17953 13175 17986
rect 5637 14721 5815 14760
rect 5671 14687 5709 14721
rect 5743 14687 5781 14721
rect 5637 14648 5815 14687
rect 5671 14614 5709 14648
rect 5743 14614 5781 14648
rect 5637 14575 5815 14614
rect 5671 14541 5709 14575
rect 5743 14541 5781 14575
rect 5637 14502 5815 14541
rect 5671 14468 5709 14502
rect 5743 14468 5781 14502
rect 5637 14429 5815 14468
rect 5671 14395 5709 14429
rect 5743 14395 5781 14429
rect 5637 14356 5815 14395
rect 5671 14322 5709 14356
rect 5743 14322 5781 14356
rect 5637 14283 5815 14322
rect 5671 14249 5709 14283
rect 5743 14249 5781 14283
rect 5637 14210 5815 14249
rect 5671 14176 5709 14210
rect 5743 14176 5781 14210
rect 5637 14137 5815 14176
rect 5671 14103 5709 14137
rect 5743 14103 5781 14137
rect 12969 17428 12997 17953
rect 12969 14103 12997 14590
rect 4717 14032 4923 14103
rect 12969 14032 13175 14103
rect 13453 17927 13458 17966
rect 13628 17927 13631 17966
rect 13453 17854 13458 17893
rect 13628 17854 13631 17893
rect 13453 17781 13458 17820
rect 13628 17781 13631 17820
rect 13453 17708 13458 17747
rect 13628 17708 13631 17747
rect 13453 17635 13458 17674
rect 13628 17635 13631 17674
rect 13453 17562 13458 17601
rect 13628 17562 13631 17601
rect 13453 17489 13458 17528
rect 13628 17489 13631 17528
rect 13453 17416 13458 17455
rect 13628 17416 13631 17455
rect 13453 17343 13458 17382
rect 13628 17343 13631 17382
rect 13453 17270 13458 17309
rect 13628 17270 13631 17309
rect 13453 17197 13458 17236
rect 13628 17197 13631 17236
rect 13453 17124 13458 17163
rect 13628 17124 13631 17163
rect 13453 17051 13458 17090
rect 13628 17051 13631 17090
rect 13453 16978 13458 17017
rect 13628 16978 13631 17017
rect 13453 16905 13458 16944
rect 13628 16905 13631 16944
rect 13453 16832 13458 16871
rect 13628 16832 13631 16871
rect 13453 16759 13458 16798
rect 13628 16759 13631 16798
rect 13453 16686 13458 16725
rect 13628 16686 13631 16725
rect 2473 13995 2513 13999
rect 2547 13995 2587 13999
rect 2621 13995 2661 13999
rect 2695 13995 2735 13999
rect 2769 13995 2809 13999
rect 2843 13995 2883 13999
rect 2917 13995 2957 13999
rect 2991 13995 3031 13999
rect 3065 13995 3105 13999
rect 3139 13995 3179 13999
rect 3213 13995 3253 13999
rect 3287 13995 3327 13999
rect 3361 13995 3401 13999
rect 3435 13995 3475 13999
rect 3509 13995 3549 13999
rect 3583 13995 3623 13999
rect 3657 13995 3697 13999
rect 3731 13995 3771 13999
rect 3805 13995 3845 13999
rect 3879 13995 3918 13999
rect 3952 13995 3991 13999
rect 4025 13995 4064 13999
rect 4098 13995 4137 13999
rect 4171 13995 4210 13999
rect 4244 13995 4283 13999
rect 4317 13995 4356 13999
rect 4390 13995 4429 13999
rect 4463 13995 4536 13999
rect 2221 13939 2225 13983
rect 2395 13949 2399 13995
rect 2221 13861 2225 13905
rect 2395 13869 2399 13915
rect 2221 13783 2225 13827
rect 2395 13789 2399 13835
rect 4702 13964 5016 13998
rect 5050 13964 5084 13998
rect 5118 13964 5418 13998
rect 5452 13964 5486 13998
rect 5520 13964 5936 13998
rect 5970 13964 6004 13998
rect 6038 13964 6338 13998
rect 6372 13964 6406 13998
rect 6440 13964 6856 13998
rect 6890 13964 6924 13998
rect 6958 13964 7258 13998
rect 7292 13964 7326 13998
rect 7360 13964 7776 13998
rect 7810 13964 7844 13998
rect 7878 13964 8178 13998
rect 8212 13964 8246 13998
rect 8280 13964 8696 13998
rect 8730 13964 8764 13998
rect 8798 13964 9098 13998
rect 9132 13964 9166 13998
rect 9200 13964 9616 13998
rect 9650 13964 9684 13998
rect 9718 13964 10018 13998
rect 10052 13964 10086 13998
rect 10120 13964 10536 13998
rect 10570 13964 10604 13998
rect 10638 13964 10938 13998
rect 10972 13964 11006 13998
rect 11040 13964 11456 13998
rect 11490 13964 11524 13998
rect 11558 13964 11858 13998
rect 11892 13964 11926 13998
rect 11960 13964 12376 13998
rect 12410 13964 12444 13998
rect 12478 13964 12778 13998
rect 12812 13964 12846 13998
rect 12880 13964 12900 13998
rect 4702 13799 12900 13964
rect 2221 13705 2225 13749
rect 2395 13708 2399 13755
rect 2221 13627 2225 13671
rect 2395 13627 2399 13674
rect 3141 13642 12900 13799
rect 3141 13608 3157 13642
rect 3191 13608 3230 13642
rect 3264 13608 3303 13642
rect 3337 13608 3376 13642
rect 3410 13608 3449 13642
rect 3483 13608 3522 13642
rect 3556 13608 3595 13642
rect 3629 13608 3668 13642
rect 3702 13608 3741 13642
rect 3775 13608 3813 13642
rect 3847 13608 3885 13642
rect 3919 13608 3957 13642
rect 3991 13608 4029 13642
rect 4063 13608 4101 13642
rect 4135 13608 4173 13642
rect 4207 13608 4245 13642
rect 4279 13608 4317 13642
rect 4351 13608 4389 13642
rect 4423 13608 4461 13642
rect 4495 13608 4533 13642
rect 4567 13608 4605 13642
rect 4639 13608 12900 13642
rect 2221 13544 2225 13593
rect 2395 13544 2399 13593
rect 2395 11095 2399 11134
rect 2221 11023 2225 11062
rect 2395 11022 2399 11061
rect 2221 10950 2225 10989
rect 2395 10949 2399 10988
rect 2221 10877 2225 10916
rect 2395 10876 2399 10915
rect 2221 10804 2225 10843
rect 2395 10803 2399 10842
rect 2221 10731 2225 10770
rect 2395 10730 2399 10769
rect 2221 10658 2225 10697
rect 2395 10657 2399 10696
rect 2221 10585 2225 10624
rect 2395 10584 2399 10623
rect 2221 10512 2225 10551
rect 2395 10511 2399 10550
rect 2221 10439 2225 10478
rect 2395 10438 2399 10477
rect 2221 10366 2225 10405
rect 2395 10365 2399 10404
rect 2221 10293 2225 10332
rect 2395 10292 2399 10331
rect 2221 10220 2225 10259
rect 2395 10219 2399 10258
rect 2221 10147 2225 10186
rect 2395 10146 2399 10185
rect 2221 10074 2225 10113
rect 2395 10073 2399 10112
rect 2221 10001 2225 10040
rect 2395 10000 2399 10039
rect 2221 9928 2225 9967
rect 2395 9927 2399 9966
rect 2221 9855 2225 9894
rect 2395 9854 2399 9893
rect 2221 9782 2225 9821
rect 2395 9781 2399 9820
rect 2221 9709 2225 9748
rect 2395 9708 2399 9747
rect 2221 9636 2225 9675
rect 2395 9635 2399 9674
rect 2221 9563 2225 9602
rect 2395 9562 2399 9601
rect 2221 9490 2225 9529
rect 2395 9489 2399 9528
rect 2221 9417 2225 9456
rect 2395 9416 2399 9455
rect 2221 9344 2225 9383
rect 2395 9343 2399 9382
rect 2617 13521 2651 13559
rect 2617 13449 2651 13487
rect 3141 13508 12900 13608
rect 3141 13474 3176 13508
rect 3210 13474 3244 13508
rect 3278 13474 3578 13508
rect 3612 13474 3646 13508
rect 3680 13474 4096 13508
rect 4130 13474 4164 13508
rect 4198 13474 4498 13508
rect 4532 13474 4566 13508
rect 4600 13474 5016 13508
rect 5050 13474 5084 13508
rect 5118 13474 5418 13508
rect 5452 13474 5486 13508
rect 5520 13474 5936 13508
rect 5970 13474 6004 13508
rect 6038 13474 6338 13508
rect 6372 13474 6406 13508
rect 6440 13474 6856 13508
rect 6890 13474 6924 13508
rect 6958 13474 7258 13508
rect 7292 13474 7326 13508
rect 7360 13474 7776 13508
rect 7810 13474 7844 13508
rect 7878 13474 8178 13508
rect 8212 13474 8246 13508
rect 8280 13474 8696 13508
rect 8730 13474 8764 13508
rect 8798 13474 9098 13508
rect 9132 13474 9166 13508
rect 9200 13474 9616 13508
rect 9650 13474 9684 13508
rect 9718 13474 10018 13508
rect 10052 13474 10086 13508
rect 10120 13474 10536 13508
rect 10570 13474 10604 13508
rect 10638 13474 10938 13508
rect 10972 13474 11006 13508
rect 11040 13474 11456 13508
rect 11490 13474 11524 13508
rect 11558 13474 11858 13508
rect 11892 13474 11926 13508
rect 11960 13474 12376 13508
rect 12410 13474 12444 13508
rect 12478 13474 12778 13508
rect 12812 13474 12846 13508
rect 12880 13474 12900 13508
rect 3141 13468 12900 13474
rect 2617 13377 2651 13415
rect 2617 13305 2651 13343
rect 2617 13233 2651 13271
rect 2617 13161 2651 13199
rect 2617 13089 2651 13127
rect 2617 13017 2651 13055
rect 2617 12945 2651 12983
rect 2617 12873 2651 12911
rect 2617 12801 2651 12839
rect 2617 12729 2651 12767
rect 2617 12657 2651 12695
rect 2617 12585 2651 12623
rect 2617 12513 2651 12551
rect 2617 12441 2651 12479
rect 2617 12369 2651 12407
rect 2617 12297 2651 12335
rect 2617 12225 2651 12263
rect 2617 12153 2651 12191
rect 2617 12081 2651 12119
rect 2617 12009 2651 12047
rect 2617 11937 2651 11975
rect 2617 11865 2651 11903
rect 2617 11793 2651 11831
rect 2617 11721 2651 11759
rect 2617 11649 2651 11687
rect 2617 11577 2651 11615
rect 2617 11505 2651 11543
rect 2617 11433 2651 11471
rect 2617 11361 2651 11399
rect 2617 11289 2651 11327
rect 2617 11217 2651 11255
rect 2617 11145 2651 11183
rect 2617 11073 2651 11111
rect 2617 11001 2651 11039
rect 2617 10929 2651 10967
rect 2617 10857 2651 10895
rect 2617 10784 2651 10823
rect 2617 10711 2651 10750
rect 2617 10638 2651 10677
rect 2617 10565 2651 10604
rect 2617 10492 2651 10531
rect 2617 10419 2651 10458
rect 2617 10346 2651 10385
rect 2617 10273 2651 10312
rect 2617 10200 2651 10239
rect 2617 10127 2651 10166
rect 2617 10054 2651 10093
rect 2617 9981 2651 10020
rect 2617 9908 2651 9947
rect 2617 9835 2651 9874
rect 2617 9762 2651 9801
rect 2617 9689 2651 9728
rect 2617 9616 2651 9655
rect 2617 9543 2651 9582
rect 2617 9470 2651 9509
rect 2617 9398 2651 9436
rect 2877 13371 3083 13386
rect 3055 10817 3083 13371
rect 2877 10778 3083 10817
rect 2911 10744 2949 10778
rect 2983 10744 3021 10778
rect 3055 10744 3083 10778
rect 2877 10705 3083 10744
rect 2911 10671 2949 10705
rect 2983 10671 3021 10705
rect 3055 10671 3083 10705
rect 2877 10632 3083 10671
rect 2911 10598 2949 10632
rect 2983 10598 3021 10632
rect 3055 10598 3083 10632
rect 2877 10559 3083 10598
rect 2911 10525 2949 10559
rect 2983 10525 3021 10559
rect 3055 10525 3083 10559
rect 2877 10486 3083 10525
rect 2911 10452 2949 10486
rect 2983 10452 3021 10486
rect 3055 10452 3083 10486
rect 2877 10413 3083 10452
rect 2911 10379 2949 10413
rect 2983 10379 3021 10413
rect 3055 10379 3083 10413
rect 2877 10340 3083 10379
rect 2911 10306 2949 10340
rect 2983 10306 3021 10340
rect 3055 10306 3083 10340
rect 2877 10267 3083 10306
rect 2911 10233 2949 10267
rect 2983 10233 3021 10267
rect 3055 10233 3083 10267
rect 2877 10194 3083 10233
rect 2911 10160 2949 10194
rect 2983 10160 3021 10194
rect 3055 10160 3083 10194
rect 2877 10121 3083 10160
rect 2911 10087 2949 10121
rect 2983 10087 3021 10121
rect 3055 10087 3083 10121
rect 2877 10048 3083 10087
rect 2911 10014 2949 10048
rect 2983 10014 3021 10048
rect 3055 10014 3083 10048
rect 2877 9975 3083 10014
rect 2911 9941 2949 9975
rect 2983 9941 3021 9975
rect 3055 9941 3083 9975
rect 2877 9902 3083 9941
rect 2911 9868 2949 9902
rect 2983 9868 3021 9902
rect 3055 9868 3083 9902
rect 2877 9829 3083 9868
rect 2911 9795 2949 9829
rect 2983 9795 3021 9829
rect 3055 9795 3083 9829
rect 2877 9756 3083 9795
rect 2911 9722 2949 9756
rect 2983 9722 3021 9756
rect 3055 9722 3083 9756
rect 2877 9683 3083 9722
rect 2911 9649 2949 9683
rect 2983 9649 3021 9683
rect 3055 9649 3083 9683
rect 2877 9610 3083 9649
rect 2911 9576 2949 9610
rect 2983 9576 3021 9610
rect 3055 9576 3083 9610
rect 2877 9537 3083 9576
rect 2911 9503 2949 9537
rect 2983 9503 3021 9537
rect 3055 9503 3083 9537
rect 12969 13362 13175 13386
rect 3797 10778 3975 10817
rect 3831 10744 3869 10778
rect 3903 10744 3941 10778
rect 3797 10705 3975 10744
rect 3831 10671 3869 10705
rect 3903 10671 3941 10705
rect 3797 10632 3975 10671
rect 3831 10598 3869 10632
rect 3903 10598 3941 10632
rect 3797 10559 3975 10598
rect 3831 10525 3869 10559
rect 3903 10525 3941 10559
rect 3797 10486 3975 10525
rect 3831 10452 3869 10486
rect 3903 10452 3941 10486
rect 3797 10413 3975 10452
rect 3831 10379 3869 10413
rect 3903 10379 3941 10413
rect 3797 10340 3975 10379
rect 3831 10306 3869 10340
rect 3903 10306 3941 10340
rect 3797 10267 3975 10306
rect 3831 10233 3869 10267
rect 3903 10233 3941 10267
rect 3797 10194 3975 10233
rect 3831 10160 3869 10194
rect 3903 10160 3941 10194
rect 3797 10121 3975 10160
rect 3831 10087 3869 10121
rect 3903 10087 3941 10121
rect 3797 10048 3975 10087
rect 3831 10014 3869 10048
rect 3903 10014 3941 10048
rect 3797 9975 3975 10014
rect 3831 9941 3869 9975
rect 3903 9941 3941 9975
rect 3797 9902 3975 9941
rect 3831 9868 3869 9902
rect 3903 9868 3941 9902
rect 3797 9829 3975 9868
rect 3831 9795 3869 9829
rect 3903 9795 3941 9829
rect 3797 9756 3975 9795
rect 3831 9722 3869 9756
rect 3903 9722 3941 9756
rect 3797 9683 3975 9722
rect 3831 9649 3869 9683
rect 3903 9649 3941 9683
rect 3797 9610 3975 9649
rect 3831 9576 3869 9610
rect 3903 9576 3941 9610
rect 3797 9537 3975 9576
rect 3831 9503 3869 9537
rect 3903 9503 3941 9537
rect 4717 10121 4895 10160
rect 4751 10087 4789 10121
rect 4823 10087 4861 10121
rect 4717 10048 4895 10087
rect 4751 10014 4789 10048
rect 4823 10014 4861 10048
rect 4717 9975 4895 10014
rect 4751 9941 4789 9975
rect 4823 9941 4861 9975
rect 4717 9902 4895 9941
rect 4751 9868 4789 9902
rect 4823 9868 4861 9902
rect 4717 9829 4895 9868
rect 4751 9795 4789 9829
rect 4823 9795 4861 9829
rect 4717 9756 4895 9795
rect 4751 9722 4789 9756
rect 4823 9722 4861 9756
rect 4717 9683 4895 9722
rect 4751 9649 4789 9683
rect 4823 9649 4861 9683
rect 4717 9610 4895 9649
rect 4751 9576 4789 9610
rect 4823 9576 4861 9610
rect 4717 9537 4895 9576
rect 4751 9503 4789 9537
rect 4823 9503 4861 9537
rect 5637 10121 5815 10160
rect 5671 10087 5709 10121
rect 5743 10087 5781 10121
rect 5637 10048 5815 10087
rect 5671 10014 5709 10048
rect 5743 10014 5781 10048
rect 5637 9975 5815 10014
rect 5671 9941 5709 9975
rect 5743 9941 5781 9975
rect 5637 9902 5815 9941
rect 5671 9868 5709 9902
rect 5743 9868 5781 9902
rect 5637 9829 5815 9868
rect 5671 9795 5709 9829
rect 5743 9795 5781 9829
rect 5637 9756 5815 9795
rect 5671 9722 5709 9756
rect 5743 9722 5781 9756
rect 5637 9683 5815 9722
rect 5671 9649 5709 9683
rect 5743 9649 5781 9683
rect 5637 9610 5815 9649
rect 5671 9576 5709 9610
rect 5743 9576 5781 9610
rect 5637 9537 5815 9576
rect 5671 9503 5709 9537
rect 5743 9503 5781 9537
rect 6557 10121 6735 10160
rect 6591 10087 6629 10121
rect 6663 10087 6701 10121
rect 6557 10048 6735 10087
rect 6591 10014 6629 10048
rect 6663 10014 6701 10048
rect 6557 9975 6735 10014
rect 6591 9941 6629 9975
rect 6663 9941 6701 9975
rect 6557 9902 6735 9941
rect 6591 9868 6629 9902
rect 6663 9868 6701 9902
rect 6557 9829 6735 9868
rect 6591 9795 6629 9829
rect 6663 9795 6701 9829
rect 6557 9756 6735 9795
rect 6591 9722 6629 9756
rect 6663 9722 6701 9756
rect 6557 9683 6735 9722
rect 6591 9649 6629 9683
rect 6663 9649 6701 9683
rect 6557 9610 6735 9649
rect 6591 9576 6629 9610
rect 6663 9576 6701 9610
rect 6557 9537 6735 9576
rect 6591 9503 6629 9537
rect 6663 9503 6701 9537
rect 7477 10121 7655 10160
rect 7511 10087 7549 10121
rect 7583 10087 7621 10121
rect 7477 10048 7655 10087
rect 7511 10014 7549 10048
rect 7583 10014 7621 10048
rect 7477 9975 7655 10014
rect 7511 9941 7549 9975
rect 7583 9941 7621 9975
rect 7477 9902 7655 9941
rect 7511 9868 7549 9902
rect 7583 9868 7621 9902
rect 7477 9829 7655 9868
rect 7511 9795 7549 9829
rect 7583 9795 7621 9829
rect 7477 9756 7655 9795
rect 7511 9722 7549 9756
rect 7583 9722 7621 9756
rect 7477 9683 7655 9722
rect 7511 9649 7549 9683
rect 7583 9649 7621 9683
rect 7477 9610 7655 9649
rect 7511 9576 7549 9610
rect 7583 9576 7621 9610
rect 7477 9537 7655 9576
rect 7511 9503 7549 9537
rect 7583 9503 7621 9537
rect 8397 10121 8575 10160
rect 8431 10087 8469 10121
rect 8503 10087 8541 10121
rect 8397 10048 8575 10087
rect 8431 10014 8469 10048
rect 8503 10014 8541 10048
rect 8397 9975 8575 10014
rect 8431 9941 8469 9975
rect 8503 9941 8541 9975
rect 8397 9902 8575 9941
rect 8431 9868 8469 9902
rect 8503 9868 8541 9902
rect 8397 9829 8575 9868
rect 8431 9795 8469 9829
rect 8503 9795 8541 9829
rect 8397 9756 8575 9795
rect 8431 9722 8469 9756
rect 8503 9722 8541 9756
rect 8397 9683 8575 9722
rect 8431 9649 8469 9683
rect 8503 9649 8541 9683
rect 8397 9610 8575 9649
rect 8431 9576 8469 9610
rect 8503 9576 8541 9610
rect 8397 9537 8575 9576
rect 8431 9503 8469 9537
rect 8503 9503 8541 9537
rect 9317 10121 9495 10160
rect 9351 10087 9389 10121
rect 9423 10087 9461 10121
rect 9317 10048 9495 10087
rect 9351 10014 9389 10048
rect 9423 10014 9461 10048
rect 9317 9975 9495 10014
rect 9351 9941 9389 9975
rect 9423 9941 9461 9975
rect 9317 9902 9495 9941
rect 9351 9868 9389 9902
rect 9423 9868 9461 9902
rect 9317 9829 9495 9868
rect 9351 9795 9389 9829
rect 9423 9795 9461 9829
rect 9317 9756 9495 9795
rect 9351 9722 9389 9756
rect 9423 9722 9461 9756
rect 9317 9683 9495 9722
rect 9351 9649 9389 9683
rect 9423 9649 9461 9683
rect 9317 9610 9495 9649
rect 9351 9576 9389 9610
rect 9423 9576 9461 9610
rect 9317 9537 9495 9576
rect 9351 9503 9389 9537
rect 9423 9503 9461 9537
rect 10237 10121 10415 10160
rect 10271 10087 10309 10121
rect 10343 10087 10381 10121
rect 10237 10048 10415 10087
rect 10271 10014 10309 10048
rect 10343 10014 10381 10048
rect 10237 9975 10415 10014
rect 10271 9941 10309 9975
rect 10343 9941 10381 9975
rect 10237 9902 10415 9941
rect 10271 9868 10309 9902
rect 10343 9868 10381 9902
rect 10237 9829 10415 9868
rect 10271 9795 10309 9829
rect 10343 9795 10381 9829
rect 10237 9756 10415 9795
rect 10271 9722 10309 9756
rect 10343 9722 10381 9756
rect 10237 9683 10415 9722
rect 10271 9649 10309 9683
rect 10343 9649 10381 9683
rect 10237 9610 10415 9649
rect 10271 9576 10309 9610
rect 10343 9576 10381 9610
rect 10237 9537 10415 9576
rect 10271 9503 10309 9537
rect 10343 9503 10381 9537
rect 11157 10121 11335 10160
rect 11191 10087 11229 10121
rect 11263 10087 11301 10121
rect 11157 10048 11335 10087
rect 11191 10014 11229 10048
rect 11263 10014 11301 10048
rect 11157 9975 11335 10014
rect 11191 9941 11229 9975
rect 11263 9941 11301 9975
rect 11157 9902 11335 9941
rect 11191 9868 11229 9902
rect 11263 9868 11301 9902
rect 11157 9829 11335 9868
rect 11191 9795 11229 9829
rect 11263 9795 11301 9829
rect 11157 9756 11335 9795
rect 11191 9722 11229 9756
rect 11263 9722 11301 9756
rect 11157 9683 11335 9722
rect 11191 9649 11229 9683
rect 11263 9649 11301 9683
rect 11157 9610 11335 9649
rect 11191 9576 11229 9610
rect 11263 9576 11301 9610
rect 11157 9537 11335 9576
rect 11191 9503 11229 9537
rect 11263 9503 11301 9537
rect 12077 10121 12255 10160
rect 12111 10087 12149 10121
rect 12183 10087 12221 10121
rect 12077 10048 12255 10087
rect 12111 10014 12149 10048
rect 12183 10014 12221 10048
rect 12077 9975 12255 10014
rect 12111 9941 12149 9975
rect 12183 9941 12221 9975
rect 12077 9902 12255 9941
rect 12111 9868 12149 9902
rect 12183 9868 12221 9902
rect 12077 9829 12255 9868
rect 12111 9795 12149 9829
rect 12183 9795 12221 9829
rect 12077 9756 12255 9795
rect 12111 9722 12149 9756
rect 12183 9722 12221 9756
rect 12077 9683 12255 9722
rect 12111 9649 12149 9683
rect 12183 9649 12221 9683
rect 12077 9610 12255 9649
rect 12111 9576 12149 9610
rect 12183 9576 12221 9610
rect 12077 9537 12255 9576
rect 12111 9503 12149 9537
rect 12183 9503 12221 9537
rect 12969 10160 12997 13362
rect 12969 10121 13175 10160
rect 12969 10087 12997 10121
rect 13031 10087 13069 10121
rect 13103 10087 13141 10121
rect 12969 10048 13175 10087
rect 12969 10014 12997 10048
rect 13031 10014 13069 10048
rect 13103 10014 13141 10048
rect 12969 9975 13175 10014
rect 12969 9941 12997 9975
rect 13031 9941 13069 9975
rect 13103 9941 13141 9975
rect 12969 9902 13175 9941
rect 12969 9868 12997 9902
rect 13031 9868 13069 9902
rect 13103 9868 13141 9902
rect 12969 9829 13175 9868
rect 12969 9795 12997 9829
rect 13031 9795 13069 9829
rect 13103 9795 13141 9829
rect 12969 9756 13175 9795
rect 12969 9722 12997 9756
rect 13031 9722 13069 9756
rect 13103 9722 13141 9756
rect 12969 9683 13175 9722
rect 12969 9649 12997 9683
rect 13031 9649 13069 9683
rect 13103 9649 13141 9683
rect 12969 9610 13175 9649
rect 12969 9576 12997 9610
rect 13031 9576 13069 9610
rect 13103 9576 13141 9610
rect 12969 9537 13175 9576
rect 12969 9503 12997 9537
rect 13031 9503 13069 9537
rect 13103 9503 13141 9537
rect 2877 9432 3083 9503
rect 12969 9432 13175 9503
rect 2617 9397 3176 9398
rect 2651 9391 3176 9397
rect 3210 9391 3244 9398
rect 3278 9391 3578 9398
rect 3612 9391 3646 9398
rect 3680 9391 4096 9398
rect 4130 9391 4164 9398
rect 4198 9391 4498 9398
rect 4532 9391 4566 9398
rect 4600 9391 5016 9398
rect 5050 9391 5084 9398
rect 5118 9391 5418 9398
rect 5452 9391 5486 9398
rect 5520 9391 5936 9398
rect 5970 9391 6004 9398
rect 6038 9391 6338 9398
rect 2651 9363 2697 9391
rect 2618 9357 2697 9363
rect 2731 9357 2770 9391
rect 2804 9357 2843 9391
rect 2877 9357 2916 9391
rect 2950 9357 2989 9391
rect 3023 9357 3061 9391
rect 3095 9357 3133 9391
rect 3167 9364 3176 9391
rect 3239 9364 3244 9391
rect 3167 9357 3205 9364
rect 3239 9357 3277 9364
rect 3311 9357 3349 9391
rect 3383 9357 3421 9391
rect 3455 9357 3493 9391
rect 3527 9357 3565 9391
rect 3612 9364 3637 9391
rect 3680 9364 3709 9391
rect 3599 9357 3637 9364
rect 3671 9357 3709 9364
rect 3743 9357 3781 9391
rect 3815 9357 3853 9391
rect 3887 9357 3925 9391
rect 3959 9357 3997 9391
rect 4031 9357 4069 9391
rect 4130 9364 4141 9391
rect 4198 9364 4213 9391
rect 4103 9357 4141 9364
rect 4175 9357 4213 9364
rect 4247 9357 4285 9391
rect 4319 9357 4357 9391
rect 4391 9357 4429 9391
rect 4463 9364 4498 9391
rect 4535 9364 4566 9391
rect 4463 9357 4501 9364
rect 4535 9357 4573 9364
rect 4607 9357 4645 9391
rect 4679 9357 4717 9391
rect 4751 9357 4789 9391
rect 4823 9357 4861 9391
rect 4895 9357 4933 9391
rect 4967 9357 5005 9391
rect 5050 9364 5077 9391
rect 5118 9364 5149 9391
rect 5039 9357 5077 9364
rect 5111 9357 5149 9364
rect 5183 9357 5221 9391
rect 5255 9357 5293 9391
rect 5327 9357 5365 9391
rect 5399 9364 5418 9391
rect 5471 9364 5486 9391
rect 5399 9357 5437 9364
rect 5471 9357 5509 9364
rect 5543 9357 5581 9391
rect 5615 9357 5653 9391
rect 5687 9357 5725 9391
rect 5759 9357 5797 9391
rect 5831 9357 5869 9391
rect 5903 9364 5936 9391
rect 5975 9364 6004 9391
rect 5903 9357 5941 9364
rect 5975 9357 6013 9364
rect 6047 9357 6085 9391
rect 6119 9357 6157 9391
rect 6191 9357 6229 9391
rect 6263 9357 6301 9391
rect 6335 9364 6338 9391
rect 6372 9391 6406 9398
rect 6440 9391 6856 9398
rect 6890 9391 6924 9398
rect 6958 9391 7258 9398
rect 7292 9391 7326 9398
rect 7360 9391 7776 9398
rect 6372 9364 6373 9391
rect 6440 9364 6445 9391
rect 6335 9357 6373 9364
rect 6407 9357 6445 9364
rect 6479 9357 6517 9391
rect 6551 9357 6589 9391
rect 6623 9357 6661 9391
rect 6695 9357 6733 9391
rect 6767 9357 6805 9391
rect 6839 9364 6856 9391
rect 6911 9364 6924 9391
rect 6839 9357 6877 9364
rect 6911 9357 6949 9364
rect 6983 9357 7021 9391
rect 7055 9357 7093 9391
rect 7127 9357 7165 9391
rect 7199 9357 7237 9391
rect 7292 9364 7309 9391
rect 7360 9364 7381 9391
rect 7271 9357 7309 9364
rect 7343 9357 7381 9364
rect 7415 9357 7453 9391
rect 7487 9357 7525 9391
rect 7559 9357 7597 9391
rect 7631 9357 7669 9391
rect 7703 9357 7741 9391
rect 7775 9364 7776 9391
rect 7810 9391 7844 9398
rect 7878 9391 8178 9398
rect 8212 9391 8246 9398
rect 8280 9391 8696 9398
rect 8730 9391 8764 9398
rect 8798 9391 9098 9398
rect 9132 9391 9166 9398
rect 9200 9391 9616 9398
rect 7810 9364 7813 9391
rect 7878 9364 7885 9391
rect 7775 9357 7813 9364
rect 7847 9357 7885 9364
rect 7919 9357 7957 9391
rect 7991 9357 8029 9391
rect 8063 9357 8101 9391
rect 8135 9357 8173 9391
rect 8212 9364 8245 9391
rect 8280 9364 8317 9391
rect 8207 9357 8245 9364
rect 8279 9357 8317 9364
rect 8351 9357 8389 9391
rect 8423 9357 8461 9391
rect 8495 9357 8533 9391
rect 8567 9357 8605 9391
rect 8639 9357 8677 9391
rect 8730 9364 8749 9391
rect 8798 9364 8821 9391
rect 8711 9357 8749 9364
rect 8783 9357 8821 9364
rect 8855 9357 8893 9391
rect 8927 9357 8965 9391
rect 8999 9357 9037 9391
rect 9071 9364 9098 9391
rect 9143 9364 9166 9391
rect 9071 9357 9109 9364
rect 9143 9357 9181 9364
rect 9215 9357 9253 9391
rect 9287 9357 9325 9391
rect 9359 9357 9397 9391
rect 9431 9357 9469 9391
rect 9503 9357 9541 9391
rect 9575 9357 9613 9391
rect 9650 9364 9684 9398
rect 9718 9391 10018 9398
rect 10052 9391 10086 9398
rect 10120 9391 10536 9398
rect 10570 9391 10604 9398
rect 10638 9391 10938 9398
rect 10972 9391 11006 9398
rect 11040 9391 11456 9398
rect 11490 9391 11524 9398
rect 11558 9391 11858 9398
rect 11892 9391 11926 9398
rect 11960 9391 12376 9398
rect 12410 9391 12444 9398
rect 12478 9391 12778 9398
rect 12812 9391 12846 9398
rect 12880 9391 12900 9398
rect 9647 9357 9685 9364
rect 9719 9357 9757 9391
rect 9791 9357 9829 9391
rect 9863 9357 9901 9391
rect 9935 9357 9973 9391
rect 10007 9364 10018 9391
rect 10079 9364 10086 9391
rect 10007 9357 10045 9364
rect 10079 9357 10117 9364
rect 10151 9357 10189 9391
rect 10223 9357 10261 9391
rect 10295 9357 10333 9391
rect 10367 9357 10405 9391
rect 10439 9357 10477 9391
rect 10511 9364 10536 9391
rect 10583 9364 10604 9391
rect 10511 9357 10549 9364
rect 10583 9357 10621 9364
rect 10655 9357 10693 9391
rect 10727 9357 10765 9391
rect 10799 9357 10837 9391
rect 10871 9357 10909 9391
rect 10972 9364 10981 9391
rect 11040 9364 11053 9391
rect 10943 9357 10981 9364
rect 11015 9357 11053 9364
rect 11087 9357 11125 9391
rect 11159 9357 11197 9391
rect 11231 9357 11269 9391
rect 11303 9357 11341 9391
rect 11375 9357 11413 9391
rect 11447 9364 11456 9391
rect 11519 9364 11524 9391
rect 11447 9357 11485 9364
rect 11519 9357 11557 9364
rect 11591 9357 11629 9391
rect 11663 9357 11701 9391
rect 11735 9357 11773 9391
rect 11807 9357 11845 9391
rect 11892 9364 11917 9391
rect 11960 9364 11989 9391
rect 11879 9357 11917 9364
rect 11951 9357 11989 9364
rect 12023 9357 12061 9391
rect 12095 9357 12133 9391
rect 12167 9357 12205 9391
rect 12239 9357 12277 9391
rect 12311 9357 12349 9391
rect 12410 9364 12421 9391
rect 12478 9364 12493 9391
rect 12383 9357 12421 9364
rect 12455 9357 12493 9364
rect 12527 9357 12565 9391
rect 12599 9357 12637 9391
rect 12671 9357 12709 9391
rect 12743 9364 12778 9391
rect 12815 9364 12846 9391
rect 12743 9357 12781 9364
rect 12815 9357 12853 9364
rect 12887 9357 12900 9391
rect 2618 9348 12900 9357
rect 2221 9271 2225 9310
rect 2327 9309 2365 9313
rect 2327 9270 2399 9309
rect 2327 9266 2365 9270
rect 2255 9237 2293 9245
rect 2327 9237 2361 9266
rect 2221 9211 2361 9237
rect 2221 9198 2225 9211
rect 2259 9198 2361 9211
rect 2259 9177 2293 9198
rect 2255 9164 2293 9177
rect 2221 9092 2293 9164
rect 13559 9092 13631 9164
rect 13775 9116 13781 9165
rect 14019 9121 14025 9165
rect 2072 9024 2077 9063
rect 1827 8953 1834 8992
rect 2005 8991 2043 9012
rect 2004 8990 2043 8991
rect 2004 8952 2077 8990
rect 2005 8951 2077 8952
rect 13775 9033 13781 9082
rect 14019 9043 14025 9087
rect 13775 8951 13781 8999
rect 14019 8966 14025 9009
rect 1827 8880 1834 8919
rect 1936 8918 1971 8944
rect 2005 8940 2043 8951
rect 8845 8940 8884 8951
rect 8918 8940 8957 8951
rect 8991 8940 9030 8951
rect 9064 8940 9103 8951
rect 9137 8940 9176 8951
rect 9210 8940 9249 8951
rect 9283 8940 9322 8951
rect 9356 8940 9395 8951
rect 9429 8940 9468 8951
rect 9502 8940 9541 8951
rect 9575 8940 9614 8951
rect 9648 8940 9687 8951
rect 9721 8940 9760 8951
rect 9794 8940 9833 8951
rect 9867 8940 9906 8951
rect 9940 8940 9979 8951
rect 10013 8940 10052 8951
rect 10086 8940 10125 8951
rect 10159 8940 10198 8951
rect 10232 8940 10271 8951
rect 10305 8940 10344 8951
rect 10378 8940 10417 8951
rect 10451 8940 10490 8951
rect 10524 8940 10563 8951
rect 10597 8940 10636 8951
rect 10670 8940 10709 8951
rect 10743 8940 10782 8951
rect 10816 8940 10855 8951
rect 10889 8940 10928 8951
rect 10962 8940 11001 8951
rect 11035 8940 11074 8951
rect 11108 8940 11147 8951
rect 11181 8940 11220 8951
rect 11254 8940 11293 8951
rect 11327 8940 11366 8951
rect 11400 8940 11439 8951
rect 11473 8940 11512 8951
rect 11546 8940 11585 8951
rect 11619 8940 11658 8951
rect 11692 8940 11731 8951
rect 11765 8940 11804 8951
rect 11838 8940 11877 8951
rect 11911 8940 11950 8951
rect 11984 8940 12023 8951
rect 12057 8940 12096 8951
rect 12130 8940 12169 8951
rect 12203 8940 12242 8951
rect 12276 8940 12315 8951
rect 12349 8940 12388 8951
rect 12422 8940 12461 8951
rect 12495 8940 12534 8951
rect 12568 8940 12607 8951
rect 12641 8940 12680 8951
rect 12714 8940 12753 8951
rect 12787 8940 12826 8951
rect 12860 8940 12899 8951
rect 12933 8940 12972 8951
rect 13006 8940 13045 8951
rect 13079 8940 13118 8951
rect 13152 8940 13191 8951
rect 13225 8940 13264 8951
rect 13298 8940 13337 8951
rect 13371 8940 13410 8951
rect 13444 8940 13483 8951
rect 13517 8940 13556 8951
rect 13590 8940 13629 8951
rect 13663 8940 13702 8951
rect 2005 8918 2038 8940
rect 1936 8879 2038 8918
rect 13700 8917 13702 8940
rect 13736 8917 13775 8951
rect 13700 8906 13781 8917
rect 13700 8879 13849 8906
rect 14019 8889 14025 8932
rect 1936 8876 1971 8879
rect 1861 8846 1899 8876
rect 1933 8872 1971 8876
rect 1933 8846 1970 8872
rect 1827 8842 1970 8846
rect 1827 8808 1834 8842
rect 1868 8808 1970 8842
rect 1827 8807 1970 8808
rect 13700 8872 13701 8879
rect 13735 8872 13774 8879
rect 13768 8845 13774 8872
rect 13808 8845 13847 8879
rect 13768 8838 13849 8845
rect 13768 8807 13917 8838
rect 14019 8812 14025 8855
rect 1861 8773 1899 8807
rect 229 8690 263 8728
rect 1827 8701 1899 8773
rect 13768 8804 13773 8807
rect 13807 8804 13846 8807
rect 13836 8773 13846 8804
rect 13880 8773 13917 8807
rect 13836 8770 13917 8773
rect 14019 8770 14025 8778
rect 13836 8736 14025 8770
rect 13836 8735 13870 8736
rect 13904 8735 14025 8736
rect 13836 8702 13846 8735
rect 13904 8702 13919 8735
rect 8989 8701 9028 8702
rect 9062 8701 9101 8702
rect 9135 8701 9174 8702
rect 9208 8701 9247 8702
rect 9281 8701 9320 8702
rect 9354 8701 9393 8702
rect 9427 8701 9466 8702
rect 9500 8701 9539 8702
rect 9573 8701 9612 8702
rect 9646 8701 9685 8702
rect 9719 8701 9758 8702
rect 9792 8701 9831 8702
rect 9865 8701 9904 8702
rect 9938 8701 9977 8702
rect 10011 8701 10050 8702
rect 10084 8701 10123 8702
rect 10157 8701 10196 8702
rect 10230 8701 10269 8702
rect 10303 8701 10342 8702
rect 10376 8701 10415 8702
rect 10449 8701 10488 8702
rect 10522 8701 10561 8702
rect 10595 8701 10634 8702
rect 10668 8701 10707 8702
rect 10741 8701 10780 8702
rect 10814 8701 10853 8702
rect 10887 8701 10926 8702
rect 10960 8701 10999 8702
rect 11033 8701 11072 8702
rect 11106 8701 11145 8702
rect 11179 8701 11218 8702
rect 11252 8701 11291 8702
rect 11325 8701 11364 8702
rect 11398 8701 11437 8702
rect 11471 8701 11510 8702
rect 11544 8701 11583 8702
rect 11617 8701 11656 8702
rect 11690 8701 11729 8702
rect 11763 8701 11802 8702
rect 11836 8701 11875 8702
rect 11909 8701 11948 8702
rect 11982 8701 12021 8702
rect 12055 8701 12094 8702
rect 12128 8701 12167 8702
rect 12201 8701 12240 8702
rect 12274 8701 12313 8702
rect 12347 8701 12386 8702
rect 12420 8701 12459 8702
rect 12493 8701 12532 8702
rect 12566 8701 12605 8702
rect 12639 8701 12678 8702
rect 12712 8701 12751 8702
rect 12785 8701 12824 8702
rect 12858 8701 12897 8702
rect 12931 8701 12970 8702
rect 13004 8701 13043 8702
rect 13077 8701 13116 8702
rect 13150 8701 13189 8702
rect 13223 8701 13262 8702
rect 13296 8701 13335 8702
rect 13369 8701 13408 8702
rect 13442 8701 13481 8702
rect 13515 8701 13554 8702
rect 13588 8701 13627 8702
rect 13661 8701 13700 8702
rect 13734 8701 13773 8702
rect 13807 8701 13846 8702
rect 13880 8701 13919 8702
rect 13953 8701 14025 8735
rect 1644 8654 1682 8688
rect 14128 8564 14166 8598
rect 14200 8564 14211 8598
rect 14145 8547 14211 8564
rect 10464 8465 10536 8499
rect 10570 8465 10609 8499
rect 10643 8465 10682 8499
rect 10716 8465 10755 8499
rect 10789 8465 10828 8499
rect 10862 8465 10901 8499
rect 10935 8465 10974 8499
rect 11008 8465 11047 8499
rect 11081 8465 11120 8499
rect 11154 8465 11193 8499
rect 11227 8465 11266 8499
rect 11300 8465 11339 8499
rect 11373 8465 11412 8499
rect 11446 8465 11485 8499
rect 11519 8465 11558 8499
rect 11592 8465 11631 8499
rect 11665 8465 11704 8499
rect 11738 8465 11777 8499
rect 11811 8465 11850 8499
rect 11884 8465 11923 8499
rect 11957 8465 11996 8499
rect 12030 8465 12069 8499
rect 12103 8465 12142 8499
rect 12176 8465 12215 8499
rect 12249 8465 12288 8499
rect 12322 8465 12361 8499
rect 12395 8465 12434 8499
rect 12468 8465 12507 8499
rect 12541 8465 12580 8499
rect 12614 8465 12653 8499
rect 12687 8465 12726 8499
rect 12760 8465 12799 8499
rect 12833 8465 12872 8499
rect 12906 8465 12945 8499
rect 12979 8465 13018 8499
rect 13052 8465 13091 8499
rect 10464 8457 13091 8465
rect 10464 8427 10604 8457
rect 10638 8427 10672 8457
rect 10706 8427 10740 8457
rect 10774 8427 10808 8457
rect 10842 8427 10876 8457
rect 10910 8427 10944 8457
rect 10978 8427 11012 8457
rect 10464 8426 10536 8427
rect 10498 8393 10536 8426
rect 10570 8423 10604 8427
rect 10643 8423 10672 8427
rect 10716 8423 10740 8427
rect 10789 8423 10808 8427
rect 10862 8423 10876 8427
rect 10935 8423 10944 8427
rect 11008 8423 11012 8427
rect 11046 8427 11080 8457
rect 11114 8427 11148 8457
rect 11182 8427 11216 8457
rect 11250 8427 11284 8457
rect 11318 8427 11352 8457
rect 11386 8427 11420 8457
rect 11454 8427 11488 8457
rect 11046 8423 11047 8427
rect 11114 8423 11120 8427
rect 11182 8423 11193 8427
rect 11250 8423 11266 8427
rect 11318 8423 11339 8427
rect 11386 8423 11412 8427
rect 11454 8423 11485 8427
rect 11522 8423 11556 8457
rect 11590 8427 11624 8457
rect 11658 8427 11692 8457
rect 11726 8427 11760 8457
rect 11794 8427 11828 8457
rect 11862 8427 11896 8457
rect 11930 8427 11964 8457
rect 11998 8427 12032 8457
rect 11592 8423 11624 8427
rect 11665 8423 11692 8427
rect 11738 8423 11760 8427
rect 11811 8423 11828 8427
rect 11884 8423 11896 8427
rect 11957 8423 11964 8427
rect 12030 8423 12032 8427
rect 12066 8427 12100 8457
rect 12134 8427 12168 8457
rect 12202 8427 12236 8457
rect 12270 8427 12304 8457
rect 12338 8427 12372 8457
rect 12406 8427 12440 8457
rect 12474 8427 12508 8457
rect 12066 8423 12069 8427
rect 12134 8423 12142 8427
rect 12202 8423 12215 8427
rect 12270 8423 12288 8427
rect 12338 8423 12361 8427
rect 12406 8423 12434 8427
rect 12474 8423 12507 8427
rect 12542 8423 12576 8457
rect 12610 8427 12644 8457
rect 12678 8427 12712 8457
rect 12746 8427 12780 8457
rect 12814 8427 12848 8457
rect 12882 8427 12916 8457
rect 12950 8427 12984 8457
rect 12614 8423 12644 8427
rect 12687 8423 12712 8427
rect 12760 8423 12780 8427
rect 12833 8423 12848 8427
rect 12906 8423 12916 8427
rect 12979 8423 12984 8427
rect 13018 8427 13052 8457
rect 10570 8393 10609 8423
rect 10643 8393 10682 8423
rect 10716 8393 10755 8423
rect 10789 8393 10828 8423
rect 10862 8393 10901 8423
rect 10935 8393 10974 8423
rect 11008 8393 11047 8423
rect 11081 8393 11120 8423
rect 11154 8393 11193 8423
rect 11227 8393 11266 8423
rect 11300 8393 11339 8423
rect 11373 8393 11412 8423
rect 11446 8393 11485 8423
rect 11519 8393 11558 8423
rect 11592 8393 11631 8423
rect 11665 8393 11704 8423
rect 11738 8393 11777 8423
rect 11811 8393 11850 8423
rect 11884 8393 11923 8423
rect 11957 8393 11996 8423
rect 12030 8393 12069 8423
rect 12103 8393 12142 8423
rect 12176 8393 12215 8423
rect 12249 8393 12288 8423
rect 12322 8393 12361 8423
rect 12395 8393 12434 8423
rect 12468 8393 12507 8423
rect 12541 8393 12580 8423
rect 12614 8393 12653 8423
rect 12687 8393 12726 8423
rect 12760 8393 12799 8423
rect 12833 8393 12872 8423
rect 12906 8393 12945 8423
rect 12979 8393 13018 8423
rect 13086 8423 13091 8457
rect 13701 8427 13773 8499
rect 13052 8393 13091 8423
rect 13701 8393 13739 8427
rect 10498 8392 13163 8393
rect 10464 8389 13163 8392
rect 10464 8355 10473 8389
rect 10507 8355 13163 8389
rect 10464 8353 10608 8355
rect 10498 8321 10536 8353
rect 10507 8319 10536 8321
rect 10570 8325 10608 8353
rect 10642 8325 10681 8355
rect 10715 8325 10754 8355
rect 10788 8325 10827 8355
rect 10861 8325 10900 8355
rect 10934 8325 10973 8355
rect 11007 8325 11046 8355
rect 11080 8325 11119 8355
rect 11153 8325 11192 8355
rect 11226 8325 11265 8355
rect 11299 8325 11338 8355
rect 11372 8325 11411 8355
rect 11445 8325 11484 8355
rect 11518 8325 11557 8355
rect 11591 8325 11630 8355
rect 11664 8325 11703 8355
rect 11737 8325 11776 8355
rect 11810 8325 11849 8355
rect 11883 8325 11922 8355
rect 11956 8325 11995 8355
rect 12029 8325 12068 8355
rect 12102 8325 12141 8355
rect 12175 8325 12214 8355
rect 12248 8325 12287 8355
rect 12321 8325 12360 8355
rect 12394 8325 12433 8355
rect 12467 8325 12506 8355
rect 12540 8325 12579 8355
rect 12613 8325 12652 8355
rect 12686 8325 12725 8355
rect 12759 8325 12798 8355
rect 12832 8325 12871 8355
rect 12905 8325 12944 8355
rect 12978 8325 13017 8355
rect 13051 8325 13090 8355
rect 10570 8319 10605 8325
rect 10642 8321 10676 8325
rect 10715 8321 10744 8325
rect 10788 8321 10812 8325
rect 10861 8321 10880 8325
rect 10934 8321 10948 8325
rect 11007 8321 11016 8325
rect 11080 8321 11084 8325
rect 10464 8287 10473 8319
rect 10507 8291 10605 8319
rect 10639 8291 10676 8321
rect 10710 8291 10744 8321
rect 10778 8291 10812 8321
rect 10846 8291 10880 8321
rect 10914 8291 10948 8321
rect 10982 8291 11016 8321
rect 11050 8291 11084 8321
rect 11118 8321 11119 8325
rect 11186 8321 11192 8325
rect 11254 8321 11265 8325
rect 11322 8321 11338 8325
rect 11390 8321 11411 8325
rect 11458 8321 11484 8325
rect 11526 8321 11557 8325
rect 11118 8291 11152 8321
rect 11186 8291 11220 8321
rect 11254 8291 11288 8321
rect 11322 8291 11356 8321
rect 11390 8291 11424 8321
rect 11458 8291 11492 8321
rect 11526 8291 11560 8321
rect 11594 8291 11628 8325
rect 11664 8321 11696 8325
rect 11737 8321 11764 8325
rect 11810 8321 11832 8325
rect 11883 8321 11900 8325
rect 11956 8321 11968 8325
rect 12029 8321 12036 8325
rect 12102 8321 12104 8325
rect 11662 8291 11696 8321
rect 11730 8291 11764 8321
rect 11798 8291 11832 8321
rect 11866 8291 11900 8321
rect 11934 8291 11968 8321
rect 12002 8291 12036 8321
rect 12070 8291 12104 8321
rect 12138 8321 12141 8325
rect 12206 8321 12214 8325
rect 12274 8321 12287 8325
rect 12342 8321 12360 8325
rect 12410 8321 12433 8325
rect 12478 8321 12506 8325
rect 12546 8321 12579 8325
rect 12138 8291 12172 8321
rect 12206 8291 12240 8321
rect 12274 8291 12308 8321
rect 12342 8291 12376 8321
rect 12410 8291 12444 8321
rect 12478 8291 12512 8321
rect 12546 8291 12580 8321
rect 12614 8291 12648 8325
rect 12686 8321 12716 8325
rect 12759 8321 12784 8325
rect 12832 8321 12852 8325
rect 12905 8321 12920 8325
rect 12978 8321 12988 8325
rect 13051 8321 13056 8325
rect 12682 8291 12716 8321
rect 12750 8291 12784 8321
rect 12818 8291 12852 8321
rect 12886 8291 12920 8321
rect 12954 8291 12988 8321
rect 13022 8291 13056 8321
rect 13124 8325 13163 8355
rect 13557 8326 13773 8393
rect 13557 8325 13595 8326
rect 13629 8325 13773 8326
rect 13090 8291 13124 8321
rect 13158 8321 13163 8325
rect 13158 8291 13192 8321
rect 13226 8291 13260 8321
rect 13294 8291 13328 8321
rect 13362 8291 13396 8321
rect 13430 8291 13464 8321
rect 13498 8291 13532 8321
rect 13566 8292 13595 8325
rect 13634 8324 13773 8325
rect 13634 8297 13732 8324
rect 13766 8297 13773 8324
rect 13566 8291 13600 8292
rect 13634 8291 13667 8297
rect 10507 8287 10642 8291
rect 10464 8282 10642 8287
rect 10464 8280 10608 8282
rect 10498 8253 10536 8280
rect 10507 8246 10536 8253
rect 10570 8257 10608 8280
rect 13595 8263 13667 8291
rect 13701 8290 13732 8297
rect 13701 8263 13739 8290
rect 10570 8246 10605 8257
rect 10464 8219 10473 8246
rect 10507 8223 10605 8246
rect 10639 8223 10642 8248
rect 10507 8219 10642 8223
rect 10464 8209 10642 8219
rect 10464 8207 10608 8209
rect 10498 8185 10536 8207
rect 10507 8173 10536 8185
rect 10570 8189 10608 8207
rect 10570 8173 10605 8189
rect 10464 8151 10473 8173
rect 10507 8155 10605 8173
rect 10639 8155 10642 8175
rect 10507 8151 10642 8155
rect 10464 8136 10642 8151
rect 10464 8134 10608 8136
rect 10498 8117 10536 8134
rect 10507 8100 10536 8117
rect 10570 8121 10608 8134
rect 10570 8100 10605 8121
rect 13600 8256 13766 8263
rect 13600 8252 13732 8256
rect 13634 8222 13732 8252
rect 13634 8218 13766 8222
rect 13600 8188 13766 8218
rect 13600 8184 13732 8188
rect 13634 8154 13732 8184
rect 13634 8150 13766 8154
rect 13600 8120 13766 8150
rect 13600 8116 13732 8120
rect 10464 8083 10473 8100
rect 10507 8087 10605 8100
rect 10639 8087 10642 8102
rect 10507 8083 10642 8087
rect 10464 8063 10642 8083
rect 10464 8061 10608 8063
rect 10498 8049 10536 8061
rect 10507 8027 10536 8049
rect 10570 8053 10608 8061
rect 10570 8027 10605 8053
rect 10464 8015 10473 8027
rect 10507 8019 10605 8027
rect 10639 8019 10642 8029
rect 10507 8015 10642 8019
rect 10464 7990 10642 8015
rect 10464 7988 10608 7990
rect 10498 7981 10536 7988
rect 10507 7954 10536 7981
rect 10570 7985 10608 7988
rect 10570 7954 10605 7985
rect 10464 7947 10473 7954
rect 10507 7951 10605 7954
rect 10639 7951 10642 7956
rect 10507 7947 10642 7951
rect 10464 7917 10642 7947
rect 626 7913 698 7917
rect 732 7913 771 7917
rect 805 7913 844 7917
rect 878 7913 917 7917
rect 951 7913 990 7917
rect 1024 7913 1063 7917
rect 1097 7913 1136 7917
rect 1170 7913 1209 7917
rect 1243 7913 1282 7917
rect 1316 7913 1355 7917
rect 1389 7913 1428 7917
rect 1462 7913 1501 7917
rect 1535 7913 1574 7917
rect 1608 7913 1647 7917
rect 1681 7913 1720 7917
rect 1754 7913 1793 7917
rect 1827 7913 1866 7917
rect 1900 7913 1939 7917
rect 1973 7913 2012 7917
rect 2046 7913 2085 7917
rect 2119 7913 2158 7917
rect 2192 7913 2231 7917
rect 2265 7913 2304 7917
rect 2338 7913 2377 7917
rect 2411 7913 2450 7917
rect 2484 7913 2523 7917
rect 2557 7913 2596 7917
rect 2630 7913 2669 7917
rect 2703 7913 2742 7917
rect 2776 7913 2815 7917
rect 2849 7913 2888 7917
rect 2922 7913 2961 7917
rect 2995 7913 3034 7917
rect 3068 7913 3107 7917
rect 3141 7913 3180 7917
rect 3214 7913 3253 7917
rect 3287 7913 3326 7917
rect 3360 7913 3399 7917
rect 3433 7913 3472 7917
rect 3506 7913 3545 7917
rect 3579 7913 3618 7917
rect 3652 7913 3691 7917
rect 3725 7913 3764 7917
rect 3798 7913 3837 7917
rect 3871 7913 3910 7917
rect 3944 7913 3983 7917
rect 4017 7913 4056 7917
rect 4090 7913 4129 7917
rect 4163 7913 4202 7917
rect 4236 7913 4275 7917
rect 4309 7913 4348 7917
rect 4382 7913 4421 7917
rect 4455 7913 4494 7917
rect 620 7879 694 7913
rect 732 7883 762 7913
rect 728 7879 762 7883
rect 620 7845 762 7879
rect 732 7811 762 7845
rect 9568 7845 9640 7917
rect 9568 7811 9606 7845
rect 732 7777 830 7811
rect 790 7773 830 7777
rect 804 7743 830 7773
rect 9500 7778 9640 7811
rect 9500 7771 9602 7778
rect 9636 7771 9640 7778
rect 9500 7743 9534 7771
rect 804 7739 843 7743
rect 877 7739 916 7743
rect 950 7739 989 7743
rect 1023 7739 1062 7743
rect 1096 7739 1135 7743
rect 1169 7739 1208 7743
rect 1242 7739 1281 7743
rect 1315 7739 1354 7743
rect 1388 7739 1427 7743
rect 1461 7739 1500 7743
rect 1534 7739 1573 7743
rect 1607 7739 1646 7743
rect 1680 7739 1719 7743
rect 1753 7739 1792 7743
rect 1826 7739 1865 7743
rect 1899 7739 1938 7743
rect 1972 7739 2011 7743
rect 2045 7739 2084 7743
rect 2118 7739 2157 7743
rect 2191 7739 2230 7743
rect 2264 7739 2303 7743
rect 2337 7739 2376 7743
rect 2410 7739 2449 7743
rect 2483 7739 2522 7743
rect 2556 7739 2595 7743
rect 2629 7739 2668 7743
rect 2702 7739 2741 7743
rect 2775 7739 2814 7743
rect 2848 7739 2887 7743
rect 2921 7739 2960 7743
rect 2994 7739 3033 7743
rect 3067 7739 3106 7743
rect 3140 7739 3179 7743
rect 3213 7739 3252 7743
rect 3286 7739 3325 7743
rect 3359 7739 3398 7743
rect 3432 7739 3471 7743
rect 3505 7739 3544 7743
rect 3578 7739 3617 7743
rect 3651 7739 3690 7743
rect 3724 7739 3763 7743
rect 3797 7739 3836 7743
rect 3870 7739 3909 7743
rect 3943 7739 3982 7743
rect 4016 7739 4055 7743
rect 4089 7739 4128 7743
rect 4162 7739 4201 7743
rect 4235 7739 4274 7743
rect 4308 7739 4347 7743
rect 4381 7739 4420 7743
rect 4454 7739 4493 7743
rect 4527 7739 4566 7743
rect 9496 7739 9534 7743
rect 9462 7737 9534 7739
rect 9568 7744 9602 7771
rect 9568 7737 9606 7744
rect 9462 7710 9640 7737
rect 9462 7699 9534 7710
rect 9496 7665 9534 7699
rect 9636 7697 9640 7710
rect 9462 7642 9534 7665
rect 9462 7625 9466 7642
rect 9636 7623 9640 7663
rect 9462 7551 9466 7591
rect 790 6044 804 6083
rect 790 5971 804 6010
rect 790 5898 804 5937
rect 790 5825 804 5864
rect 947 7485 1019 7519
rect 1053 7485 1059 7519
rect 1125 7485 1127 7519
rect 1161 7485 1163 7519
rect 1229 7485 1235 7519
rect 1297 7485 1307 7519
rect 1365 7485 1379 7519
rect 1433 7485 1451 7519
rect 1501 7485 1523 7519
rect 1569 7485 1595 7519
rect 1637 7485 1667 7519
rect 1705 7485 1739 7519
rect 1773 7485 1807 7519
rect 1845 7485 1875 7519
rect 1917 7485 1943 7519
rect 1989 7485 2011 7519
rect 2061 7485 2079 7519
rect 2133 7485 2147 7519
rect 2205 7485 2215 7519
rect 2277 7485 2283 7519
rect 2349 7485 2351 7519
rect 2385 7485 2387 7519
rect 2453 7485 2459 7519
rect 2521 7485 2531 7519
rect 2589 7485 2603 7519
rect 2657 7485 2675 7519
rect 2725 7485 2747 7519
rect 2793 7485 2819 7519
rect 2861 7485 2891 7519
rect 2929 7485 2963 7519
rect 2997 7485 3031 7519
rect 3069 7485 3099 7519
rect 3141 7485 3167 7519
rect 3213 7485 3235 7519
rect 3285 7485 3303 7519
rect 3357 7485 3371 7519
rect 3429 7485 3439 7519
rect 3501 7485 3507 7519
rect 3573 7485 3575 7519
rect 3609 7485 3611 7519
rect 3677 7485 3683 7519
rect 3745 7485 3755 7519
rect 3813 7485 3827 7519
rect 3881 7485 3899 7519
rect 3949 7485 3971 7519
rect 4017 7485 4043 7519
rect 4085 7485 4115 7519
rect 4153 7485 4187 7519
rect 4221 7485 4255 7519
rect 4293 7485 4323 7519
rect 4365 7485 4391 7519
rect 4437 7485 4459 7519
rect 4509 7485 4527 7519
rect 4581 7485 4595 7519
rect 4653 7485 4663 7519
rect 4725 7485 4731 7519
rect 4797 7485 4799 7519
rect 4833 7485 4835 7519
rect 4901 7485 4907 7519
rect 4969 7485 4979 7519
rect 5037 7485 5051 7519
rect 5105 7485 5123 7519
rect 5173 7485 5195 7519
rect 5241 7485 5267 7519
rect 5309 7485 5339 7519
rect 5377 7485 5411 7519
rect 5445 7485 5479 7519
rect 5517 7485 5547 7519
rect 5589 7485 5615 7519
rect 5661 7485 5683 7519
rect 5733 7485 5751 7519
rect 5805 7485 5819 7519
rect 5877 7485 5887 7519
rect 5949 7485 5955 7519
rect 6021 7485 6023 7519
rect 6057 7485 6059 7519
rect 6125 7485 6131 7519
rect 6193 7485 6203 7519
rect 6261 7485 6275 7519
rect 6329 7485 6347 7519
rect 6397 7485 6419 7519
rect 6465 7485 6491 7519
rect 6533 7485 6563 7519
rect 6601 7485 6635 7519
rect 6669 7485 6703 7519
rect 6741 7485 6771 7519
rect 6813 7485 6839 7519
rect 6885 7485 6907 7519
rect 6957 7485 6975 7519
rect 7029 7485 7043 7519
rect 7101 7485 7111 7519
rect 7173 7485 7179 7519
rect 7245 7485 7247 7519
rect 7281 7485 7283 7519
rect 7349 7485 7355 7519
rect 7417 7485 7427 7519
rect 7485 7485 7499 7519
rect 7553 7485 7571 7519
rect 7621 7485 7643 7519
rect 7689 7485 7715 7519
rect 7757 7485 7787 7519
rect 7825 7485 7859 7519
rect 7893 7485 7927 7519
rect 7965 7485 7995 7519
rect 8037 7485 8063 7519
rect 8109 7485 8131 7519
rect 8181 7485 8199 7519
rect 8253 7485 8267 7519
rect 8325 7485 8335 7519
rect 8397 7485 8403 7519
rect 8469 7485 8471 7519
rect 8505 7485 8507 7519
rect 8573 7485 8579 7519
rect 8641 7485 8651 7519
rect 8709 7485 8723 7519
rect 8777 7485 8795 7519
rect 8845 7485 8867 7519
rect 8913 7485 8939 7519
rect 8981 7485 9012 7519
rect 9049 7485 9083 7519
rect 9119 7485 9191 7519
rect 947 7451 981 7485
rect 9151 7450 9191 7485
rect 947 7383 981 7413
rect 1268 7428 1284 7446
rect 1318 7428 1353 7446
rect 1387 7428 1422 7446
rect 1456 7428 1491 7446
rect 1268 7394 1269 7428
rect 1318 7412 1342 7428
rect 1387 7412 1415 7428
rect 1456 7412 1488 7428
rect 1525 7412 1560 7446
rect 1594 7428 1629 7446
rect 1663 7428 1698 7446
rect 1732 7428 1767 7446
rect 1801 7428 1836 7446
rect 1870 7428 1905 7446
rect 1939 7428 1974 7446
rect 2008 7428 2043 7446
rect 2077 7428 2112 7446
rect 2146 7428 2181 7446
rect 1595 7412 1629 7428
rect 1668 7412 1698 7428
rect 1741 7412 1767 7428
rect 1814 7412 1836 7428
rect 1887 7412 1905 7428
rect 1960 7412 1974 7428
rect 2033 7412 2043 7428
rect 2106 7412 2112 7428
rect 2179 7412 2181 7428
rect 2215 7428 2250 7446
rect 2284 7428 2319 7446
rect 2353 7428 2388 7446
rect 2422 7428 2457 7446
rect 2491 7428 2526 7446
rect 2560 7428 2595 7446
rect 2629 7428 2664 7446
rect 2698 7428 2733 7446
rect 2215 7412 2218 7428
rect 2284 7412 2291 7428
rect 2353 7412 2364 7428
rect 2422 7412 2437 7428
rect 2491 7412 2510 7428
rect 2560 7412 2583 7428
rect 2629 7412 2656 7428
rect 2698 7412 2729 7428
rect 2767 7412 2802 7446
rect 2836 7412 2871 7446
rect 2905 7428 2940 7446
rect 2974 7428 3009 7446
rect 3043 7428 3078 7446
rect 3112 7428 3147 7446
rect 3181 7428 3216 7446
rect 3250 7428 3285 7446
rect 3319 7428 3354 7446
rect 3388 7428 3423 7446
rect 2909 7412 2940 7428
rect 2982 7412 3009 7428
rect 3055 7412 3078 7428
rect 3128 7412 3147 7428
rect 3201 7412 3216 7428
rect 3274 7412 3285 7428
rect 3347 7412 3354 7428
rect 3420 7412 3423 7428
rect 3457 7428 3492 7446
rect 3526 7428 3561 7446
rect 3595 7428 3630 7446
rect 3664 7428 3699 7446
rect 3733 7428 3768 7446
rect 3802 7428 3837 7446
rect 3871 7428 3906 7446
rect 3940 7428 3975 7446
rect 4009 7428 4044 7446
rect 3457 7412 3459 7428
rect 3526 7412 3532 7428
rect 3595 7412 3605 7428
rect 3664 7412 3678 7428
rect 3733 7412 3751 7428
rect 3802 7412 3824 7428
rect 3871 7412 3897 7428
rect 3940 7412 3970 7428
rect 4009 7412 4043 7428
rect 4078 7412 4113 7446
rect 4147 7428 4182 7446
rect 4216 7428 4251 7446
rect 4285 7428 4320 7446
rect 4354 7428 4389 7446
rect 4423 7428 4458 7446
rect 4492 7428 4527 7446
rect 4561 7428 4596 7446
rect 4630 7428 4665 7446
rect 4150 7412 4182 7428
rect 4223 7412 4251 7428
rect 4296 7412 4320 7428
rect 4369 7412 4389 7428
rect 4442 7412 4458 7428
rect 4515 7412 4527 7428
rect 4588 7412 4596 7428
rect 4661 7412 4665 7428
rect 4699 7428 4734 7446
rect 4699 7412 4700 7428
rect 1303 7394 1342 7412
rect 1376 7394 1415 7412
rect 1449 7394 1488 7412
rect 1522 7394 1561 7412
rect 1595 7394 1634 7412
rect 1668 7394 1707 7412
rect 1741 7394 1780 7412
rect 1814 7394 1853 7412
rect 1887 7394 1926 7412
rect 1960 7394 1999 7412
rect 2033 7394 2072 7412
rect 2106 7394 2145 7412
rect 2179 7394 2218 7412
rect 2252 7394 2291 7412
rect 2325 7394 2364 7412
rect 2398 7394 2437 7412
rect 2471 7394 2510 7412
rect 2544 7394 2583 7412
rect 2617 7394 2656 7412
rect 2690 7394 2729 7412
rect 2763 7394 2802 7412
rect 2836 7394 2875 7412
rect 2909 7394 2948 7412
rect 2982 7394 3021 7412
rect 3055 7394 3094 7412
rect 3128 7394 3167 7412
rect 3201 7394 3240 7412
rect 3274 7394 3313 7412
rect 3347 7394 3386 7412
rect 3420 7394 3459 7412
rect 3493 7394 3532 7412
rect 3566 7394 3605 7412
rect 3639 7394 3678 7412
rect 3712 7394 3751 7412
rect 3785 7394 3824 7412
rect 3858 7394 3897 7412
rect 3931 7394 3970 7412
rect 4004 7394 4043 7412
rect 4077 7394 4116 7412
rect 4150 7394 4189 7412
rect 4223 7394 4262 7412
rect 4296 7394 4335 7412
rect 4369 7394 4408 7412
rect 4442 7394 4481 7412
rect 4515 7394 4554 7412
rect 4588 7394 4627 7412
rect 4661 7394 4700 7412
rect 4768 7428 4803 7446
rect 4837 7428 4872 7446
rect 4906 7428 4941 7446
rect 4975 7428 5010 7446
rect 5044 7428 5079 7446
rect 5113 7428 5148 7446
rect 5182 7428 5217 7446
rect 5251 7428 5286 7446
rect 4768 7412 4773 7428
rect 4837 7412 4846 7428
rect 4906 7412 4919 7428
rect 4975 7412 4992 7428
rect 5044 7412 5065 7428
rect 5113 7412 5138 7428
rect 5182 7412 5211 7428
rect 5251 7412 5284 7428
rect 5320 7412 5355 7446
rect 5389 7428 5424 7446
rect 5458 7428 5493 7446
rect 5527 7428 5562 7446
rect 5596 7428 5630 7446
rect 5664 7428 5698 7446
rect 5732 7428 5766 7446
rect 5800 7428 5834 7446
rect 5391 7412 5424 7428
rect 5464 7412 5493 7428
rect 5537 7412 5562 7428
rect 5610 7412 5630 7428
rect 5683 7412 5698 7428
rect 5756 7412 5766 7428
rect 5829 7412 5834 7428
rect 5868 7428 5902 7446
rect 4734 7394 4773 7412
rect 4807 7394 4846 7412
rect 4880 7394 4919 7412
rect 4953 7394 4992 7412
rect 5026 7394 5065 7412
rect 5099 7394 5138 7412
rect 5172 7394 5211 7412
rect 5245 7394 5284 7412
rect 5318 7394 5357 7412
rect 5391 7394 5430 7412
rect 5464 7394 5503 7412
rect 5537 7394 5576 7412
rect 5610 7394 5649 7412
rect 5683 7394 5722 7412
rect 5756 7394 5795 7412
rect 5829 7394 5868 7412
rect 5936 7428 5970 7446
rect 6004 7428 6038 7446
rect 6072 7428 6106 7446
rect 6140 7428 6174 7446
rect 6208 7428 6242 7446
rect 6276 7428 6310 7446
rect 5936 7412 5941 7428
rect 6004 7412 6014 7428
rect 6072 7412 6087 7428
rect 6140 7412 6160 7428
rect 6208 7412 6233 7428
rect 6276 7412 6306 7428
rect 6344 7412 6378 7446
rect 6412 7428 6446 7446
rect 6480 7428 6514 7446
rect 6548 7428 6582 7446
rect 6616 7428 6650 7446
rect 6684 7428 6718 7446
rect 6752 7428 6786 7446
rect 6820 7428 6854 7446
rect 6888 7428 6922 7446
rect 6956 7428 6990 7446
rect 6413 7412 6446 7428
rect 6485 7412 6514 7428
rect 6557 7412 6582 7428
rect 6629 7412 6650 7428
rect 6701 7412 6718 7428
rect 6773 7412 6786 7428
rect 6845 7412 6854 7428
rect 6917 7412 6922 7428
rect 6989 7412 6990 7428
rect 7024 7428 7058 7446
rect 7092 7428 7126 7446
rect 7160 7428 7194 7446
rect 7228 7428 7262 7446
rect 7296 7428 7330 7446
rect 7364 7428 7398 7446
rect 7432 7428 7466 7446
rect 7500 7428 7534 7446
rect 7024 7412 7027 7428
rect 7092 7412 7099 7428
rect 7160 7412 7171 7428
rect 7228 7412 7243 7428
rect 7296 7412 7315 7428
rect 7364 7412 7387 7428
rect 7432 7412 7459 7428
rect 7500 7412 7531 7428
rect 7568 7412 7602 7446
rect 7636 7428 7670 7446
rect 7704 7428 7738 7446
rect 7772 7428 7806 7446
rect 7840 7428 7874 7446
rect 7908 7428 7942 7446
rect 7976 7428 8010 7446
rect 8044 7428 8078 7446
rect 8112 7428 8146 7446
rect 8180 7428 8214 7446
rect 7637 7412 7670 7428
rect 7709 7412 7738 7428
rect 7781 7412 7806 7428
rect 7853 7412 7874 7428
rect 7925 7412 7942 7428
rect 7997 7412 8010 7428
rect 8069 7412 8078 7428
rect 8141 7412 8146 7428
rect 8213 7412 8214 7428
rect 8248 7428 8282 7446
rect 8316 7428 8350 7446
rect 8384 7428 8418 7446
rect 8452 7428 8486 7446
rect 8520 7428 8554 7446
rect 8588 7428 8622 7446
rect 8656 7428 8690 7446
rect 8724 7428 8758 7446
rect 8248 7412 8251 7428
rect 8316 7412 8323 7428
rect 8384 7412 8395 7428
rect 8452 7412 8467 7428
rect 8520 7412 8539 7428
rect 8588 7412 8611 7428
rect 8656 7412 8683 7428
rect 8724 7412 8755 7428
rect 8792 7412 8826 7446
rect 8860 7428 8894 7446
rect 8928 7428 8962 7446
rect 8996 7428 9012 7446
rect 8861 7412 8894 7428
rect 8933 7412 8962 7428
rect 5902 7394 5941 7412
rect 5975 7394 6014 7412
rect 6048 7394 6087 7412
rect 6121 7394 6160 7412
rect 6194 7394 6233 7412
rect 6267 7394 6306 7412
rect 6340 7394 6379 7412
rect 6413 7394 6451 7412
rect 6485 7394 6523 7412
rect 6557 7394 6595 7412
rect 6629 7394 6667 7412
rect 6701 7394 6739 7412
rect 6773 7394 6811 7412
rect 6845 7394 6883 7412
rect 6917 7394 6955 7412
rect 6989 7394 7027 7412
rect 7061 7394 7099 7412
rect 7133 7394 7171 7412
rect 7205 7394 7243 7412
rect 7277 7394 7315 7412
rect 7349 7394 7387 7412
rect 7421 7394 7459 7412
rect 7493 7394 7531 7412
rect 7565 7394 7603 7412
rect 7637 7394 7675 7412
rect 7709 7394 7747 7412
rect 7781 7394 7819 7412
rect 7853 7394 7891 7412
rect 7925 7394 7963 7412
rect 7997 7394 8035 7412
rect 8069 7394 8107 7412
rect 8141 7394 8179 7412
rect 8213 7394 8251 7412
rect 8285 7394 8323 7412
rect 8357 7394 8395 7412
rect 8429 7394 8467 7412
rect 8501 7394 8539 7412
rect 8573 7394 8611 7412
rect 8645 7394 8683 7412
rect 8717 7394 8755 7412
rect 8789 7394 8827 7412
rect 8861 7394 8899 7412
rect 8933 7394 8971 7412
rect 9005 7394 9012 7428
rect 9185 7445 9191 7450
rect 9151 7411 9157 7416
rect 947 7315 981 7338
rect 9151 7382 9191 7411
rect 9185 7371 9191 7382
rect 9151 7337 9157 7348
rect 9151 7314 9191 7337
rect 947 7247 981 7263
rect 947 7179 981 7188
rect 947 7111 981 7113
rect 947 7072 981 7077
rect 947 6997 981 7009
rect 947 6922 981 6941
rect 947 6847 981 6873
rect 947 6772 981 6805
rect 947 6703 981 6737
rect 1223 7224 1257 7264
rect 1223 7150 1257 7190
rect 1223 7076 1257 7116
rect 1223 7002 1257 7042
rect 1223 6927 1257 6968
rect 1223 6852 1257 6893
rect 1223 6777 1257 6818
rect 1223 6702 1257 6743
rect 1535 7224 1569 7264
rect 1535 7150 1569 7190
rect 1535 7076 1569 7116
rect 1535 7001 1569 7042
rect 1535 6926 1569 6967
rect 1535 6851 1569 6892
rect 1535 6776 1569 6817
rect 1535 6701 1569 6742
rect 1847 7224 1881 7264
rect 1847 7150 1881 7190
rect 1847 7076 1881 7116
rect 1847 7002 1881 7042
rect 1847 6927 1881 6968
rect 1847 6852 1881 6893
rect 1847 6777 1881 6818
rect 1847 6702 1881 6743
rect 2159 7224 2193 7264
rect 2159 7150 2193 7190
rect 2159 7076 2193 7116
rect 2159 7001 2193 7042
rect 2159 6926 2193 6967
rect 2159 6851 2193 6892
rect 2159 6776 2193 6817
rect 2159 6701 2193 6742
rect 2471 7224 2505 7264
rect 2471 7150 2505 7190
rect 2471 7076 2505 7116
rect 2471 7002 2505 7042
rect 2471 6927 2505 6968
rect 2471 6852 2505 6893
rect 2471 6777 2505 6818
rect 2471 6702 2505 6743
rect 2783 7224 2817 7264
rect 2783 7150 2817 7190
rect 2783 7076 2817 7116
rect 2783 7001 2817 7042
rect 2783 6926 2817 6967
rect 2783 6851 2817 6892
rect 2783 6776 2817 6817
rect 2783 6701 2817 6742
rect 3095 7224 3129 7264
rect 3095 7150 3129 7190
rect 3095 7076 3129 7116
rect 3095 7002 3129 7042
rect 3095 6927 3129 6968
rect 3095 6852 3129 6893
rect 3095 6777 3129 6818
rect 3095 6702 3129 6743
rect 3407 7224 3441 7264
rect 3407 7150 3441 7190
rect 3407 7076 3441 7116
rect 3407 7001 3441 7042
rect 3407 6926 3441 6967
rect 3407 6851 3441 6892
rect 3407 6776 3441 6817
rect 3407 6701 3441 6742
rect 3719 7224 3753 7264
rect 3719 7150 3753 7190
rect 3719 7076 3753 7116
rect 3719 7002 3753 7042
rect 3719 6927 3753 6968
rect 3719 6852 3753 6893
rect 3719 6777 3753 6818
rect 3719 6702 3753 6743
rect 4031 7224 4065 7264
rect 4031 7150 4065 7190
rect 4031 7076 4065 7116
rect 4031 7001 4065 7042
rect 4031 6926 4065 6967
rect 4031 6851 4065 6892
rect 4031 6776 4065 6817
rect 4031 6701 4065 6742
rect 4343 7224 4377 7264
rect 4343 7150 4377 7190
rect 4343 7076 4377 7116
rect 4343 7002 4377 7042
rect 4343 6927 4377 6968
rect 4343 6852 4377 6893
rect 4343 6777 4377 6818
rect 4343 6702 4377 6743
rect 4655 7224 4689 7264
rect 4655 7150 4689 7190
rect 4655 7076 4689 7116
rect 4655 7001 4689 7042
rect 4655 6926 4689 6967
rect 4655 6851 4689 6892
rect 4655 6776 4689 6817
rect 4655 6701 4689 6742
rect 4967 7224 5001 7264
rect 4967 7150 5001 7190
rect 4967 7076 5001 7116
rect 4967 7002 5001 7042
rect 4967 6927 5001 6968
rect 4967 6852 5001 6893
rect 4967 6777 5001 6818
rect 4967 6702 5001 6743
rect 5279 7224 5313 7264
rect 5279 7150 5313 7190
rect 5279 7076 5313 7116
rect 5279 7001 5313 7042
rect 5279 6926 5313 6967
rect 5279 6851 5313 6892
rect 5279 6776 5313 6817
rect 5279 6701 5313 6742
rect 5591 7224 5625 7264
rect 5591 7150 5625 7190
rect 5591 7076 5625 7116
rect 5591 7002 5625 7042
rect 5591 6927 5625 6968
rect 5591 6852 5625 6893
rect 5591 6777 5625 6818
rect 5591 6702 5625 6743
rect 5903 7224 5937 7264
rect 5903 7150 5937 7190
rect 5903 7076 5937 7116
rect 5903 7001 5937 7042
rect 5903 6926 5937 6967
rect 5903 6851 5937 6892
rect 5903 6776 5937 6817
rect 5903 6701 5937 6742
rect 6215 7224 6249 7264
rect 6215 7150 6249 7190
rect 6215 7076 6249 7116
rect 6215 7002 6249 7042
rect 6215 6927 6249 6968
rect 6215 6852 6249 6893
rect 6215 6777 6249 6818
rect 6215 6702 6249 6743
rect 6527 7224 6561 7264
rect 6527 7150 6561 7190
rect 6527 7076 6561 7116
rect 6527 7001 6561 7042
rect 6527 6926 6561 6967
rect 6527 6851 6561 6892
rect 6527 6776 6561 6817
rect 6527 6701 6561 6742
rect 6839 7224 6873 7264
rect 6839 7150 6873 7190
rect 6839 7076 6873 7116
rect 6839 7002 6873 7042
rect 6839 6927 6873 6968
rect 6839 6852 6873 6893
rect 6839 6777 6873 6818
rect 6839 6702 6873 6743
rect 7151 7224 7185 7264
rect 7151 7150 7185 7190
rect 7151 7076 7185 7116
rect 7151 7001 7185 7042
rect 7151 6926 7185 6967
rect 7151 6851 7185 6892
rect 7151 6776 7185 6817
rect 7151 6701 7185 6742
rect 7463 7224 7497 7264
rect 7463 7150 7497 7190
rect 7463 7076 7497 7116
rect 7463 7002 7497 7042
rect 7463 6927 7497 6968
rect 7463 6852 7497 6893
rect 7463 6777 7497 6818
rect 7463 6702 7497 6743
rect 7775 7224 7809 7264
rect 7775 7150 7809 7190
rect 7775 7076 7809 7116
rect 7775 7001 7809 7042
rect 7775 6926 7809 6967
rect 7775 6851 7809 6892
rect 7775 6776 7809 6817
rect 7775 6701 7809 6742
rect 8087 7224 8121 7264
rect 8087 7150 8121 7190
rect 8087 7076 8121 7116
rect 8087 7001 8121 7042
rect 8087 6926 8121 6967
rect 8087 6851 8121 6892
rect 8087 6776 8121 6817
rect 8087 6701 8121 6742
rect 8399 7224 8433 7264
rect 8399 7150 8433 7190
rect 8399 7076 8433 7116
rect 8399 7002 8433 7042
rect 8399 6927 8433 6968
rect 8399 6852 8433 6893
rect 8399 6777 8433 6818
rect 8399 6702 8433 6743
rect 8711 7224 8745 7264
rect 8711 7150 8745 7190
rect 8711 7076 8745 7116
rect 8711 7001 8745 7042
rect 8711 6926 8745 6967
rect 8711 6851 8745 6892
rect 8711 6776 8745 6817
rect 8711 6701 8745 6742
rect 9023 7224 9057 7264
rect 9023 7150 9057 7190
rect 9023 7076 9057 7116
rect 9023 7002 9057 7042
rect 9023 6927 9057 6968
rect 9023 6852 9057 6893
rect 9023 6777 9057 6818
rect 9023 6702 9057 6743
rect 9185 7297 9191 7314
rect 9151 7263 9157 7280
rect 9151 7246 9191 7263
rect 9185 7223 9191 7246
rect 9151 7189 9157 7212
rect 9151 7178 9191 7189
rect 9185 7149 9191 7178
rect 9151 7115 9157 7144
rect 9151 7110 9191 7115
rect 9185 7076 9191 7110
rect 9151 7075 9191 7076
rect 9151 7042 9157 7075
rect 9185 7008 9191 7041
rect 9151 7001 9191 7008
rect 9151 6974 9157 7001
rect 9185 6940 9191 6967
rect 9151 6926 9191 6940
rect 9151 6906 9157 6926
rect 9185 6872 9191 6892
rect 9151 6851 9191 6872
rect 9151 6838 9157 6851
rect 9185 6804 9191 6817
rect 9151 6776 9191 6804
rect 9151 6770 9157 6776
rect 9185 6736 9191 6742
rect 9151 6702 9191 6736
rect 9185 6701 9191 6702
rect 9151 6667 9157 6668
rect 947 6635 981 6663
rect 947 6567 981 6588
rect 9151 6634 9191 6667
rect 9185 6626 9191 6634
rect 9151 6592 9157 6600
rect 947 6499 981 6513
rect 947 6431 981 6438
rect 947 6363 981 6364
rect 947 6324 981 6329
rect 947 6250 981 6261
rect 947 6176 981 6193
rect 947 6102 981 6125
rect 947 6028 981 6057
rect 947 5954 981 5989
rect 1379 6500 1413 6538
rect 1379 6427 1413 6466
rect 1379 6354 1413 6393
rect 1379 6281 1413 6320
rect 1379 6208 1413 6247
rect 1379 6135 1413 6174
rect 1379 6062 1413 6101
rect 1379 5989 1413 6028
rect 1691 6499 1725 6538
rect 1691 6426 1725 6465
rect 1691 6353 1725 6392
rect 1691 6280 1725 6319
rect 1691 6207 1725 6246
rect 1691 6134 1725 6173
rect 1691 6061 1725 6100
rect 1691 5988 1725 6027
rect 2003 6500 2037 6538
rect 2003 6427 2037 6466
rect 2003 6354 2037 6393
rect 2003 6281 2037 6320
rect 2003 6208 2037 6247
rect 2003 6135 2037 6174
rect 2003 6062 2037 6101
rect 2003 5989 2037 6028
rect 2315 6499 2349 6538
rect 2315 6426 2349 6465
rect 2315 6353 2349 6392
rect 2315 6280 2349 6319
rect 2315 6207 2349 6246
rect 2315 6134 2349 6173
rect 2315 6061 2349 6100
rect 2315 5988 2349 6027
rect 2627 6500 2661 6538
rect 2627 6427 2661 6466
rect 2627 6354 2661 6393
rect 2627 6281 2661 6320
rect 2627 6208 2661 6247
rect 2627 6135 2661 6174
rect 2627 6062 2661 6101
rect 2627 5989 2661 6028
rect 2939 6499 2973 6538
rect 2939 6426 2973 6465
rect 2939 6353 2973 6392
rect 2939 6280 2973 6319
rect 2939 6207 2973 6246
rect 2939 6134 2973 6173
rect 2939 6061 2973 6100
rect 2939 5988 2973 6027
rect 3251 6499 3285 6538
rect 3251 6426 3285 6465
rect 3251 6353 3285 6392
rect 3251 6280 3285 6319
rect 3251 6207 3285 6246
rect 3251 6134 3285 6173
rect 3251 6061 3285 6100
rect 3251 5988 3285 6027
rect 3563 6499 3597 6538
rect 3563 6426 3597 6465
rect 3563 6353 3597 6392
rect 3563 6280 3597 6319
rect 3563 6207 3597 6246
rect 3563 6134 3597 6173
rect 3563 6061 3597 6100
rect 3563 5988 3597 6027
rect 3875 6500 3909 6538
rect 3875 6427 3909 6466
rect 3875 6354 3909 6393
rect 3875 6281 3909 6320
rect 3875 6208 3909 6247
rect 3875 6135 3909 6174
rect 3875 6062 3909 6101
rect 3875 5989 3909 6028
rect 4187 6499 4221 6538
rect 4187 6426 4221 6465
rect 4187 6353 4221 6392
rect 4187 6280 4221 6319
rect 4187 6207 4221 6246
rect 4187 6134 4221 6173
rect 4187 6061 4221 6100
rect 4187 5988 4221 6027
rect 4499 6500 4533 6538
rect 4499 6427 4533 6466
rect 4499 6354 4533 6393
rect 4499 6281 4533 6320
rect 4499 6208 4533 6247
rect 4499 6135 4533 6174
rect 4499 6062 4533 6101
rect 4499 5989 4533 6028
rect 4811 6499 4845 6538
rect 4811 6426 4845 6465
rect 4811 6353 4845 6392
rect 4811 6280 4845 6319
rect 4811 6207 4845 6246
rect 4811 6134 4845 6173
rect 4811 6061 4845 6100
rect 4811 5988 4845 6027
rect 5123 6500 5157 6538
rect 5123 6427 5157 6466
rect 5123 6354 5157 6393
rect 5123 6281 5157 6320
rect 5123 6208 5157 6247
rect 5123 6135 5157 6174
rect 5123 6062 5157 6101
rect 5123 5989 5157 6028
rect 5435 6499 5469 6538
rect 5435 6426 5469 6465
rect 5435 6353 5469 6392
rect 5435 6280 5469 6319
rect 5435 6207 5469 6246
rect 5435 6134 5469 6173
rect 5435 6061 5469 6100
rect 5435 5988 5469 6027
rect 5747 6500 5781 6538
rect 5747 6427 5781 6466
rect 5747 6354 5781 6393
rect 5747 6281 5781 6320
rect 5747 6208 5781 6247
rect 5747 6135 5781 6174
rect 5747 6062 5781 6101
rect 5747 5989 5781 6028
rect 6059 6499 6093 6538
rect 6059 6426 6093 6465
rect 6059 6353 6093 6392
rect 6059 6280 6093 6319
rect 6059 6207 6093 6246
rect 6059 6134 6093 6173
rect 6059 6061 6093 6100
rect 6059 5988 6093 6027
rect 6371 6500 6405 6538
rect 6371 6427 6405 6466
rect 6371 6354 6405 6393
rect 6371 6281 6405 6320
rect 6371 6208 6405 6247
rect 6371 6135 6405 6174
rect 6371 6062 6405 6101
rect 6371 5989 6405 6028
rect 6683 6499 6717 6538
rect 6683 6426 6717 6465
rect 6683 6353 6717 6392
rect 6683 6280 6717 6319
rect 6683 6207 6717 6246
rect 6683 6134 6717 6173
rect 6683 6061 6717 6100
rect 6683 5988 6717 6027
rect 6995 6500 7029 6538
rect 6995 6427 7029 6466
rect 6995 6354 7029 6393
rect 6995 6281 7029 6320
rect 6995 6208 7029 6247
rect 6995 6135 7029 6174
rect 6995 6062 7029 6101
rect 6995 5989 7029 6028
rect 7307 6499 7341 6538
rect 7307 6426 7341 6465
rect 7307 6353 7341 6392
rect 7307 6280 7341 6319
rect 7307 6207 7341 6246
rect 7307 6134 7341 6173
rect 7307 6061 7341 6100
rect 7307 5988 7341 6027
rect 7619 6500 7653 6538
rect 7619 6427 7653 6466
rect 7619 6354 7653 6393
rect 7619 6281 7653 6320
rect 7619 6208 7653 6247
rect 7619 6135 7653 6174
rect 7619 6062 7653 6101
rect 7619 5989 7653 6028
rect 7931 6499 7965 6538
rect 7931 6426 7965 6465
rect 7931 6353 7965 6392
rect 7931 6280 7965 6319
rect 7931 6207 7965 6246
rect 7931 6134 7965 6173
rect 7931 6061 7965 6100
rect 7931 5988 7965 6027
rect 8243 6499 8277 6538
rect 8243 6426 8277 6465
rect 8243 6353 8277 6392
rect 8243 6280 8277 6319
rect 8243 6207 8277 6246
rect 8243 6134 8277 6173
rect 8243 6061 8277 6100
rect 8243 5988 8277 6027
rect 8555 6500 8589 6538
rect 8555 6427 8589 6466
rect 8555 6354 8589 6393
rect 8555 6281 8589 6320
rect 8555 6208 8589 6247
rect 8555 6135 8589 6174
rect 8555 6062 8589 6101
rect 8555 5989 8589 6028
rect 8867 6499 8901 6538
rect 8867 6426 8901 6465
rect 8867 6353 8901 6392
rect 8867 6280 8901 6319
rect 8867 6207 8901 6246
rect 8867 6134 8901 6173
rect 8867 6061 8901 6100
rect 8867 5988 8901 6027
rect 9151 6566 9191 6592
rect 9185 6551 9191 6566
rect 9151 6517 9157 6532
rect 9151 6498 9191 6517
rect 9185 6476 9191 6498
rect 9151 6442 9157 6464
rect 9151 6430 9191 6442
rect 9185 6401 9191 6430
rect 9151 6367 9157 6396
rect 9151 6362 9191 6367
rect 9185 6328 9191 6362
rect 9151 6326 9191 6328
rect 9151 6294 9157 6326
rect 9185 6260 9191 6292
rect 9151 6251 9191 6260
rect 9151 6226 9157 6251
rect 9185 6192 9191 6217
rect 9151 6176 9191 6192
rect 9151 6158 9157 6176
rect 9185 6124 9191 6142
rect 9151 6101 9191 6124
rect 9151 6090 9157 6101
rect 9185 6056 9191 6067
rect 9151 6026 9191 6056
rect 9151 6022 9157 6026
rect 9185 5988 9191 5992
rect 9151 5954 9191 5988
rect 947 5886 981 5920
rect 9185 5951 9191 5954
rect 9151 5917 9157 5920
rect 9151 5886 9191 5917
rect 9636 7549 9640 7589
rect 9462 7477 9466 7517
rect 9636 7475 9640 7515
rect 9462 7403 9466 7443
rect 9636 7401 9640 7441
rect 9462 7329 9466 7369
rect 9636 7327 9640 7367
rect 9462 7255 9466 7295
rect 9636 7253 9640 7293
rect 9462 7181 9466 7221
rect 9636 7180 9640 7219
rect 9462 7107 9466 7147
rect 9636 7107 9640 7146
rect 9462 7034 9466 7073
rect 9636 7034 9640 7073
rect 9462 6961 9466 7000
rect 9636 6961 9640 7000
rect 9462 6888 9466 6927
rect 9636 6888 9640 6927
rect 9462 6815 9466 6854
rect 9636 6815 9640 6854
rect 9462 6742 9466 6781
rect 9636 6742 9640 6781
rect 9462 6669 9466 6708
rect 9636 6669 9640 6708
rect 9462 6596 9466 6635
rect 9636 6596 9640 6635
rect 9462 6523 9466 6562
rect 9636 6523 9640 6562
rect 9462 6450 9466 6489
rect 9636 6450 9640 6489
rect 9462 6377 9466 6416
rect 9636 6377 9640 6416
rect 9462 6304 9466 6343
rect 9636 6304 9640 6343
rect 9462 6231 9466 6270
rect 9636 6231 9640 6270
rect 9462 6158 9466 6197
rect 9636 6158 9640 6197
rect 9462 6085 9466 6124
rect 9636 6085 9640 6124
rect 9462 6012 9466 6051
rect 9636 6012 9640 6051
rect 9462 5939 9466 5978
rect 9636 5939 9640 5978
rect 10464 7915 10605 7917
rect 10498 7913 10536 7915
rect 10507 7881 10536 7913
rect 10570 7883 10605 7915
rect 10570 7881 10642 7883
rect 10464 7879 10473 7881
rect 10507 7879 10642 7881
rect 10464 7849 10642 7879
rect 10464 7845 10605 7849
rect 10464 7842 10473 7845
rect 10507 7842 10605 7845
rect 10639 7844 10642 7849
rect 10507 7811 10536 7842
rect 10498 7808 10536 7811
rect 10570 7815 10605 7842
rect 10570 7810 10608 7815
rect 10570 7808 10642 7810
rect 10464 7781 10642 7808
rect 10464 7777 10605 7781
rect 10464 7769 10473 7777
rect 10507 7769 10605 7777
rect 10639 7771 10642 7781
rect 10507 7743 10536 7769
rect 10498 7735 10536 7743
rect 10570 7747 10605 7769
rect 10570 7737 10608 7747
rect 10570 7735 10642 7737
rect 10464 7713 10642 7735
rect 10464 7709 10605 7713
rect 10464 7696 10473 7709
rect 10507 7696 10605 7709
rect 10639 7698 10642 7713
rect 10507 7675 10536 7696
rect 10498 7662 10536 7675
rect 10570 7679 10605 7696
rect 10570 7664 10608 7679
rect 10570 7662 10642 7664
rect 10464 7645 10642 7662
rect 10464 7641 10605 7645
rect 10464 7623 10473 7641
rect 10507 7623 10605 7641
rect 10639 7625 10642 7645
rect 10507 7607 10536 7623
rect 10498 7589 10536 7607
rect 10570 7611 10605 7623
rect 10570 7591 10608 7611
rect 10570 7589 10642 7591
rect 10464 7577 10642 7589
rect 10464 7573 10605 7577
rect 10464 7550 10473 7573
rect 10507 7550 10605 7573
rect 10639 7552 10642 7577
rect 10507 7539 10536 7550
rect 10498 7516 10536 7539
rect 10570 7543 10605 7550
rect 10570 7518 10608 7543
rect 10570 7516 10642 7518
rect 10464 7509 10642 7516
rect 10464 7505 10605 7509
rect 10464 7477 10473 7505
rect 10507 7477 10605 7505
rect 10639 7479 10642 7509
rect 10507 7471 10536 7477
rect 10498 7443 10536 7471
rect 10570 7475 10605 7477
rect 10570 7445 10608 7475
rect 10570 7443 10642 7445
rect 10464 7441 10642 7443
rect 10464 7437 10605 7441
rect 10464 7404 10473 7437
rect 10507 7407 10605 7437
rect 10639 7407 10642 7441
rect 10507 7406 10642 7407
rect 10507 7404 10608 7406
rect 10507 7403 10536 7404
rect 10498 7370 10536 7403
rect 10570 7373 10608 7404
rect 10570 7370 10605 7373
rect 10464 7369 10605 7370
rect 10464 7335 10473 7369
rect 10507 7339 10605 7369
rect 10639 7339 10642 7372
rect 10507 7335 10642 7339
rect 10464 7333 10642 7335
rect 10464 7331 10608 7333
rect 10498 7301 10536 7331
rect 10507 7297 10536 7301
rect 10570 7305 10608 7331
rect 10570 7297 10605 7305
rect 10464 7267 10473 7297
rect 10507 7271 10605 7297
rect 10639 7271 10642 7299
rect 10507 7267 10642 7271
rect 10464 7260 10642 7267
rect 10464 7258 10608 7260
rect 10498 7233 10536 7258
rect 10507 7224 10536 7233
rect 10570 7237 10608 7258
rect 10570 7224 10605 7237
rect 10464 7199 10473 7224
rect 10507 7203 10605 7224
rect 10639 7203 10642 7226
rect 10507 7199 10642 7203
rect 10464 7187 10642 7199
rect 10464 7185 10608 7187
rect 10498 7165 10536 7185
rect 10507 7151 10536 7165
rect 10570 7169 10608 7185
rect 10570 7151 10605 7169
rect 10464 7131 10473 7151
rect 10507 7135 10605 7151
rect 10639 7135 10642 7153
rect 10507 7131 10642 7135
rect 10464 7113 10642 7131
rect 10464 7112 10608 7113
rect 10498 7097 10536 7112
rect 10507 7078 10536 7097
rect 10570 7101 10608 7112
rect 10570 7078 10605 7101
rect 10464 7063 10473 7078
rect 10507 7067 10605 7078
rect 10639 7067 10642 7079
rect 10507 7063 10642 7067
rect 10464 7039 10642 7063
rect 10498 7029 10536 7039
rect 10507 7005 10536 7029
rect 10570 7033 10608 7039
rect 10570 7005 10605 7033
rect 10464 6995 10473 7005
rect 10507 6999 10605 7005
rect 10639 6999 10642 7005
rect 10507 6995 10642 6999
rect 10464 6965 10642 6995
rect 10498 6961 10536 6965
rect 10507 6931 10536 6961
rect 10570 6931 10605 6965
rect 10464 6927 10473 6931
rect 10507 6927 10642 6931
rect 10464 6897 10642 6927
rect 10464 6893 10605 6897
rect 10464 6891 10473 6893
rect 10507 6891 10605 6893
rect 10639 6891 10642 6897
rect 10507 6859 10536 6891
rect 10498 6857 10536 6859
rect 10570 6863 10605 6891
rect 10570 6857 10608 6863
rect 10464 6829 10642 6857
rect 10464 6825 10605 6829
rect 10464 6817 10473 6825
rect 10507 6817 10605 6825
rect 10639 6817 10642 6829
rect 10507 6791 10536 6817
rect 10498 6783 10536 6791
rect 10570 6795 10605 6817
rect 10570 6783 10608 6795
rect 10464 6761 10642 6783
rect 10464 6757 10605 6761
rect 10464 6743 10473 6757
rect 10507 6743 10605 6757
rect 10639 6743 10642 6761
rect 10507 6723 10536 6743
rect 10498 6709 10536 6723
rect 10570 6727 10605 6743
rect 10570 6709 10608 6727
rect 10464 6693 10642 6709
rect 10464 6689 10605 6693
rect 10464 6669 10473 6689
rect 10507 6669 10605 6689
rect 10639 6669 10642 6693
rect 10507 6655 10536 6669
rect 10498 6635 10536 6655
rect 10570 6659 10605 6669
rect 10570 6635 10608 6659
rect 10464 6625 10642 6635
rect 10464 6621 10605 6625
rect 10464 6595 10473 6621
rect 10507 6595 10605 6621
rect 10639 6595 10642 6625
rect 10507 6587 10536 6595
rect 10498 6561 10536 6587
rect 10570 6591 10605 6595
rect 10570 6561 10608 6591
rect 10464 6557 10642 6561
rect 10464 6553 10605 6557
rect 10464 6521 10473 6553
rect 10507 6523 10605 6553
rect 10639 6523 10642 6557
rect 10507 6521 10642 6523
rect 10507 6519 10536 6521
rect 10498 6487 10536 6519
rect 10570 6489 10608 6521
rect 10570 6487 10605 6489
rect 10464 6485 10605 6487
rect 10464 6451 10473 6485
rect 10507 6455 10605 6485
rect 10639 6455 10642 6487
rect 10507 6451 10642 6455
rect 10464 6428 10642 6451
rect 10498 6394 10536 6428
rect 10570 6394 10608 6428
rect 10464 6350 10642 6394
rect 10792 8082 10864 8116
rect 10912 8082 10936 8116
rect 10980 8082 11008 8116
rect 11048 8082 11080 8116
rect 11116 8082 11150 8116
rect 11186 8082 11218 8116
rect 11258 8082 11286 8116
rect 11330 8082 11354 8116
rect 11402 8082 11422 8116
rect 11474 8082 11490 8116
rect 11546 8082 11558 8116
rect 11618 8082 11626 8116
rect 11690 8082 11694 8116
rect 11796 8082 11800 8116
rect 11864 8082 11872 8116
rect 11932 8082 11944 8116
rect 12000 8082 12016 8116
rect 12068 8082 12088 8116
rect 12136 8082 12160 8116
rect 12204 8082 12232 8116
rect 12272 8082 12304 8116
rect 12340 8082 12374 8116
rect 12410 8082 12442 8116
rect 12482 8082 12510 8116
rect 12554 8082 12578 8116
rect 12626 8082 12646 8116
rect 12698 8082 12714 8116
rect 12770 8082 12782 8116
rect 12842 8082 12850 8116
rect 12914 8082 12918 8116
rect 13020 8082 13024 8116
rect 13088 8082 13096 8116
rect 13156 8082 13169 8116
rect 13224 8082 13242 8116
rect 13292 8082 13315 8116
rect 13360 8082 13428 8116
rect 13634 8096 13732 8116
rect 10792 8048 10826 8082
rect 10792 7980 10826 8014
rect 13387 8041 13428 8082
rect 13421 8033 13428 8041
rect 13387 7999 13394 8007
rect 10988 7954 10995 7988
rect 11038 7954 11070 7988
rect 11108 7954 11144 7988
rect 11179 7954 11214 7988
rect 11254 7954 11284 7988
rect 11329 7954 11354 7988
rect 11404 7954 11423 7988
rect 11479 7954 11492 7988
rect 11553 7954 11561 7988
rect 11627 7954 11630 7988
rect 11664 7954 11667 7988
rect 11733 7954 11741 7988
rect 11802 7954 11815 7988
rect 11871 7954 11889 7988
rect 11940 7954 11963 7988
rect 12009 7954 12037 7988
rect 12078 7954 12111 7988
rect 12147 7954 12182 7988
rect 12219 7954 12251 7988
rect 12293 7954 12320 7988
rect 12367 7954 12389 7988
rect 12441 7954 12458 7988
rect 12515 7954 12527 7988
rect 12589 7954 12596 7988
rect 12663 7954 12665 7988
rect 12699 7954 12703 7988
rect 12768 7954 12777 7988
rect 12837 7954 12851 7988
rect 12906 7954 12925 7988
rect 12975 7954 12999 7988
rect 13044 7954 13073 7988
rect 13113 7954 13147 7988
rect 13182 7954 13217 7988
rect 13255 7954 13267 7988
rect 13387 7966 13428 7999
rect 13421 7965 13428 7966
rect 10792 7912 10826 7946
rect 10792 7858 10826 7878
rect 13387 7931 13394 7932
rect 13387 7897 13428 7931
rect 13387 7891 13394 7897
rect 10792 7784 10826 7810
rect 10792 7710 10826 7742
rect 10792 7640 10826 7674
rect 10792 7572 10826 7602
rect 10792 7504 10826 7529
rect 10792 7436 10826 7456
rect 10792 7368 10826 7383
rect 10792 7300 10826 7310
rect 10939 7785 10973 7824
rect 10939 7712 10973 7751
rect 10939 7639 10973 7678
rect 10939 7566 10973 7605
rect 10939 7493 10973 7532
rect 10939 7420 10973 7459
rect 10939 7346 10973 7386
rect 10939 7272 10973 7312
rect 11251 7785 11285 7824
rect 11251 7712 11285 7751
rect 11251 7639 11285 7678
rect 11251 7566 11285 7605
rect 11251 7493 11285 7532
rect 11251 7420 11285 7459
rect 11251 7346 11285 7386
rect 11251 7272 11285 7312
rect 11563 7785 11597 7824
rect 11563 7712 11597 7751
rect 11563 7639 11597 7678
rect 11563 7566 11597 7605
rect 11563 7493 11597 7532
rect 11563 7420 11597 7459
rect 11563 7346 11597 7386
rect 11563 7272 11597 7312
rect 11875 7785 11909 7824
rect 11875 7712 11909 7751
rect 11875 7639 11909 7678
rect 11875 7566 11909 7605
rect 11875 7493 11909 7532
rect 11875 7420 11909 7459
rect 11875 7346 11909 7386
rect 11875 7272 11909 7312
rect 12187 7785 12221 7824
rect 12187 7712 12221 7751
rect 12187 7639 12221 7678
rect 12187 7566 12221 7605
rect 12187 7493 12221 7532
rect 12187 7420 12221 7459
rect 12187 7346 12221 7386
rect 12187 7272 12221 7312
rect 12499 7785 12533 7824
rect 12499 7712 12533 7751
rect 12499 7639 12533 7678
rect 12499 7566 12533 7605
rect 12499 7493 12533 7532
rect 12499 7420 12533 7459
rect 12499 7346 12533 7386
rect 12499 7272 12533 7312
rect 12811 7785 12845 7824
rect 12811 7712 12845 7751
rect 12811 7639 12845 7678
rect 12811 7566 12845 7605
rect 12811 7493 12845 7532
rect 12811 7420 12845 7459
rect 12811 7346 12845 7386
rect 12811 7272 12845 7312
rect 13123 7785 13157 7824
rect 13123 7712 13157 7751
rect 13123 7639 13157 7678
rect 13123 7566 13157 7605
rect 13123 7493 13157 7532
rect 13123 7420 13157 7459
rect 13123 7346 13157 7386
rect 13123 7272 13157 7312
rect 13421 7857 13428 7863
rect 13387 7829 13428 7857
rect 13387 7816 13394 7829
rect 13421 7782 13428 7795
rect 13387 7761 13428 7782
rect 13387 7741 13394 7761
rect 13421 7707 13428 7727
rect 13387 7693 13428 7707
rect 13387 7666 13394 7693
rect 13421 7632 13428 7659
rect 13387 7625 13428 7632
rect 13387 7591 13394 7625
rect 13421 7557 13428 7591
rect 13387 7523 13394 7557
rect 13387 7516 13428 7523
rect 13421 7489 13428 7516
rect 13387 7455 13394 7482
rect 13387 7441 13428 7455
rect 13421 7421 13428 7441
rect 13387 7387 13394 7407
rect 13387 7365 13428 7387
rect 13421 7353 13428 7365
rect 13387 7319 13394 7331
rect 13387 7289 13428 7319
rect 13421 7285 13428 7289
rect 10792 7232 10826 7237
rect 13394 7217 13428 7251
rect 10792 7164 10826 7198
rect 13421 7179 13428 7183
rect 10792 7096 10826 7130
rect 10792 7028 10826 7062
rect 10792 6960 10826 6994
rect 10792 6892 10826 6926
rect 10792 6824 10826 6858
rect 10792 6756 10826 6790
rect 10792 6688 10826 6722
rect 10792 6620 10826 6654
rect 10792 6552 10826 6586
rect 11093 7080 11127 7120
rect 11093 7006 11127 7046
rect 11093 6932 11127 6972
rect 11093 6858 11127 6898
rect 11093 6783 11127 6824
rect 11093 6708 11127 6749
rect 11093 6633 11127 6674
rect 11093 6558 11127 6599
rect 11405 7080 11439 7120
rect 11405 7006 11439 7046
rect 11405 6932 11439 6972
rect 11405 6858 11439 6898
rect 11405 6783 11439 6824
rect 11405 6708 11439 6749
rect 11405 6633 11439 6674
rect 11405 6558 11439 6599
rect 11717 7080 11751 7120
rect 11717 7006 11751 7046
rect 11717 6932 11751 6972
rect 11717 6858 11751 6898
rect 11717 6783 11751 6824
rect 11717 6708 11751 6749
rect 11717 6633 11751 6674
rect 11717 6558 11751 6599
rect 12029 7080 12063 7120
rect 12029 7006 12063 7046
rect 12029 6932 12063 6972
rect 12029 6858 12063 6898
rect 12029 6783 12063 6824
rect 12029 6708 12063 6749
rect 12029 6633 12063 6674
rect 12029 6558 12063 6599
rect 12341 7080 12375 7120
rect 12341 7006 12375 7046
rect 12341 6932 12375 6972
rect 12341 6858 12375 6898
rect 12341 6783 12375 6824
rect 12341 6708 12375 6749
rect 12341 6633 12375 6674
rect 12341 6558 12375 6599
rect 12653 7080 12687 7120
rect 12653 7006 12687 7046
rect 12653 6932 12687 6972
rect 12653 6858 12687 6898
rect 12653 6783 12687 6824
rect 12653 6708 12687 6749
rect 12653 6633 12687 6674
rect 12653 6558 12687 6599
rect 12965 7080 12999 7120
rect 12965 7006 12999 7046
rect 12965 6932 12999 6972
rect 12965 6858 12999 6898
rect 12965 6783 12999 6824
rect 12965 6708 12999 6749
rect 12965 6633 12999 6674
rect 12965 6558 12999 6599
rect 13277 7080 13311 7120
rect 13277 7006 13311 7046
rect 13277 6932 13311 6972
rect 13277 6858 13311 6898
rect 13277 6783 13311 6824
rect 13277 6708 13311 6749
rect 13277 6633 13311 6674
rect 13277 6558 13311 6599
rect 13387 7149 13428 7179
rect 13387 7139 13394 7149
rect 13421 7105 13428 7115
rect 13387 7081 13428 7105
rect 13387 7065 13394 7081
rect 13421 7031 13428 7047
rect 13387 7013 13428 7031
rect 13387 6991 13394 7013
rect 13421 6957 13428 6979
rect 13387 6945 13428 6957
rect 13387 6917 13394 6945
rect 13421 6883 13428 6911
rect 13387 6877 13428 6883
rect 13387 6843 13394 6877
rect 13421 6809 13428 6843
rect 13387 6775 13394 6809
rect 13387 6769 13428 6775
rect 13421 6741 13428 6769
rect 13387 6707 13394 6735
rect 13387 6695 13428 6707
rect 13421 6673 13428 6695
rect 13387 6639 13394 6661
rect 13387 6621 13428 6639
rect 13421 6605 13428 6621
rect 13387 6571 13394 6587
rect 13387 6547 13428 6571
rect 13421 6537 13428 6547
rect 10792 6401 10826 6518
rect 13387 6503 13394 6513
rect 13387 6473 13428 6503
rect 13421 6469 13428 6473
rect 13387 6435 13394 6439
rect 13387 6401 13428 6435
rect 10792 6367 10860 6401
rect 10898 6367 10928 6401
rect 10971 6367 10996 6401
rect 11044 6367 11064 6401
rect 11117 6367 11132 6401
rect 11189 6367 11200 6401
rect 11261 6367 11268 6401
rect 11333 6367 11336 6401
rect 11370 6367 11371 6401
rect 11438 6367 11443 6401
rect 11506 6367 11515 6401
rect 11574 6367 11587 6401
rect 11642 6367 11659 6401
rect 11710 6367 11731 6401
rect 11778 6367 11803 6401
rect 11846 6367 11875 6401
rect 11914 6367 11947 6401
rect 11982 6367 12016 6401
rect 12053 6367 12084 6401
rect 12125 6367 12152 6401
rect 12197 6367 12220 6401
rect 12269 6367 12288 6401
rect 12341 6367 12356 6401
rect 12413 6367 12424 6401
rect 12485 6367 12492 6401
rect 12557 6367 12560 6401
rect 12594 6367 12595 6401
rect 12662 6367 12667 6401
rect 12730 6367 12739 6401
rect 12798 6367 12811 6401
rect 12866 6367 12883 6401
rect 12934 6367 12955 6401
rect 13002 6367 13027 6401
rect 13070 6367 13099 6401
rect 13138 6367 13171 6401
rect 13206 6367 13240 6401
rect 13277 6367 13308 6401
rect 13349 6367 13428 6401
rect 13634 8082 13667 8096
rect 13629 8062 13667 8082
rect 13701 8086 13732 8096
rect 13701 8062 13739 8086
rect 13595 8052 13773 8062
rect 13595 8048 13732 8052
rect 13595 8022 13600 8048
rect 13634 8022 13732 8048
rect 13766 8022 13773 8052
rect 13634 8014 13667 8022
rect 13629 7988 13667 8014
rect 13701 8018 13732 8022
rect 13701 7988 13739 8018
rect 13595 7984 13773 7988
rect 13595 7980 13732 7984
rect 13595 7948 13600 7980
rect 13634 7950 13732 7980
rect 13766 7950 13773 7984
rect 13634 7948 13773 7950
rect 13634 7946 13667 7948
rect 13629 7914 13667 7946
rect 13701 7916 13739 7948
rect 13701 7914 13732 7916
rect 13595 7912 13732 7914
rect 13595 7878 13600 7912
rect 13634 7882 13732 7912
rect 13766 7882 13773 7914
rect 13634 7878 13773 7882
rect 13595 7874 13773 7878
rect 13629 7844 13667 7874
rect 13634 7840 13667 7844
rect 13701 7848 13739 7874
rect 13701 7840 13732 7848
rect 13595 7810 13600 7840
rect 13634 7814 13732 7840
rect 13766 7814 13773 7840
rect 13634 7810 13773 7814
rect 13595 7800 13773 7810
rect 13629 7776 13667 7800
rect 13634 7766 13667 7776
rect 13701 7780 13739 7800
rect 13701 7766 13732 7780
rect 13595 7742 13600 7766
rect 13634 7746 13732 7766
rect 13766 7746 13773 7766
rect 13634 7742 13773 7746
rect 13595 7726 13773 7742
rect 13629 7708 13667 7726
rect 13634 7692 13667 7708
rect 13701 7712 13739 7726
rect 13701 7692 13732 7712
rect 13595 7674 13600 7692
rect 13634 7678 13732 7692
rect 13766 7678 13773 7692
rect 13634 7674 13773 7678
rect 13595 7652 13773 7674
rect 13629 7640 13667 7652
rect 13634 7618 13667 7640
rect 13701 7644 13739 7652
rect 13701 7618 13732 7644
rect 13595 7606 13600 7618
rect 13634 7610 13732 7618
rect 13766 7610 13773 7618
rect 13634 7606 13773 7610
rect 13595 7578 13773 7606
rect 13629 7572 13667 7578
rect 13634 7544 13667 7572
rect 13701 7576 13739 7578
rect 13701 7544 13732 7576
rect 13595 7538 13600 7544
rect 13634 7542 13732 7544
rect 13766 7542 13773 7544
rect 13634 7538 13773 7542
rect 13595 7508 13773 7538
rect 13595 7504 13732 7508
rect 13766 7504 13773 7508
rect 13634 7470 13667 7504
rect 13701 7474 13732 7504
rect 13701 7470 13739 7474
rect 13595 7440 13773 7470
rect 13595 7436 13732 7440
rect 13595 7430 13600 7436
rect 13634 7431 13732 7436
rect 13766 7431 13773 7440
rect 13634 7402 13667 7431
rect 13629 7397 13667 7402
rect 13701 7406 13732 7431
rect 13701 7397 13739 7406
rect 13629 7396 13773 7397
rect 13595 7372 13773 7396
rect 13595 7368 13732 7372
rect 13595 7356 13600 7368
rect 13634 7358 13732 7368
rect 13766 7358 13773 7372
rect 13634 7334 13667 7358
rect 13629 7324 13667 7334
rect 13701 7338 13732 7358
rect 13701 7324 13739 7338
rect 13629 7322 13773 7324
rect 13595 7304 13773 7322
rect 13595 7300 13732 7304
rect 13595 7283 13600 7300
rect 13634 7285 13732 7300
rect 13766 7285 13773 7304
rect 13634 7266 13667 7285
rect 13629 7251 13667 7266
rect 13701 7270 13732 7285
rect 13701 7251 13739 7270
rect 13629 7249 13773 7251
rect 13595 7236 13773 7249
rect 13595 7232 13732 7236
rect 13595 7210 13600 7232
rect 13634 7212 13732 7232
rect 13766 7212 13773 7236
rect 13634 7198 13667 7212
rect 13629 7178 13667 7198
rect 13701 7202 13732 7212
rect 13701 7178 13739 7202
rect 13629 7176 13773 7178
rect 13595 7168 13773 7176
rect 13595 7164 13732 7168
rect 13595 7137 13600 7164
rect 13634 7139 13732 7164
rect 13766 7139 13773 7168
rect 13634 7130 13667 7139
rect 13629 7105 13667 7130
rect 13701 7134 13732 7139
rect 13701 7105 13739 7134
rect 13629 7103 13773 7105
rect 13595 7100 13773 7103
rect 13595 7096 13732 7100
rect 13595 7064 13600 7096
rect 13634 7066 13732 7096
rect 13766 7066 13773 7100
rect 13634 7062 13667 7066
rect 13629 7032 13667 7062
rect 13701 7032 13739 7066
rect 13629 7030 13732 7032
rect 13595 7028 13732 7030
rect 13595 6994 13600 7028
rect 13634 6998 13732 7028
rect 13766 6998 13773 7032
rect 13634 6994 13773 6998
rect 13595 6993 13773 6994
rect 13595 6991 13667 6993
rect 13629 6960 13667 6991
rect 13634 6959 13667 6960
rect 13701 6964 13739 6993
rect 13701 6959 13732 6964
rect 13595 6926 13600 6957
rect 13634 6930 13732 6959
rect 13766 6930 13773 6959
rect 13634 6926 13773 6930
rect 13595 6920 13773 6926
rect 13595 6918 13667 6920
rect 13629 6892 13667 6918
rect 13634 6886 13667 6892
rect 13701 6896 13739 6920
rect 13701 6886 13732 6896
rect 13595 6858 13600 6884
rect 13634 6862 13732 6886
rect 13766 6862 13773 6886
rect 13634 6858 13773 6862
rect 13595 6847 13773 6858
rect 13595 6845 13667 6847
rect 13629 6824 13667 6845
rect 13634 6813 13667 6824
rect 13701 6828 13739 6847
rect 13701 6813 13732 6828
rect 13595 6790 13600 6811
rect 13634 6794 13732 6813
rect 13766 6794 13773 6813
rect 13634 6790 13773 6794
rect 13595 6774 13773 6790
rect 13595 6772 13667 6774
rect 13629 6756 13667 6772
rect 13634 6740 13667 6756
rect 13701 6760 13739 6774
rect 13701 6740 13732 6760
rect 13595 6722 13600 6738
rect 13634 6726 13732 6740
rect 13766 6726 13773 6740
rect 13634 6722 13773 6726
rect 13595 6701 13773 6722
rect 13595 6699 13667 6701
rect 13629 6688 13667 6699
rect 13634 6667 13667 6688
rect 13701 6692 13739 6701
rect 13701 6667 13732 6692
rect 13595 6654 13600 6665
rect 13634 6658 13732 6667
rect 13766 6658 13773 6667
rect 13634 6654 13773 6658
rect 13595 6628 13773 6654
rect 13595 6626 13667 6628
rect 13629 6620 13667 6626
rect 13634 6594 13667 6620
rect 13701 6624 13739 6628
rect 13701 6594 13732 6624
rect 13595 6586 13600 6592
rect 13634 6590 13732 6594
rect 13766 6590 13773 6594
rect 13634 6586 13773 6590
rect 13595 6556 13773 6586
rect 13595 6555 13732 6556
rect 13766 6555 13773 6556
rect 13595 6553 13667 6555
rect 13629 6552 13667 6553
rect 13634 6521 13667 6552
rect 13701 6522 13732 6555
rect 13701 6521 13739 6522
rect 13595 6518 13600 6519
rect 13634 6518 13773 6521
rect 13595 6488 13773 6518
rect 13595 6484 13732 6488
rect 13595 6480 13600 6484
rect 13634 6482 13732 6484
rect 13766 6482 13773 6488
rect 13634 6450 13667 6482
rect 13629 6448 13667 6450
rect 13701 6454 13732 6482
rect 13701 6448 13739 6454
rect 13629 6446 13773 6448
rect 13595 6420 13773 6446
rect 13595 6416 13732 6420
rect 13595 6407 13600 6416
rect 13634 6409 13732 6416
rect 13766 6409 13773 6420
rect 13634 6382 13667 6409
rect 13629 6375 13667 6382
rect 13701 6386 13732 6409
rect 13701 6375 13739 6386
rect 13629 6373 13773 6375
rect 10498 6329 10536 6350
rect 10507 6316 10536 6329
rect 10570 6348 10642 6350
rect 10570 6329 10608 6348
rect 10570 6316 10605 6329
rect 10464 6295 10473 6316
rect 10507 6295 10605 6316
rect 10639 6295 10642 6314
rect 10464 6272 10642 6295
rect 10498 6261 10536 6272
rect 10507 6238 10536 6261
rect 10570 6268 10642 6272
rect 10570 6238 10608 6268
rect 10464 6227 10473 6238
rect 10507 6234 10608 6238
rect 10507 6227 10642 6234
rect 10464 6212 10642 6227
rect 13595 6352 13773 6373
rect 13595 6348 13732 6352
rect 13595 6334 13600 6348
rect 13634 6336 13732 6348
rect 13766 6336 13773 6352
rect 13634 6314 13667 6336
rect 13629 6302 13667 6314
rect 13701 6318 13732 6336
rect 13701 6302 13739 6318
rect 13629 6300 13773 6302
rect 13595 6284 13773 6300
rect 13595 6280 13732 6284
rect 13595 6261 13600 6280
rect 13634 6263 13732 6280
rect 13766 6263 13773 6284
rect 13634 6246 13667 6263
rect 13629 6229 13667 6246
rect 13701 6250 13732 6263
rect 13701 6229 13739 6250
rect 13629 6227 13773 6229
rect 13595 6216 13773 6227
rect 13595 6212 13732 6216
rect 10464 6194 10605 6212
rect 10498 6193 10536 6194
rect 10507 6160 10536 6193
rect 10570 6178 10605 6194
rect 10639 6188 10673 6212
rect 10707 6188 10741 6212
rect 10775 6188 10809 6212
rect 10843 6188 10877 6212
rect 10911 6188 10945 6212
rect 10979 6188 11013 6212
rect 11047 6188 11081 6212
rect 11115 6188 11149 6212
rect 11074 6178 11081 6188
rect 11147 6178 11149 6188
rect 11183 6188 11217 6212
rect 11251 6188 11285 6212
rect 11319 6188 11353 6212
rect 11387 6188 11421 6212
rect 11455 6188 11489 6212
rect 11523 6188 11557 6212
rect 11591 6188 11625 6212
rect 11183 6178 11186 6188
rect 11251 6178 11259 6188
rect 11319 6178 11332 6188
rect 11387 6178 11405 6188
rect 11455 6178 11478 6188
rect 11523 6178 11551 6188
rect 11591 6178 11624 6188
rect 11659 6178 11693 6212
rect 11727 6188 11761 6212
rect 11795 6188 11829 6212
rect 11863 6188 11897 6212
rect 11931 6188 11965 6212
rect 11999 6188 12033 6212
rect 12067 6188 12101 6212
rect 11731 6178 11761 6188
rect 11804 6178 11829 6188
rect 11877 6178 11897 6188
rect 11950 6178 11965 6188
rect 12023 6178 12033 6188
rect 12096 6178 12101 6188
rect 12135 6188 12169 6212
rect 10570 6160 10608 6178
rect 10464 6159 10473 6160
rect 10507 6159 10608 6160
rect 10464 6116 10608 6159
rect 11074 6154 11113 6178
rect 11147 6154 11186 6178
rect 11220 6154 11259 6178
rect 11293 6154 11332 6178
rect 11366 6154 11405 6178
rect 11439 6154 11478 6178
rect 11512 6154 11551 6178
rect 11585 6154 11624 6178
rect 11658 6154 11697 6178
rect 11731 6154 11770 6178
rect 11804 6154 11843 6178
rect 11877 6154 11916 6178
rect 11950 6154 11989 6178
rect 12023 6154 12062 6178
rect 12096 6154 12135 6178
rect 12203 6188 12237 6212
rect 12271 6188 12305 6212
rect 12339 6188 12373 6212
rect 12407 6188 12441 6212
rect 12475 6188 12509 6212
rect 12543 6188 12577 6212
rect 12203 6178 12208 6188
rect 12271 6178 12281 6188
rect 12339 6178 12354 6188
rect 12407 6178 12427 6188
rect 12475 6178 12500 6188
rect 12543 6178 12573 6188
rect 12611 6178 12645 6212
rect 12679 6188 12713 6212
rect 12747 6188 12781 6212
rect 12815 6188 12849 6212
rect 12883 6188 12917 6212
rect 12951 6188 12985 6212
rect 13019 6188 13053 6212
rect 13087 6188 13121 6212
rect 12680 6178 12713 6188
rect 12753 6178 12781 6188
rect 12826 6178 12849 6188
rect 12899 6178 12917 6188
rect 12972 6178 12985 6188
rect 13045 6178 13053 6188
rect 13118 6178 13121 6188
rect 13155 6188 13189 6212
rect 13223 6188 13257 6212
rect 13291 6188 13325 6212
rect 13359 6188 13393 6212
rect 13427 6188 13461 6212
rect 13495 6188 13529 6212
rect 13563 6188 13600 6212
rect 13634 6190 13732 6212
rect 13766 6190 13773 6216
rect 13155 6178 13157 6188
rect 13223 6178 13230 6188
rect 13291 6178 13303 6188
rect 13359 6178 13376 6188
rect 13427 6178 13449 6188
rect 13495 6178 13522 6188
rect 13563 6178 13595 6188
rect 13634 6178 13667 6190
rect 12169 6154 12208 6178
rect 12242 6154 12281 6178
rect 12315 6154 12354 6178
rect 12388 6154 12427 6178
rect 12461 6154 12500 6178
rect 12534 6154 12573 6178
rect 12607 6154 12646 6178
rect 12680 6154 12719 6178
rect 12753 6154 12792 6178
rect 12826 6154 12865 6178
rect 12899 6154 12938 6178
rect 12972 6154 13011 6178
rect 13045 6154 13084 6178
rect 13118 6154 13157 6178
rect 13191 6154 13230 6178
rect 13264 6154 13303 6178
rect 13337 6154 13376 6178
rect 13410 6154 13449 6178
rect 13483 6154 13522 6178
rect 13556 6154 13595 6178
rect 13629 6156 13667 6178
rect 13701 6182 13732 6190
rect 13701 6156 13739 6182
rect 13629 6154 13773 6156
rect 11074 6148 13773 6154
rect 11074 6116 13732 6148
rect 13766 6117 13773 6148
rect 10498 6082 10536 6116
rect 10464 6010 10536 6082
rect 11146 6082 11185 6116
rect 11219 6082 11258 6116
rect 11292 6082 11331 6116
rect 11365 6082 11404 6116
rect 11438 6082 11477 6116
rect 11511 6082 11550 6116
rect 11584 6082 11623 6116
rect 11657 6082 11696 6116
rect 11730 6082 11769 6116
rect 11803 6082 11842 6116
rect 11876 6082 11915 6116
rect 11949 6082 11988 6116
rect 12022 6082 12061 6116
rect 12095 6082 12134 6116
rect 12168 6082 12207 6116
rect 12241 6082 12280 6116
rect 12314 6082 12353 6116
rect 12387 6082 12426 6116
rect 12460 6082 12499 6116
rect 12533 6082 12572 6116
rect 12606 6082 12645 6116
rect 12679 6082 12718 6116
rect 12752 6082 12791 6116
rect 12825 6082 12864 6116
rect 12898 6082 12937 6116
rect 12971 6082 13010 6116
rect 13044 6082 13083 6116
rect 13117 6082 13156 6116
rect 13190 6082 13229 6116
rect 13263 6082 13302 6116
rect 13336 6082 13375 6116
rect 13409 6082 13448 6116
rect 13482 6082 13521 6116
rect 13555 6082 13594 6116
rect 13628 6082 13667 6116
rect 13701 6114 13732 6116
rect 13701 6083 13739 6114
rect 13701 6082 13773 6083
rect 11146 6080 13773 6082
rect 11146 6046 11153 6080
rect 11187 6046 11221 6080
rect 11255 6046 11289 6080
rect 11323 6046 11357 6080
rect 11391 6046 11425 6080
rect 11459 6046 11493 6080
rect 11527 6046 11561 6080
rect 11595 6046 11629 6080
rect 11663 6046 11697 6080
rect 11731 6046 11765 6080
rect 11799 6046 11833 6080
rect 11867 6046 11901 6080
rect 11935 6046 11969 6080
rect 12003 6046 12037 6080
rect 12071 6046 12105 6080
rect 12139 6046 12173 6080
rect 12207 6046 12241 6080
rect 12275 6046 12309 6080
rect 12343 6046 12377 6080
rect 12411 6046 12445 6080
rect 12479 6046 12513 6080
rect 12547 6046 12581 6080
rect 12615 6046 12649 6080
rect 12683 6046 12717 6080
rect 12751 6046 12785 6080
rect 12819 6046 12853 6080
rect 12887 6046 12921 6080
rect 12955 6046 12989 6080
rect 13023 6046 13057 6080
rect 13091 6046 13125 6080
rect 13159 6046 13193 6080
rect 13227 6046 13261 6080
rect 13295 6046 13329 6080
rect 13363 6046 13397 6080
rect 13431 6046 13465 6080
rect 13499 6046 13533 6080
rect 13567 6046 13601 6080
rect 13635 6046 13773 6080
rect 11146 6044 13773 6046
rect 11146 6010 11185 6044
rect 11219 6010 11258 6044
rect 11292 6010 11331 6044
rect 11365 6010 11404 6044
rect 11438 6010 11477 6044
rect 11511 6010 11550 6044
rect 11584 6010 11623 6044
rect 11657 6010 11696 6044
rect 11730 6010 11769 6044
rect 11803 6010 11842 6044
rect 11876 6010 11915 6044
rect 11949 6010 11988 6044
rect 12022 6010 12061 6044
rect 12095 6010 12134 6044
rect 12168 6010 12207 6044
rect 12241 6010 12280 6044
rect 12314 6010 12353 6044
rect 12387 6010 12426 6044
rect 12460 6010 12499 6044
rect 12533 6010 12572 6044
rect 12606 6010 12645 6044
rect 12679 6010 12718 6044
rect 12752 6010 12791 6044
rect 12825 6010 12864 6044
rect 12898 6010 12937 6044
rect 12971 6010 13010 6044
rect 13044 6010 13083 6044
rect 13117 6010 13156 6044
rect 13190 6010 13229 6044
rect 13263 6010 13302 6044
rect 13336 6010 13375 6044
rect 13409 6010 13448 6044
rect 13482 6010 13521 6044
rect 13555 6010 13594 6044
rect 13628 6010 13667 6044
rect 13701 6010 13773 6044
rect 10464 5950 13773 6010
rect 10464 5916 10473 5950
rect 10507 5916 10546 5950
rect 10580 5916 10619 5950
rect 10653 5916 10692 5950
rect 10726 5916 10765 5950
rect 10799 5916 10838 5950
rect 10872 5916 10911 5950
rect 10945 5916 10984 5950
rect 11018 5916 11057 5950
rect 11091 5916 11130 5950
rect 11164 5916 11203 5950
rect 11237 5916 11276 5950
rect 11310 5916 11349 5950
rect 11383 5916 11422 5950
rect 11456 5916 11495 5950
rect 11529 5916 11568 5950
rect 11602 5916 11641 5950
rect 11675 5916 11714 5950
rect 11748 5916 11787 5950
rect 11821 5916 11860 5950
rect 11894 5916 11933 5950
rect 11967 5916 12005 5950
rect 12039 5916 12077 5950
rect 12111 5916 12149 5950
rect 12183 5916 12221 5950
rect 12255 5916 12293 5950
rect 12327 5916 12365 5950
rect 12399 5916 12437 5950
rect 12471 5916 12509 5950
rect 12543 5916 12581 5950
rect 12615 5916 12653 5950
rect 12687 5916 12725 5950
rect 12759 5916 12797 5950
rect 12831 5916 12869 5950
rect 12903 5916 12941 5950
rect 12975 5916 13013 5950
rect 13047 5916 13085 5950
rect 13119 5916 13157 5950
rect 13191 5916 13229 5950
rect 13263 5916 13301 5950
rect 13335 5916 13373 5950
rect 13407 5916 13445 5950
rect 13479 5916 13517 5950
rect 13551 5916 13589 5950
rect 13623 5916 13661 5950
rect 13695 5916 13733 5950
rect 13767 5916 13773 5950
rect 947 5852 1015 5886
rect 1049 5880 1083 5886
rect 1117 5880 1151 5886
rect 1185 5880 1219 5886
rect 1253 5880 1287 5886
rect 1321 5880 1355 5886
rect 1389 5880 1423 5886
rect 1457 5880 1491 5886
rect 1053 5852 1083 5880
rect 1126 5852 1151 5880
rect 1199 5852 1219 5880
rect 1271 5852 1287 5880
rect 1343 5852 1355 5880
rect 1415 5852 1423 5880
rect 1487 5852 1491 5880
rect 1525 5880 1559 5886
rect 947 5846 1019 5852
rect 1053 5846 1092 5852
rect 1126 5846 1165 5852
rect 1199 5846 1237 5852
rect 1271 5846 1309 5852
rect 1343 5846 1381 5852
rect 1415 5846 1453 5852
rect 1487 5846 1525 5852
rect 1593 5880 1627 5886
rect 1661 5880 1695 5886
rect 1729 5880 1763 5886
rect 1797 5880 1831 5886
rect 1865 5880 1899 5886
rect 1933 5880 1967 5886
rect 2001 5880 2035 5886
rect 2069 5880 2103 5886
rect 1593 5852 1597 5880
rect 1661 5852 1669 5880
rect 1729 5852 1741 5880
rect 1797 5852 1813 5880
rect 1865 5852 1885 5880
rect 1933 5852 1957 5880
rect 2001 5852 2029 5880
rect 2069 5852 2101 5880
rect 2137 5852 2171 5886
rect 2205 5880 2239 5886
rect 2273 5880 2307 5886
rect 2341 5880 2375 5886
rect 2409 5880 2443 5886
rect 2477 5880 2511 5886
rect 2545 5880 2579 5886
rect 2613 5880 2647 5886
rect 2681 5880 2715 5886
rect 2207 5852 2239 5880
rect 2279 5852 2307 5880
rect 2351 5852 2375 5880
rect 2423 5852 2443 5880
rect 2495 5852 2511 5880
rect 2567 5852 2579 5880
rect 2639 5852 2647 5880
rect 2711 5852 2715 5880
rect 2749 5880 2783 5886
rect 1559 5846 1597 5852
rect 1631 5846 1669 5852
rect 1703 5846 1741 5852
rect 1775 5846 1813 5852
rect 1847 5846 1885 5852
rect 1919 5846 1957 5852
rect 1991 5846 2029 5852
rect 2063 5846 2101 5852
rect 2135 5846 2173 5852
rect 2207 5846 2245 5852
rect 2279 5846 2317 5852
rect 2351 5846 2389 5852
rect 2423 5846 2461 5852
rect 2495 5846 2533 5852
rect 2567 5846 2605 5852
rect 2639 5846 2677 5852
rect 2711 5846 2749 5852
rect 2817 5880 2851 5886
rect 2885 5880 2919 5886
rect 2953 5880 2987 5886
rect 3021 5880 3055 5886
rect 3089 5880 3123 5886
rect 3157 5880 3191 5886
rect 3225 5880 3259 5886
rect 3293 5880 3327 5886
rect 2817 5852 2821 5880
rect 2885 5852 2893 5880
rect 2953 5852 2965 5880
rect 3021 5852 3037 5880
rect 3089 5852 3109 5880
rect 3157 5852 3181 5880
rect 3225 5852 3253 5880
rect 3293 5852 3325 5880
rect 3361 5852 3395 5886
rect 3429 5880 3463 5886
rect 3497 5880 3531 5886
rect 3565 5880 3599 5886
rect 3633 5880 3667 5886
rect 3701 5880 3735 5886
rect 3769 5880 3803 5886
rect 3837 5880 3871 5886
rect 3905 5880 3939 5886
rect 3431 5852 3463 5880
rect 3503 5852 3531 5880
rect 3575 5852 3599 5880
rect 3647 5852 3667 5880
rect 3719 5852 3735 5880
rect 3791 5852 3803 5880
rect 3863 5852 3871 5880
rect 3935 5852 3939 5880
rect 3973 5880 4007 5886
rect 2783 5846 2821 5852
rect 2855 5846 2893 5852
rect 2927 5846 2965 5852
rect 2999 5846 3037 5852
rect 3071 5846 3109 5852
rect 3143 5846 3181 5852
rect 3215 5846 3253 5852
rect 3287 5846 3325 5852
rect 3359 5846 3397 5852
rect 3431 5846 3469 5852
rect 3503 5846 3541 5852
rect 3575 5846 3613 5852
rect 3647 5846 3685 5852
rect 3719 5846 3757 5852
rect 3791 5846 3829 5852
rect 3863 5846 3901 5852
rect 3935 5846 3973 5852
rect 4041 5880 4075 5886
rect 4109 5880 4143 5886
rect 4177 5880 4211 5886
rect 4245 5880 4279 5886
rect 4313 5880 4347 5886
rect 4381 5880 4415 5886
rect 4449 5880 4483 5886
rect 4517 5880 4551 5886
rect 4041 5852 4045 5880
rect 4109 5852 4117 5880
rect 4177 5852 4189 5880
rect 4245 5852 4261 5880
rect 4313 5852 4333 5880
rect 4381 5852 4405 5880
rect 4449 5852 4477 5880
rect 4517 5852 4549 5880
rect 4585 5852 4619 5886
rect 4653 5880 4687 5886
rect 4721 5880 4755 5886
rect 4789 5880 4823 5886
rect 4857 5880 4891 5886
rect 4925 5880 4959 5886
rect 4993 5880 5027 5886
rect 5061 5880 5095 5886
rect 5129 5880 5163 5886
rect 4655 5852 4687 5880
rect 4727 5852 4755 5880
rect 4799 5852 4823 5880
rect 4871 5852 4891 5880
rect 4943 5852 4959 5880
rect 5015 5852 5027 5880
rect 5087 5852 5095 5880
rect 5159 5852 5163 5880
rect 5197 5880 5231 5886
rect 4007 5846 4045 5852
rect 4079 5846 4117 5852
rect 4151 5846 4189 5852
rect 4223 5846 4261 5852
rect 4295 5846 4333 5852
rect 4367 5846 4405 5852
rect 4439 5846 4477 5852
rect 4511 5846 4549 5852
rect 4583 5846 4621 5852
rect 4655 5846 4693 5852
rect 4727 5846 4765 5852
rect 4799 5846 4837 5852
rect 4871 5846 4909 5852
rect 4943 5846 4981 5852
rect 5015 5846 5053 5852
rect 5087 5846 5125 5852
rect 5159 5846 5197 5852
rect 5265 5880 5299 5886
rect 5333 5880 5367 5886
rect 5401 5880 5435 5886
rect 5469 5880 5503 5886
rect 5537 5880 5571 5886
rect 5605 5880 5639 5886
rect 5673 5880 5707 5886
rect 5741 5880 5775 5886
rect 5265 5852 5269 5880
rect 5333 5852 5341 5880
rect 5401 5852 5413 5880
rect 5469 5852 5485 5880
rect 5537 5852 5557 5880
rect 5605 5852 5629 5880
rect 5673 5852 5701 5880
rect 5741 5852 5773 5880
rect 5809 5852 5843 5886
rect 5877 5880 5911 5886
rect 5945 5880 5979 5886
rect 6013 5880 6047 5886
rect 6081 5880 6115 5886
rect 6149 5880 6183 5886
rect 6217 5880 6251 5886
rect 6285 5880 6319 5886
rect 6353 5880 6387 5886
rect 5879 5852 5911 5880
rect 5951 5852 5979 5880
rect 6023 5852 6047 5880
rect 6095 5852 6115 5880
rect 6167 5852 6183 5880
rect 6239 5852 6251 5880
rect 6311 5852 6319 5880
rect 6383 5852 6387 5880
rect 6421 5880 6455 5886
rect 5231 5846 5269 5852
rect 5303 5846 5341 5852
rect 5375 5846 5413 5852
rect 5447 5846 5485 5852
rect 5519 5846 5557 5852
rect 5591 5846 5629 5852
rect 5663 5846 5701 5852
rect 5735 5846 5773 5852
rect 5807 5846 5845 5852
rect 5879 5846 5917 5852
rect 5951 5846 5989 5852
rect 6023 5846 6061 5852
rect 6095 5846 6133 5852
rect 6167 5846 6205 5852
rect 6239 5846 6277 5852
rect 6311 5846 6349 5852
rect 6383 5846 6421 5852
rect 6489 5880 6523 5886
rect 6557 5880 6591 5886
rect 6625 5880 6659 5886
rect 6693 5880 6727 5886
rect 6761 5880 6795 5886
rect 6829 5880 6863 5886
rect 6897 5880 6931 5886
rect 6965 5880 6999 5886
rect 6489 5852 6493 5880
rect 6557 5852 6565 5880
rect 6625 5852 6637 5880
rect 6693 5852 6709 5880
rect 6761 5852 6781 5880
rect 6829 5852 6853 5880
rect 6897 5852 6925 5880
rect 6965 5852 6997 5880
rect 7033 5852 7067 5886
rect 7101 5880 7135 5886
rect 7169 5880 7203 5886
rect 7237 5880 7271 5886
rect 7305 5880 7339 5886
rect 7373 5880 7407 5886
rect 7441 5880 7475 5886
rect 7509 5880 7543 5886
rect 7577 5880 7611 5886
rect 7103 5852 7135 5880
rect 7175 5852 7203 5880
rect 7247 5852 7271 5880
rect 7319 5852 7339 5880
rect 7391 5852 7407 5880
rect 7463 5852 7475 5880
rect 7535 5852 7543 5880
rect 7607 5852 7611 5880
rect 7645 5880 7679 5886
rect 6455 5846 6493 5852
rect 6527 5846 6565 5852
rect 6599 5846 6637 5852
rect 6671 5846 6709 5852
rect 6743 5846 6781 5852
rect 6815 5846 6853 5852
rect 6887 5846 6925 5852
rect 6959 5846 6997 5852
rect 7031 5846 7069 5852
rect 7103 5846 7141 5852
rect 7175 5846 7213 5852
rect 7247 5846 7285 5852
rect 7319 5846 7357 5852
rect 7391 5846 7429 5852
rect 7463 5846 7501 5852
rect 7535 5846 7573 5852
rect 7607 5846 7645 5852
rect 7713 5880 7747 5886
rect 7781 5880 7815 5886
rect 7849 5880 7883 5886
rect 7917 5880 7951 5886
rect 7985 5880 8019 5886
rect 8053 5880 8087 5886
rect 8121 5880 8155 5886
rect 8189 5880 8223 5886
rect 7713 5852 7717 5880
rect 7781 5852 7789 5880
rect 7849 5852 7861 5880
rect 7917 5852 7933 5880
rect 7985 5852 8005 5880
rect 8053 5852 8077 5880
rect 8121 5852 8149 5880
rect 8189 5852 8221 5880
rect 8257 5852 8291 5886
rect 8325 5880 8359 5886
rect 8393 5880 8427 5886
rect 8461 5880 8495 5886
rect 8529 5880 8563 5886
rect 8597 5880 8631 5886
rect 8665 5880 8699 5886
rect 8733 5880 8767 5886
rect 8801 5880 8835 5886
rect 8327 5852 8359 5880
rect 8399 5852 8427 5880
rect 8471 5852 8495 5880
rect 8543 5852 8563 5880
rect 8615 5852 8631 5880
rect 8687 5852 8699 5880
rect 8759 5852 8767 5880
rect 8831 5852 8835 5880
rect 8869 5880 8903 5886
rect 7679 5846 7717 5852
rect 7751 5846 7789 5852
rect 7823 5846 7861 5852
rect 7895 5846 7933 5852
rect 7967 5846 8005 5852
rect 8039 5846 8077 5852
rect 8111 5846 8149 5852
rect 8183 5846 8221 5852
rect 8255 5846 8293 5852
rect 8327 5846 8365 5852
rect 8399 5846 8437 5852
rect 8471 5846 8509 5852
rect 8543 5846 8581 5852
rect 8615 5846 8653 5852
rect 8687 5846 8725 5852
rect 8759 5846 8797 5852
rect 8831 5846 8869 5852
rect 8937 5880 8971 5886
rect 9005 5880 9039 5886
rect 9073 5880 9191 5886
rect 8937 5852 8941 5880
rect 9005 5852 9013 5880
rect 9073 5852 9085 5880
rect 8903 5846 8941 5852
rect 8975 5846 9013 5852
rect 9047 5846 9085 5852
rect 9119 5846 9191 5880
rect 10464 5860 13773 5916
rect 10832 5847 10964 5860
rect 10998 5847 11032 5860
rect 790 5752 804 5791
rect 790 5703 804 5718
rect 620 5680 804 5703
rect 620 5646 626 5680
rect 660 5646 698 5680
rect 732 5679 804 5680
rect 732 5646 770 5679
rect 620 5645 770 5646
rect 620 5631 804 5645
rect 654 5607 688 5631
rect 722 5607 804 5631
rect 660 5597 688 5607
rect 732 5606 804 5607
rect 9462 5764 9466 5809
rect 9636 5766 9640 5809
rect 9462 5685 9466 5730
rect 9636 5690 9640 5732
rect 9462 5606 9466 5651
rect 9636 5614 9640 5656
rect 732 5602 770 5606
rect 5700 5602 5739 5606
rect 5773 5602 5812 5606
rect 5846 5602 5885 5606
rect 5919 5602 5958 5606
rect 5992 5602 6031 5606
rect 6065 5602 6104 5606
rect 6138 5602 6177 5606
rect 6211 5602 6250 5606
rect 6284 5602 6323 5606
rect 6357 5602 6396 5606
rect 6430 5602 6469 5606
rect 6503 5602 6542 5606
rect 6576 5602 6615 5606
rect 6649 5602 6688 5606
rect 6722 5602 6761 5606
rect 6795 5602 6834 5606
rect 6868 5602 6907 5606
rect 6941 5602 6980 5606
rect 7014 5602 7053 5606
rect 7087 5602 7126 5606
rect 7160 5602 7199 5606
rect 7233 5602 7272 5606
rect 7306 5602 7345 5606
rect 7379 5602 7418 5606
rect 7452 5602 7491 5606
rect 7525 5602 7564 5606
rect 7598 5602 7637 5606
rect 7671 5602 7710 5606
rect 7744 5602 7783 5606
rect 7817 5602 7856 5606
rect 7890 5602 7929 5606
rect 7963 5602 8002 5606
rect 8036 5602 8075 5606
rect 8109 5602 8148 5606
rect 8182 5602 8221 5606
rect 8255 5602 8294 5606
rect 8328 5602 8367 5606
rect 8401 5602 8440 5606
rect 8474 5602 8513 5606
rect 8547 5602 8586 5606
rect 8620 5602 8659 5606
rect 8693 5602 8732 5606
rect 8766 5602 8805 5606
rect 8839 5602 8878 5606
rect 8912 5602 8951 5606
rect 8985 5602 9024 5606
rect 9058 5602 9097 5606
rect 9131 5602 9170 5606
rect 9204 5602 9243 5606
rect 9277 5602 9316 5606
rect 9350 5602 9389 5606
rect 9423 5602 9462 5606
rect 620 5573 626 5597
rect 660 5573 698 5597
rect 732 5573 756 5602
rect 620 5563 756 5573
rect 654 5534 756 5563
rect 9426 5572 9462 5602
rect 9426 5568 9466 5572
rect 9426 5534 9534 5568
rect 9636 5538 9640 5580
rect 620 5500 626 5529
rect 660 5500 688 5534
rect 620 5432 688 5500
rect 9495 5500 9534 5534
rect 9636 5500 9640 5504
rect 9494 5466 9640 5500
rect 9494 5462 9528 5466
rect 9562 5462 9640 5466
rect 9495 5432 9528 5462
rect 626 5428 698 5432
rect 5772 5428 5811 5432
rect 5845 5428 5884 5432
rect 5918 5428 5957 5432
rect 5991 5428 6030 5432
rect 6064 5428 6103 5432
rect 6137 5428 6176 5432
rect 6210 5428 6249 5432
rect 6283 5428 6322 5432
rect 6356 5428 6395 5432
rect 6429 5428 6468 5432
rect 6502 5428 6541 5432
rect 6575 5428 6614 5432
rect 6648 5428 6687 5432
rect 6721 5428 6760 5432
rect 6794 5428 6833 5432
rect 6867 5428 6906 5432
rect 6940 5428 6979 5432
rect 7013 5428 7052 5432
rect 7086 5428 7125 5432
rect 7159 5428 7198 5432
rect 7232 5428 7271 5432
rect 7305 5428 7344 5432
rect 7378 5428 7417 5432
rect 7451 5428 7490 5432
rect 7524 5428 7563 5432
rect 7597 5428 7636 5432
rect 7670 5428 7709 5432
rect 7743 5428 7782 5432
rect 7816 5428 7855 5432
rect 7889 5428 7928 5432
rect 7962 5428 8001 5432
rect 8035 5428 8074 5432
rect 8108 5428 8147 5432
rect 8181 5428 8220 5432
rect 8254 5428 8293 5432
rect 8327 5428 8366 5432
rect 8400 5428 8439 5432
rect 8473 5428 8512 5432
rect 8546 5428 8585 5432
rect 8619 5428 8658 5432
rect 8692 5428 8731 5432
rect 8765 5428 8804 5432
rect 8838 5428 8877 5432
rect 8911 5428 8950 5432
rect 8984 5428 9023 5432
rect 9057 5428 9096 5432
rect 9130 5428 9169 5432
rect 9203 5428 9242 5432
rect 9276 5428 9315 5432
rect 9349 5428 9388 5432
rect 9422 5428 9461 5432
rect 9495 5428 9534 5432
rect 9568 5428 9640 5462
rect 10832 5792 10904 5847
rect 10832 5775 10836 5792
rect 14058 5775 14126 5860
rect 10832 5699 10836 5741
rect 10938 5724 10976 5741
rect 13990 5703 14020 5758
rect 12522 5669 12561 5690
rect 12595 5669 12634 5690
rect 12668 5669 12707 5690
rect 12741 5669 12780 5690
rect 12814 5669 12853 5690
rect 12887 5669 12926 5690
rect 12960 5669 12999 5690
rect 13033 5669 13072 5690
rect 13106 5669 13145 5690
rect 13179 5669 13218 5690
rect 13252 5669 13291 5690
rect 13325 5669 13364 5690
rect 13398 5669 13437 5690
rect 13471 5669 13510 5690
rect 13544 5669 13583 5690
rect 13617 5669 13656 5690
rect 13690 5669 13729 5690
rect 13763 5669 13802 5690
rect 13836 5669 13875 5690
rect 13909 5669 13948 5690
rect 10832 5623 10836 5665
rect 11006 5628 11010 5669
rect 10832 5548 10836 5589
rect 11006 5553 11010 5594
rect 10832 5473 10836 5514
rect 11006 5478 11010 5519
rect 10832 5398 10836 5439
rect 11006 5403 11010 5444
rect 10832 5323 10836 5364
rect 11006 5328 11010 5369
rect 10832 5248 10836 5289
rect 11006 5253 11010 5294
rect 10832 5173 10836 5214
rect 11006 5178 11010 5219
rect 10832 5098 10836 5139
rect 11006 5103 11010 5144
rect 10832 5023 10836 5064
rect 11006 5028 11010 5069
rect 10832 4948 10836 4989
rect 11006 4953 11010 4994
rect 10832 4873 10836 4914
rect 11006 4878 11010 4919
rect 10832 4798 10836 4839
rect 11006 4803 11010 4844
rect 10832 4723 10836 4764
rect 11006 4728 11010 4769
rect 11364 5537 12562 5543
rect 11364 5503 11468 5537
rect 11502 5503 11536 5537
rect 11574 5503 11604 5537
rect 11646 5503 11672 5537
rect 11718 5503 11740 5537
rect 11790 5503 11808 5537
rect 11862 5503 11876 5537
rect 11934 5503 11944 5537
rect 12006 5503 12012 5537
rect 12078 5503 12080 5537
rect 12114 5503 12116 5537
rect 12182 5503 12188 5537
rect 12250 5503 12260 5537
rect 12318 5503 12332 5537
rect 12386 5503 12404 5537
rect 12454 5503 12476 5537
rect 12522 5503 12562 5537
rect 11364 5497 12562 5503
rect 11364 5462 11410 5497
rect 11364 5415 11370 5462
rect 11404 5415 11410 5462
rect 11364 5390 11410 5415
rect 11364 5347 11370 5390
rect 11404 5347 11410 5390
rect 11364 5318 11410 5347
rect 11364 5279 11370 5318
rect 11404 5279 11410 5318
rect 12516 5462 12562 5497
rect 12516 5415 12522 5462
rect 12556 5415 12562 5462
rect 12516 5390 12562 5415
rect 12516 5347 12522 5390
rect 12556 5347 12562 5390
rect 12516 5318 12562 5347
rect 11364 5246 11410 5279
rect 11364 5211 11370 5246
rect 11404 5211 11410 5246
rect 11364 5177 11410 5211
rect 11364 5140 11370 5177
rect 11404 5140 11410 5177
rect 11364 5109 11410 5140
rect 11364 5068 11370 5109
rect 11404 5068 11410 5109
rect 11364 5041 11410 5068
rect 11364 4996 11370 5041
rect 11404 4996 11410 5041
rect 11364 4973 11410 4996
rect 11364 4924 11370 4973
rect 11404 4924 11410 4973
rect 11364 4905 11410 4924
rect 11364 4852 11370 4905
rect 11404 4852 11410 4905
rect 11364 4837 11410 4852
rect 11364 4780 11370 4837
rect 11404 4780 11410 4837
rect 11364 4769 11410 4780
rect 11364 4708 11370 4769
rect 11404 4708 11410 4769
rect 11364 4701 11410 4708
rect 11364 4696 11370 4701
rect 10832 4670 10836 4689
rect 10832 4648 10904 4670
rect 11006 4653 11010 4694
rect 2330 4576 2402 4648
rect 10428 4616 10467 4648
rect 10501 4616 10540 4648
rect 10574 4616 10613 4648
rect 10647 4616 10686 4648
rect 10720 4616 10759 4648
rect 10793 4616 10832 4648
rect 10866 4616 10904 4648
rect 2364 4548 2402 4576
rect 10870 4602 10904 4616
rect 11006 4602 11010 4619
rect 10870 4578 11010 4602
rect 10870 4576 10976 4578
rect 10870 4548 10904 4576
rect 10938 4568 10976 4576
rect 2330 4503 2334 4542
rect 2436 4514 2472 4542
rect 2436 4480 2474 4514
rect 10938 4534 10972 4568
rect 11006 4534 11010 4544
rect 10938 4470 11010 4534
rect 11404 4696 11410 4701
rect 11511 5246 11557 5286
rect 11511 5212 11517 5246
rect 11551 5212 11557 5246
rect 11511 5174 11557 5212
rect 11511 5140 11517 5174
rect 11551 5140 11557 5174
rect 11511 5102 11557 5140
rect 11511 5068 11517 5102
rect 11551 5068 11557 5102
rect 11511 5030 11557 5068
rect 11511 4996 11517 5030
rect 11551 4996 11557 5030
rect 11511 4958 11557 4996
rect 11511 4924 11517 4958
rect 11551 4924 11557 4958
rect 11511 4886 11557 4924
rect 11511 4852 11517 4886
rect 11551 4852 11557 4886
rect 11511 4814 11557 4852
rect 11511 4780 11517 4814
rect 11551 4780 11557 4814
rect 11511 4742 11557 4780
rect 11511 4708 11517 4742
rect 11551 4708 11557 4742
rect 11511 4696 11557 4708
rect 12370 5246 12416 5286
rect 12370 5212 12376 5246
rect 12410 5212 12416 5246
rect 12370 5174 12416 5212
rect 12370 5140 12376 5174
rect 12410 5140 12416 5174
rect 12370 5102 12416 5140
rect 12370 5068 12376 5102
rect 12410 5068 12416 5102
rect 12370 5030 12416 5068
rect 12370 4996 12376 5030
rect 12410 4996 12416 5030
rect 12370 4958 12416 4996
rect 12370 4924 12376 4958
rect 12410 4924 12416 4958
rect 12370 4886 12416 4924
rect 12370 4852 12376 4886
rect 12410 4852 12416 4886
rect 12370 4814 12416 4852
rect 12370 4780 12376 4814
rect 12410 4780 12416 4814
rect 12370 4742 12416 4780
rect 12370 4708 12376 4742
rect 12410 4708 12416 4742
rect 12370 4696 12416 4708
rect 12516 5279 12522 5318
rect 12556 5279 12562 5318
rect 12516 5246 12562 5279
rect 12516 5211 12522 5246
rect 12556 5211 12562 5246
rect 12516 5177 12562 5211
rect 12516 5140 12522 5177
rect 12556 5140 12562 5177
rect 12516 5109 12562 5140
rect 12516 5068 12522 5109
rect 12556 5068 12562 5109
rect 12516 5041 12562 5068
rect 12516 4996 12522 5041
rect 12556 4996 12562 5041
rect 12516 4973 12562 4996
rect 12516 4924 12522 4973
rect 12556 4924 12562 4973
rect 12516 4905 12562 4924
rect 12516 4852 12522 4905
rect 12556 4852 12562 4905
rect 12516 4837 12562 4852
rect 12516 4780 12522 4837
rect 12556 4780 12562 4837
rect 12516 4769 12562 4780
rect 12516 4708 12522 4769
rect 12556 4708 12562 4769
rect 12516 4701 12562 4708
rect 12516 4696 12522 4701
rect 11370 4633 11404 4667
rect 11370 4565 11404 4599
rect 11370 4497 11404 4531
rect 2330 4430 2334 4469
rect 2504 4446 2540 4470
rect 10938 4446 11006 4470
rect 2504 4431 2508 4446
rect 2330 4357 2334 4396
rect 2504 4358 2508 4397
rect 2330 4284 2334 4323
rect 2504 4285 2508 4324
rect 11370 4429 11404 4463
rect 11370 4361 11404 4395
rect 12556 4696 12562 4701
rect 13948 5414 13956 5453
rect 13948 5341 13956 5380
rect 13948 5268 13956 5307
rect 13948 5195 13956 5234
rect 13948 5122 13956 5161
rect 13948 5049 13956 5088
rect 13948 4976 13956 5015
rect 13948 4903 13956 4942
rect 13948 4830 13956 4869
rect 13948 4757 13956 4796
rect 12522 4633 12556 4667
rect 12522 4565 12556 4599
rect 12522 4497 12556 4531
rect 13948 4684 13956 4723
rect 13948 4611 13956 4650
rect 13948 4538 13956 4577
rect 12522 4429 12556 4463
rect 11563 4387 12363 4393
rect 11563 4353 11597 4387
rect 11663 4353 11669 4387
rect 11731 4353 11741 4387
rect 11799 4353 11813 4387
rect 11867 4353 11885 4387
rect 11935 4353 11957 4387
rect 12003 4353 12029 4387
rect 12071 4353 12101 4387
rect 12139 4353 12173 4387
rect 12207 4353 12241 4387
rect 12279 4353 12309 4387
rect 12351 4353 12363 4387
rect 11563 4347 12363 4353
rect 12522 4361 12556 4395
rect 11370 4293 11404 4327
rect 12522 4293 12556 4327
rect 2330 4211 2334 4250
rect 2504 4212 2508 4251
rect 2330 4138 2334 4177
rect 2504 4139 2508 4178
rect 2330 4065 2334 4104
rect 2504 4066 2508 4105
rect 2330 3992 2334 4031
rect 2504 3993 2508 4032
rect 2330 3919 2334 3958
rect 2504 3920 2508 3959
rect 2330 3846 2334 3885
rect 2504 3847 2508 3886
rect 2330 3773 2334 3812
rect 2504 3774 2508 3813
rect 2330 3700 2334 3739
rect 2504 3701 2508 3740
rect 2330 3627 2334 3666
rect 2504 3628 2508 3667
rect 2330 3554 2334 3593
rect 2504 3555 2508 3594
rect 2330 3481 2334 3520
rect 2504 3482 2508 3521
rect 2330 3408 2334 3447
rect 2504 3409 2508 3448
rect 2330 3335 2334 3374
rect 2504 3336 2508 3375
rect 2330 3262 2334 3301
rect 2504 3263 2508 3302
rect 13953 4172 13956 4213
rect 13953 4097 13956 4138
rect 13953 4022 13956 4063
rect 13953 3947 13956 3988
rect 13953 3872 13956 3913
rect 13953 3797 13956 3838
rect 13953 3722 13956 3763
rect 13953 3647 13956 3688
rect 13953 3571 13956 3613
rect 13953 3495 13956 3537
rect 13953 3419 13956 3461
rect 13953 3343 13956 3385
rect 13953 3267 13956 3309
rect 2330 3189 2334 3228
rect 2504 3190 2508 3229
rect 2330 3116 2334 3155
rect 2504 3117 2508 3156
rect 2330 3043 2334 3082
rect 2504 3044 2508 3083
rect 2330 2970 2334 3009
rect 2504 2971 2508 3010
rect 2504 2898 2508 2937
rect 13953 2908 13956 2949
rect 13953 2833 13956 2874
rect 13953 2758 13956 2799
rect 13953 2683 13956 2724
rect 13953 2608 13956 2649
rect 13953 2533 13956 2574
rect 13953 2458 13956 2499
rect 13953 2383 13956 2424
rect 13953 2307 13956 2349
rect 13953 2231 13956 2273
rect 13953 2155 13956 2197
rect 13953 2079 13956 2121
rect 13953 2003 13956 2045
rect 13953 1708 13956 1749
rect 13953 1633 13956 1674
rect 13953 1558 13956 1599
rect 13953 1483 13956 1524
rect 13953 1408 13956 1449
rect 13953 1333 13956 1374
rect 13953 1258 13956 1299
rect 13953 1183 13956 1224
rect 13953 1107 13956 1149
rect 13953 1031 13956 1073
rect 13953 955 13956 997
rect 13953 879 13956 921
rect 13953 803 13956 845
rect 13952 466 13956 520
rect 14126 472 14130 520
rect 13952 378 13956 432
rect 14126 389 14130 438
rect 2508 374 2547 378
rect 2581 374 2620 378
rect 2654 374 2693 378
rect 2727 374 2766 378
rect 2800 374 2839 378
rect 2873 374 2912 378
rect 2946 374 2985 378
rect 3019 374 3058 378
rect 3092 374 3131 378
rect 3165 374 3204 378
rect 3238 374 3277 378
rect 3311 374 3350 378
rect 3384 374 3423 378
rect 3457 374 3496 378
rect 3530 374 3569 378
rect 3603 374 3642 378
rect 3676 374 3715 378
rect 3749 374 3788 378
rect 3822 374 3861 378
rect 3895 374 3934 378
rect 3968 374 4007 378
rect 4041 374 4080 378
rect 4114 374 4153 378
rect 4187 374 4226 378
rect 4260 374 4299 378
rect 4333 374 4372 378
rect 4406 374 4445 378
rect 4479 374 4518 378
rect 4552 374 4591 378
rect 4625 374 4664 378
rect 2436 306 2470 344
rect 13986 306 14024 340
rect 14126 306 14130 355
rect 2330 200 2402 272
rect 2436 200 2475 204
rect 2509 200 2548 204
rect 2582 200 2621 204
rect 2655 200 2694 204
rect 2728 200 2767 204
rect 2801 200 2840 204
rect 2874 200 2913 204
rect 2947 200 2986 204
rect 3020 200 3059 204
rect 3093 200 3132 204
rect 3166 200 3205 204
rect 3239 200 3278 204
rect 3312 200 3351 204
rect 3385 200 3424 204
rect 3458 200 3497 204
rect 3531 200 3570 204
rect 3604 200 3643 204
rect 3677 200 3716 204
rect 3750 200 3789 204
rect 3823 200 3862 204
rect 3896 200 3935 204
rect 3969 200 4008 204
rect 4042 200 4081 204
rect 4115 200 4154 204
rect 4188 200 4227 204
rect 4261 200 4300 204
rect 4334 200 4373 204
rect 4407 200 4446 204
rect 4480 200 4519 204
rect 4553 200 4592 204
rect 14058 200 14130 272
<< viali >>
rect 1902 39905 1936 39939
rect 1975 39933 2009 39939
rect 2048 39933 2082 39939
rect 2121 39933 2155 39939
rect 2194 39933 2228 39939
rect 2267 39933 2301 39939
rect 2340 39933 2374 39939
rect 2413 39933 2447 39939
rect 2486 39933 2520 39939
rect 2559 39933 2593 39939
rect 2632 39933 2666 39939
rect 2705 39933 2739 39939
rect 2778 39933 2812 39939
rect 2851 39933 2885 39939
rect 2924 39933 2958 39939
rect 2997 39933 3031 39939
rect 3070 39933 3104 39939
rect 3143 39933 3177 39939
rect 3216 39933 3250 39939
rect 3289 39933 3323 39939
rect 3362 39933 3396 39939
rect 3435 39933 3469 39939
rect 3508 39933 3542 39939
rect 3581 39933 3615 39939
rect 3654 39933 3688 39939
rect 3727 39933 3761 39939
rect 3800 39933 3834 39939
rect 3873 39933 3907 39939
rect 3946 39933 3980 39939
rect 4019 39933 4053 39939
rect 4092 39933 4126 39939
rect 4165 39933 4199 39939
rect 4238 39933 4272 39939
rect 4311 39933 4345 39939
rect 4384 39933 4418 39939
rect 4457 39933 4491 39939
rect 4530 39933 4564 39939
rect 4603 39933 4637 39939
rect 4676 39933 4710 39939
rect 4749 39933 4783 39939
rect 4822 39933 4856 39939
rect 4895 39933 4929 39939
rect 4968 39933 5002 39939
rect 5041 39933 5075 39939
rect 5114 39933 5148 39939
rect 5187 39933 5221 39939
rect 5260 39933 5294 39939
rect 5333 39933 5367 39939
rect 5406 39933 5440 39939
rect 5479 39933 5513 39939
rect 5552 39933 5586 39939
rect 5625 39933 5659 39939
rect 5698 39933 5732 39939
rect 5771 39933 5805 39939
rect 5844 39933 5878 39939
rect 5917 39933 5951 39939
rect 5990 39933 6024 39939
rect 6063 39933 6097 39939
rect 6136 39933 6170 39939
rect 6209 39933 6243 39939
rect 6282 39933 6316 39939
rect 6355 39933 6389 39939
rect 6428 39933 6462 39939
rect 6501 39933 6535 39939
rect 6574 39933 6608 39939
rect 6647 39933 13953 39939
rect 1975 39905 1983 39933
rect 1983 39905 2009 39933
rect 2048 39905 2082 39933
rect 2121 39905 2155 39933
rect 2194 39905 2228 39933
rect 2267 39905 2301 39933
rect 2340 39905 2374 39933
rect 2413 39905 2447 39933
rect 2486 39905 2520 39933
rect 2559 39905 2593 39933
rect 2632 39905 2666 39933
rect 2705 39905 2739 39933
rect 2778 39905 2812 39933
rect 2851 39905 2885 39933
rect 2924 39905 2958 39933
rect 2997 39905 3031 39933
rect 3070 39905 3104 39933
rect 3143 39905 3177 39933
rect 3216 39905 3250 39933
rect 3289 39905 3323 39933
rect 3362 39905 3396 39933
rect 3435 39905 3469 39933
rect 3508 39905 3542 39933
rect 3581 39905 3615 39933
rect 3654 39905 3688 39933
rect 3727 39905 3761 39933
rect 3800 39905 3834 39933
rect 3873 39905 3907 39933
rect 3946 39905 3980 39933
rect 4019 39905 4053 39933
rect 4092 39905 4126 39933
rect 4165 39905 4199 39933
rect 4238 39905 4272 39933
rect 4311 39905 4345 39933
rect 4384 39905 4418 39933
rect 4457 39905 4491 39933
rect 4530 39905 4564 39933
rect 4603 39905 4637 39933
rect 4676 39905 4710 39933
rect 4749 39905 4783 39933
rect 4822 39905 4856 39933
rect 4895 39905 4929 39933
rect 4968 39905 5002 39933
rect 5041 39905 5075 39933
rect 5114 39905 5148 39933
rect 5187 39905 5221 39933
rect 5260 39905 5294 39933
rect 5333 39905 5367 39933
rect 5406 39905 5440 39933
rect 5479 39905 5513 39933
rect 5552 39905 5586 39933
rect 5625 39905 5659 39933
rect 5698 39905 5732 39933
rect 5771 39905 5805 39933
rect 5844 39905 5878 39933
rect 5917 39905 5951 39933
rect 5990 39905 6024 39933
rect 6063 39905 6097 39933
rect 6136 39905 6170 39933
rect 6209 39905 6243 39933
rect 6282 39905 6316 39933
rect 6355 39905 6389 39933
rect 6428 39905 6462 39933
rect 6501 39905 6535 39933
rect 6574 39905 6608 39933
rect 1830 39865 1936 39867
rect 1830 35873 1834 39865
rect 1834 39795 1936 39865
rect 1975 39833 2009 39867
rect 2048 39833 2082 39867
rect 2121 39833 2155 39867
rect 2194 39833 2228 39867
rect 2267 39833 2301 39867
rect 2340 39833 2374 39867
rect 2413 39833 2447 39867
rect 2486 39833 2520 39867
rect 2559 39833 2593 39867
rect 2632 39833 2666 39867
rect 2705 39833 2739 39867
rect 2778 39833 2812 39867
rect 2851 39833 2885 39867
rect 2924 39833 2958 39867
rect 2997 39833 3031 39867
rect 3070 39833 3104 39867
rect 3143 39833 3177 39867
rect 3216 39833 3250 39867
rect 3289 39833 3323 39867
rect 3362 39833 3396 39867
rect 3435 39833 3469 39867
rect 3508 39833 3542 39867
rect 3581 39833 3615 39867
rect 3654 39833 3688 39867
rect 3727 39833 3761 39867
rect 3800 39833 3834 39867
rect 3873 39833 3907 39867
rect 3946 39833 3980 39867
rect 4019 39833 4053 39867
rect 4092 39833 4126 39867
rect 4165 39833 4199 39867
rect 4238 39833 4272 39867
rect 4311 39833 4345 39867
rect 4384 39833 4418 39867
rect 4457 39833 4491 39867
rect 4530 39833 4564 39867
rect 4603 39833 4637 39867
rect 4676 39833 4710 39867
rect 4749 39833 4783 39867
rect 4822 39833 4856 39867
rect 4895 39833 4929 39867
rect 4968 39833 5002 39867
rect 5041 39833 5075 39867
rect 5114 39833 5148 39867
rect 5187 39833 5221 39867
rect 5260 39833 5294 39867
rect 5333 39833 5367 39867
rect 5406 39833 5440 39867
rect 5479 39833 5513 39867
rect 5552 39833 5586 39867
rect 5625 39833 5659 39867
rect 5698 39833 5732 39867
rect 5771 39833 5805 39867
rect 5844 39833 5878 39867
rect 5917 39833 5951 39867
rect 5990 39833 6024 39867
rect 6063 39833 6097 39867
rect 6136 39833 6170 39867
rect 6209 39833 6243 39867
rect 6282 39833 6316 39867
rect 6355 39833 6389 39867
rect 6428 39833 6462 39867
rect 6501 39833 6535 39867
rect 6574 39833 6608 39867
rect 6647 39833 13951 39933
rect 13951 39833 13953 39933
rect 13991 39833 14025 39867
rect 14449 39842 14483 39876
rect 14521 39842 14555 39876
rect 1834 39729 2004 39795
rect 2004 39729 2008 39795
rect 2047 39761 2081 39795
rect 2120 39763 2154 39795
rect 2120 39761 2153 39763
rect 2153 39761 2154 39763
rect 2193 39761 2227 39795
rect 2266 39761 2300 39795
rect 2339 39761 2373 39795
rect 2412 39761 2446 39795
rect 2485 39761 2519 39795
rect 2558 39761 2592 39795
rect 2631 39761 2665 39795
rect 2704 39761 2738 39795
rect 2777 39761 2811 39795
rect 2850 39761 2884 39795
rect 2923 39761 2957 39795
rect 2996 39761 3030 39795
rect 3069 39761 3103 39795
rect 3142 39761 3176 39795
rect 3215 39761 3249 39795
rect 3288 39761 3322 39795
rect 3361 39761 3395 39795
rect 3434 39761 3468 39795
rect 3507 39761 3541 39795
rect 3580 39761 3614 39795
rect 3653 39761 3687 39795
rect 3726 39761 3760 39795
rect 3799 39761 3833 39795
rect 3872 39761 3906 39795
rect 3945 39761 3979 39795
rect 4018 39761 4052 39795
rect 4091 39761 4125 39795
rect 4164 39761 4198 39795
rect 4237 39761 4271 39795
rect 4310 39761 4344 39795
rect 4383 39761 4417 39795
rect 4456 39761 4490 39795
rect 4529 39761 4563 39795
rect 4602 39761 4636 39795
rect 4675 39761 4709 39795
rect 4748 39761 4782 39795
rect 4821 39761 4855 39795
rect 4894 39761 4928 39795
rect 4967 39761 5001 39795
rect 5040 39761 5074 39795
rect 5113 39761 5147 39795
rect 5186 39761 5220 39795
rect 5259 39761 5293 39795
rect 5332 39761 5366 39795
rect 5405 39761 5439 39795
rect 5478 39761 5512 39795
rect 5551 39761 5585 39795
rect 5624 39761 5658 39795
rect 5697 39761 5731 39795
rect 5770 39761 5804 39795
rect 5843 39761 5877 39795
rect 5916 39761 5950 39795
rect 5989 39761 6023 39795
rect 6062 39761 6096 39795
rect 6135 39761 6169 39795
rect 6208 39761 6242 39795
rect 6281 39761 6315 39795
rect 6354 39761 6388 39795
rect 6427 39761 6461 39795
rect 6500 39761 6534 39795
rect 6573 39761 6607 39795
rect 6646 39761 6680 39795
rect 6719 39763 13881 39833
rect 6719 39761 13815 39763
rect 13815 39761 13881 39763
rect 1834 39723 2008 39729
rect 1834 35873 2072 39723
rect 2072 35873 2080 39723
rect 2119 39689 2153 39723
rect 2192 39695 2226 39723
rect 2265 39695 2299 39723
rect 2338 39695 2372 39723
rect 2411 39695 2445 39723
rect 2484 39695 2518 39723
rect 2557 39695 2591 39723
rect 2630 39695 2664 39723
rect 2703 39695 2737 39723
rect 2776 39695 2810 39723
rect 2849 39695 2883 39723
rect 2922 39695 2956 39723
rect 2995 39695 3029 39723
rect 3068 39695 3102 39723
rect 3141 39695 3175 39723
rect 3214 39695 3248 39723
rect 3287 39695 3321 39723
rect 3360 39695 3394 39723
rect 3433 39695 3467 39723
rect 3506 39695 3540 39723
rect 3579 39695 3613 39723
rect 3652 39695 3686 39723
rect 3725 39695 3759 39723
rect 3798 39695 3832 39723
rect 3871 39695 3905 39723
rect 3944 39695 3978 39723
rect 4017 39695 4051 39723
rect 4090 39695 4124 39723
rect 4163 39695 4197 39723
rect 4236 39695 4270 39723
rect 4309 39695 4343 39723
rect 4382 39695 4416 39723
rect 4455 39695 4489 39723
rect 4528 39695 4562 39723
rect 4601 39695 4635 39723
rect 4674 39695 4708 39723
rect 4747 39695 4781 39723
rect 4820 39695 4854 39723
rect 4893 39695 4927 39723
rect 4966 39695 5000 39723
rect 5039 39695 5073 39723
rect 5112 39695 5146 39723
rect 5185 39695 5219 39723
rect 5258 39695 5292 39723
rect 5331 39695 5365 39723
rect 5404 39695 5438 39723
rect 5477 39695 5511 39723
rect 5550 39695 5584 39723
rect 5623 39695 5657 39723
rect 5696 39695 5730 39723
rect 5769 39695 5803 39723
rect 5842 39695 5876 39723
rect 5915 39695 5949 39723
rect 5988 39695 6022 39723
rect 6061 39695 6095 39723
rect 6134 39695 6168 39723
rect 6207 39695 6241 39723
rect 6280 39695 6314 39723
rect 6353 39695 6387 39723
rect 6426 39695 6460 39723
rect 6499 39695 6533 39723
rect 6572 39695 6606 39723
rect 6645 39695 6679 39723
rect 6718 39695 6752 39723
rect 6791 39695 13809 39761
rect 13919 39760 13953 39794
rect 13991 39778 14019 39794
rect 14019 39778 14025 39794
rect 13991 39760 14025 39778
rect 2192 39689 2226 39695
rect 2265 39689 2299 39695
rect 2338 39689 2372 39695
rect 2411 39689 2445 39695
rect 2484 39689 2518 39695
rect 2557 39689 2591 39695
rect 2630 39689 2664 39695
rect 2703 39689 2737 39695
rect 2776 39689 2810 39695
rect 2849 39689 2883 39695
rect 2922 39689 2956 39695
rect 2995 39689 3029 39695
rect 3068 39689 3102 39695
rect 3141 39689 3175 39695
rect 3214 39689 3248 39695
rect 3287 39689 3321 39695
rect 3360 39689 3394 39695
rect 3433 39689 3467 39695
rect 3506 39689 3540 39695
rect 3579 39689 3613 39695
rect 3652 39689 3686 39695
rect 3725 39689 3759 39695
rect 3798 39689 3832 39695
rect 3871 39689 3905 39695
rect 3944 39689 3978 39695
rect 4017 39689 4051 39695
rect 4090 39689 4124 39695
rect 4163 39689 4197 39695
rect 4236 39689 4270 39695
rect 4309 39689 4343 39695
rect 4382 39689 4416 39695
rect 4455 39689 4489 39695
rect 4528 39689 4562 39695
rect 4601 39689 4635 39695
rect 4674 39689 4708 39695
rect 4747 39689 4781 39695
rect 4820 39689 4854 39695
rect 4893 39689 4927 39695
rect 4966 39689 5000 39695
rect 5039 39689 5073 39695
rect 5112 39689 5146 39695
rect 5185 39689 5219 39695
rect 5258 39689 5292 39695
rect 5331 39689 5365 39695
rect 5404 39689 5438 39695
rect 5477 39689 5511 39695
rect 5550 39689 5584 39695
rect 5623 39689 5657 39695
rect 5696 39689 5730 39695
rect 5769 39689 5803 39695
rect 5842 39689 5876 39695
rect 5915 39689 5949 39695
rect 5988 39689 6022 39695
rect 6061 39689 6095 39695
rect 6134 39689 6168 39695
rect 6207 39689 6241 39695
rect 6280 39689 6314 39695
rect 6353 39689 6387 39695
rect 6426 39689 6460 39695
rect 6499 39689 6533 39695
rect 6572 39689 6606 39695
rect 6645 39689 6679 39695
rect 6718 39689 6752 39695
rect 6791 39689 13809 39695
rect 13847 39688 13881 39722
rect 13919 39687 13953 39721
rect 13991 39687 14019 39721
rect 14019 39687 14025 39721
rect 13775 39616 13809 39650
rect 13847 39615 13849 39649
rect 13849 39615 13881 39649
rect 13919 39614 13953 39648
rect 13991 39614 14019 39648
rect 14019 39614 14025 39648
rect 1830 35800 1834 35834
rect 1834 35800 1864 35834
rect 1902 35800 1936 35834
rect 1974 35800 2008 35834
rect 2046 35800 2072 35834
rect 2072 35800 2080 35834
rect 1830 35727 1834 35761
rect 1834 35727 1864 35761
rect 1902 35727 1936 35761
rect 1974 35727 2008 35761
rect 2046 35727 2072 35761
rect 2072 35727 2080 35761
rect 1830 35654 1834 35688
rect 1834 35654 1864 35688
rect 1902 35654 1936 35688
rect 1974 35654 2008 35688
rect 2046 35654 2072 35688
rect 2072 35654 2080 35688
rect 1830 35581 1834 35615
rect 1834 35581 1864 35615
rect 1902 35581 1936 35615
rect 1974 35581 2008 35615
rect 2046 35581 2072 35615
rect 2072 35581 2080 35615
rect 1830 35508 1834 35542
rect 1834 35508 1864 35542
rect 1902 35508 1936 35542
rect 1974 35508 2008 35542
rect 2046 35508 2072 35542
rect 2072 35508 2080 35542
rect 1830 35435 1834 35469
rect 1834 35435 1864 35469
rect 1902 35435 1936 35469
rect 1974 35435 2008 35469
rect 2046 35435 2072 35469
rect 2072 35435 2080 35469
rect 1830 35362 1834 35396
rect 1834 35362 1864 35396
rect 1902 35362 1936 35396
rect 1974 35362 2008 35396
rect 2046 35362 2072 35396
rect 2072 35362 2080 35396
rect 1830 35289 1834 35323
rect 1834 35289 1864 35323
rect 1902 35289 1936 35323
rect 1974 35289 2008 35323
rect 2046 35289 2072 35323
rect 2072 35289 2080 35323
rect 1830 35216 1834 35250
rect 1834 35216 1864 35250
rect 1902 35216 1936 35250
rect 1974 35216 2008 35250
rect 2046 35216 2072 35250
rect 2072 35216 2080 35250
rect 1830 35143 1834 35177
rect 1834 35143 1864 35177
rect 1902 35143 1936 35177
rect 1974 35143 2008 35177
rect 2046 35143 2072 35177
rect 2072 35143 2080 35177
rect 1830 35070 1834 35104
rect 1834 35070 1864 35104
rect 1902 35070 1936 35104
rect 1974 35070 2008 35104
rect 2046 35070 2072 35104
rect 2072 35070 2080 35104
rect 1830 34997 1834 35031
rect 1834 34997 1864 35031
rect 1902 34997 1936 35031
rect 1974 34997 2008 35031
rect 2046 34997 2072 35031
rect 2072 34997 2080 35031
rect 1830 34924 1834 34958
rect 1834 34924 1864 34958
rect 1902 34924 1936 34958
rect 1974 34924 2008 34958
rect 2046 34924 2072 34958
rect 2072 34924 2080 34958
rect 1830 34851 1834 34885
rect 1834 34851 1864 34885
rect 1902 34851 1936 34885
rect 1974 34851 2008 34885
rect 2046 34851 2072 34885
rect 2072 34851 2080 34885
rect 1830 34778 1834 34812
rect 1834 34778 1864 34812
rect 1902 34778 1936 34812
rect 1974 34778 2008 34812
rect 2046 34778 2072 34812
rect 2072 34778 2080 34812
rect 1830 34705 1834 34739
rect 1834 34705 1864 34739
rect 1902 34705 1936 34739
rect 1974 34705 2008 34739
rect 2046 34705 2072 34739
rect 2072 34705 2080 34739
rect 1830 34632 1834 34666
rect 1834 34632 1864 34666
rect 1902 34632 1936 34666
rect 1974 34632 2008 34666
rect 2046 34632 2072 34666
rect 2072 34632 2080 34666
rect 1830 34559 1834 34593
rect 1834 34559 1864 34593
rect 1902 34559 1936 34593
rect 1974 34559 2008 34593
rect 2046 34559 2072 34593
rect 2072 34559 2080 34593
rect 1830 34486 1834 34520
rect 1834 34486 1864 34520
rect 1902 34486 1936 34520
rect 1974 34486 2008 34520
rect 2046 34486 2072 34520
rect 2072 34486 2080 34520
rect 1830 34413 1834 34447
rect 1834 34413 1864 34447
rect 1902 34413 1936 34447
rect 1974 34413 2008 34447
rect 2046 34413 2072 34447
rect 2072 34413 2080 34447
rect 1830 34340 1834 34374
rect 1834 34340 1864 34374
rect 1902 34340 1936 34374
rect 1974 34340 2008 34374
rect 2046 34340 2072 34374
rect 2072 34340 2080 34374
rect 1830 34267 1834 34301
rect 1834 34267 1864 34301
rect 1902 34267 1936 34301
rect 1974 34267 2008 34301
rect 2046 34267 2072 34301
rect 2072 34267 2080 34301
rect 1830 34194 1834 34228
rect 1834 34194 1864 34228
rect 1902 34194 1936 34228
rect 1974 34194 2008 34228
rect 2046 34194 2072 34228
rect 2072 34194 2080 34228
rect 2292 39542 2326 39545
rect 2365 39542 13559 39545
rect 2292 39511 2306 39542
rect 2306 39511 2326 39542
rect 2220 37855 2225 39473
rect 2225 39401 2326 39473
rect 2365 39440 2374 39542
rect 2374 39440 13559 39542
rect 13597 39458 13631 39473
rect 2365 39439 2442 39440
rect 2442 39439 13492 39440
rect 13492 39439 13559 39440
rect 13597 39439 13628 39458
rect 13628 39439 13631 39458
rect 2225 37855 2395 39401
rect 2395 37855 2398 39401
rect 2437 39372 2442 39439
rect 2442 39372 13487 39439
rect 13525 39390 13559 39400
rect 13597 39390 13631 39400
rect 2437 39367 13487 39372
rect 13525 39366 13526 39390
rect 13526 39366 13559 39390
rect 13597 39366 13628 39390
rect 13628 39366 13631 39390
rect 13453 39322 13487 39328
rect 13525 39322 13526 39327
rect 13526 39322 13559 39327
rect 13453 39294 13458 39322
rect 13458 39294 13487 39322
rect 13525 39293 13559 39322
rect 13597 39293 13628 39327
rect 13628 39293 13631 39327
rect 13453 39221 13458 39255
rect 13458 39221 13487 39255
rect 13525 39220 13559 39254
rect 13597 39220 13628 39254
rect 13628 39220 13631 39254
rect 13453 39148 13458 39182
rect 13458 39148 13487 39182
rect 13525 39147 13559 39181
rect 13597 39147 13628 39181
rect 13628 39147 13631 39181
rect 3176 39074 3210 39108
rect 3248 39074 3278 39108
rect 3278 39074 3282 39108
rect 3578 39074 3612 39108
rect 3650 39074 3680 39108
rect 3680 39074 3684 39108
rect 4096 39074 4130 39108
rect 4168 39074 4198 39108
rect 4198 39074 4202 39108
rect 4498 39074 4532 39108
rect 4570 39074 4600 39108
rect 4600 39074 4604 39108
rect 5016 39074 5050 39108
rect 5088 39074 5118 39108
rect 5118 39074 5122 39108
rect 5418 39074 5452 39108
rect 5490 39074 5520 39108
rect 5520 39074 5524 39108
rect 5936 39074 5970 39108
rect 6008 39074 6038 39108
rect 6038 39074 6042 39108
rect 6338 39074 6372 39108
rect 6410 39074 6440 39108
rect 6440 39074 6444 39108
rect 6856 39074 6890 39108
rect 6928 39074 6958 39108
rect 6958 39074 6962 39108
rect 7258 39074 7292 39108
rect 7330 39074 7360 39108
rect 7360 39074 7364 39108
rect 7776 39074 7810 39108
rect 7848 39074 7878 39108
rect 7878 39074 7882 39108
rect 8178 39074 8212 39108
rect 8250 39074 8280 39108
rect 8280 39074 8284 39108
rect 8696 39074 8730 39108
rect 8768 39074 8798 39108
rect 8798 39074 8802 39108
rect 9098 39074 9132 39108
rect 9170 39074 9200 39108
rect 9200 39074 9204 39108
rect 9616 39074 9650 39108
rect 9688 39074 9718 39108
rect 9718 39074 9722 39108
rect 10018 39074 10052 39108
rect 10090 39074 10120 39108
rect 10120 39074 10124 39108
rect 10536 39074 10570 39108
rect 10608 39074 10638 39108
rect 10638 39074 10642 39108
rect 10938 39074 10972 39108
rect 11010 39074 11040 39108
rect 11040 39074 11044 39108
rect 11456 39074 11490 39108
rect 11528 39074 11558 39108
rect 11558 39074 11562 39108
rect 11858 39074 11892 39108
rect 11930 39074 11960 39108
rect 11960 39074 11964 39108
rect 12376 39074 12410 39108
rect 12448 39074 12478 39108
rect 12478 39074 12482 39108
rect 12778 39074 12812 39108
rect 12850 39074 12880 39108
rect 12880 39074 12884 39108
rect 13453 39075 13458 39109
rect 13458 39075 13487 39109
rect 2220 37782 2225 37816
rect 2225 37782 2254 37816
rect 2292 37782 2326 37816
rect 2364 37782 2395 37816
rect 2395 37782 2398 37816
rect 2220 37709 2225 37743
rect 2225 37709 2254 37743
rect 2292 37709 2326 37743
rect 2364 37709 2395 37743
rect 2395 37709 2398 37743
rect 2220 37636 2225 37670
rect 2225 37636 2254 37670
rect 2292 37636 2326 37670
rect 2364 37636 2395 37670
rect 2395 37636 2398 37670
rect 2220 37563 2225 37597
rect 2225 37563 2254 37597
rect 2292 37563 2326 37597
rect 2364 37563 2395 37597
rect 2395 37563 2398 37597
rect 2220 37490 2225 37524
rect 2225 37490 2254 37524
rect 2292 37490 2326 37524
rect 2364 37490 2395 37524
rect 2395 37490 2398 37524
rect 2220 37417 2225 37451
rect 2225 37417 2254 37451
rect 2292 37417 2326 37451
rect 2364 37417 2395 37451
rect 2395 37417 2398 37451
rect 2220 37344 2225 37378
rect 2225 37344 2254 37378
rect 2292 37344 2326 37378
rect 2364 37344 2395 37378
rect 2395 37344 2398 37378
rect 2220 37271 2225 37305
rect 2225 37271 2254 37305
rect 2292 37271 2326 37305
rect 2364 37271 2395 37305
rect 2395 37271 2398 37305
rect 2220 37198 2225 37232
rect 2225 37198 2254 37232
rect 2292 37198 2326 37232
rect 2364 37198 2395 37232
rect 2395 37198 2398 37232
rect 2220 37125 2225 37159
rect 2225 37125 2254 37159
rect 2292 37125 2326 37159
rect 2364 37125 2395 37159
rect 2395 37125 2398 37159
rect 2220 37052 2225 37086
rect 2225 37052 2254 37086
rect 2292 37052 2326 37086
rect 2364 37052 2395 37086
rect 2395 37052 2398 37086
rect 13525 39074 13559 39108
rect 13597 39074 13628 39108
rect 13628 39074 13631 39108
rect 2877 37541 3055 39015
rect 2877 37468 2911 37502
rect 2949 37468 2983 37502
rect 3021 37468 3055 37502
rect 2877 37395 2911 37429
rect 2949 37395 2983 37429
rect 3021 37395 3055 37429
rect 2877 37322 2911 37356
rect 2949 37322 2983 37356
rect 3021 37322 3055 37356
rect 2877 37249 2911 37283
rect 2949 37249 2983 37283
rect 3021 37249 3055 37283
rect 2877 37176 2911 37210
rect 2949 37176 2983 37210
rect 3021 37176 3055 37210
rect 2877 37103 2911 37137
rect 2949 37103 2983 37137
rect 3021 37103 3055 37137
rect 3797 37541 3975 39015
rect 3797 37468 3831 37502
rect 3869 37468 3903 37502
rect 3941 37468 3975 37502
rect 3797 37395 3831 37429
rect 3869 37395 3903 37429
rect 3941 37395 3975 37429
rect 3797 37322 3831 37356
rect 3869 37322 3903 37356
rect 3941 37322 3975 37356
rect 3797 37249 3831 37283
rect 3869 37249 3903 37283
rect 3941 37249 3975 37283
rect 3797 37176 3831 37210
rect 3869 37176 3903 37210
rect 3941 37176 3975 37210
rect 3797 37103 3831 37137
rect 3869 37103 3903 37137
rect 3941 37103 3975 37137
rect 4717 38972 4751 39006
rect 4789 38972 4823 39006
rect 4861 38972 4895 39006
rect 4717 38898 4751 38932
rect 4789 38898 4823 38932
rect 4861 38898 4895 38932
rect 4717 38824 4751 38858
rect 4789 38824 4823 38858
rect 4861 38824 4895 38858
rect 4717 38750 4751 38784
rect 4789 38750 4823 38784
rect 4861 38750 4895 38784
rect 4717 38676 4751 38710
rect 4789 38676 4823 38710
rect 4861 38676 4895 38710
rect 4717 38602 4751 38636
rect 4789 38602 4823 38636
rect 4861 38602 4895 38636
rect 4717 38528 4751 38562
rect 4789 38528 4823 38562
rect 4861 38528 4895 38562
rect 4717 38453 4751 38487
rect 4789 38453 4823 38487
rect 4861 38453 4895 38487
rect 4717 38378 4751 38412
rect 4789 38378 4823 38412
rect 4861 38378 4895 38412
rect 4717 38303 4751 38337
rect 4789 38303 4823 38337
rect 4861 38303 4895 38337
rect 4717 38228 4751 38262
rect 4789 38228 4823 38262
rect 4861 38228 4895 38262
rect 4717 38153 4751 38187
rect 4789 38153 4823 38187
rect 4861 38153 4895 38187
rect 4717 38078 4751 38112
rect 4789 38078 4823 38112
rect 4861 38078 4895 38112
rect 4717 38003 4751 38037
rect 4789 38003 4823 38037
rect 4861 38003 4895 38037
rect 4717 37928 4751 37962
rect 4789 37928 4823 37962
rect 4861 37928 4895 37962
rect 4717 37853 4751 37887
rect 4789 37853 4823 37887
rect 4861 37853 4895 37887
rect 4717 37778 4751 37812
rect 4789 37778 4823 37812
rect 4861 37778 4895 37812
rect 4717 37703 4751 37737
rect 4789 37703 4823 37737
rect 4861 37703 4895 37737
rect 4717 37628 4751 37662
rect 4789 37628 4823 37662
rect 4861 37628 4895 37662
rect 4717 37553 4751 37587
rect 4789 37553 4823 37587
rect 4861 37553 4895 37587
rect 4717 37478 4751 37512
rect 4789 37478 4823 37512
rect 4861 37478 4895 37512
rect 4717 37403 4751 37437
rect 4789 37403 4823 37437
rect 4861 37403 4895 37437
rect 4717 37328 4751 37362
rect 4789 37328 4823 37362
rect 4861 37328 4895 37362
rect 4717 37253 4751 37287
rect 4789 37253 4823 37287
rect 4861 37253 4895 37287
rect 4717 37178 4751 37212
rect 4789 37178 4823 37212
rect 4861 37178 4895 37212
rect 4717 37103 4751 37137
rect 4789 37103 4823 37137
rect 4861 37103 4895 37137
rect 5637 38972 5671 39006
rect 5709 38972 5743 39006
rect 5781 38972 5815 39006
rect 5637 38898 5671 38932
rect 5709 38898 5743 38932
rect 5781 38898 5815 38932
rect 5637 38824 5671 38858
rect 5709 38824 5743 38858
rect 5781 38824 5815 38858
rect 5637 38750 5671 38784
rect 5709 38750 5743 38784
rect 5781 38750 5815 38784
rect 5637 38676 5671 38710
rect 5709 38676 5743 38710
rect 5781 38676 5815 38710
rect 5637 38602 5671 38636
rect 5709 38602 5743 38636
rect 5781 38602 5815 38636
rect 5637 38528 5671 38562
rect 5709 38528 5743 38562
rect 5781 38528 5815 38562
rect 5637 38453 5671 38487
rect 5709 38453 5743 38487
rect 5781 38453 5815 38487
rect 5637 38378 5671 38412
rect 5709 38378 5743 38412
rect 5781 38378 5815 38412
rect 5637 38303 5671 38337
rect 5709 38303 5743 38337
rect 5781 38303 5815 38337
rect 5637 38228 5671 38262
rect 5709 38228 5743 38262
rect 5781 38228 5815 38262
rect 5637 38153 5671 38187
rect 5709 38153 5743 38187
rect 5781 38153 5815 38187
rect 5637 38078 5671 38112
rect 5709 38078 5743 38112
rect 5781 38078 5815 38112
rect 5637 38003 5671 38037
rect 5709 38003 5743 38037
rect 5781 38003 5815 38037
rect 5637 37928 5671 37962
rect 5709 37928 5743 37962
rect 5781 37928 5815 37962
rect 5637 37853 5671 37887
rect 5709 37853 5743 37887
rect 5781 37853 5815 37887
rect 5637 37778 5671 37812
rect 5709 37778 5743 37812
rect 5781 37778 5815 37812
rect 5637 37703 5671 37737
rect 5709 37703 5743 37737
rect 5781 37703 5815 37737
rect 5637 37628 5671 37662
rect 5709 37628 5743 37662
rect 5781 37628 5815 37662
rect 5637 37553 5671 37587
rect 5709 37553 5743 37587
rect 5781 37553 5815 37587
rect 5637 37478 5671 37512
rect 5709 37478 5743 37512
rect 5781 37478 5815 37512
rect 5637 37403 5671 37437
rect 5709 37403 5743 37437
rect 5781 37403 5815 37437
rect 5637 37328 5671 37362
rect 5709 37328 5743 37362
rect 5781 37328 5815 37362
rect 5637 37253 5671 37287
rect 5709 37253 5743 37287
rect 5781 37253 5815 37287
rect 5637 37178 5671 37212
rect 5709 37178 5743 37212
rect 5781 37178 5815 37212
rect 5637 37103 5671 37137
rect 5709 37103 5743 37137
rect 5781 37103 5815 37137
rect 6557 38972 6591 39006
rect 6629 38972 6663 39006
rect 6701 38972 6735 39006
rect 6557 38898 6591 38932
rect 6629 38898 6663 38932
rect 6701 38898 6735 38932
rect 6557 38824 6591 38858
rect 6629 38824 6663 38858
rect 6701 38824 6735 38858
rect 6557 38750 6591 38784
rect 6629 38750 6663 38784
rect 6701 38750 6735 38784
rect 6557 38676 6591 38710
rect 6629 38676 6663 38710
rect 6701 38676 6735 38710
rect 6557 38602 6591 38636
rect 6629 38602 6663 38636
rect 6701 38602 6735 38636
rect 6557 38528 6591 38562
rect 6629 38528 6663 38562
rect 6701 38528 6735 38562
rect 6557 38453 6591 38487
rect 6629 38453 6663 38487
rect 6701 38453 6735 38487
rect 6557 38378 6591 38412
rect 6629 38378 6663 38412
rect 6701 38378 6735 38412
rect 6557 38303 6591 38337
rect 6629 38303 6663 38337
rect 6701 38303 6735 38337
rect 6557 38228 6591 38262
rect 6629 38228 6663 38262
rect 6701 38228 6735 38262
rect 6557 38153 6591 38187
rect 6629 38153 6663 38187
rect 6701 38153 6735 38187
rect 6557 38078 6591 38112
rect 6629 38078 6663 38112
rect 6701 38078 6735 38112
rect 6557 38003 6591 38037
rect 6629 38003 6663 38037
rect 6701 38003 6735 38037
rect 6557 37928 6591 37962
rect 6629 37928 6663 37962
rect 6701 37928 6735 37962
rect 6557 37853 6591 37887
rect 6629 37853 6663 37887
rect 6701 37853 6735 37887
rect 6557 37778 6591 37812
rect 6629 37778 6663 37812
rect 6701 37778 6735 37812
rect 6557 37703 6591 37737
rect 6629 37703 6663 37737
rect 6701 37703 6735 37737
rect 6557 37628 6591 37662
rect 6629 37628 6663 37662
rect 6701 37628 6735 37662
rect 6557 37553 6591 37587
rect 6629 37553 6663 37587
rect 6701 37553 6735 37587
rect 6557 37478 6591 37512
rect 6629 37478 6663 37512
rect 6701 37478 6735 37512
rect 6557 37403 6591 37437
rect 6629 37403 6663 37437
rect 6701 37403 6735 37437
rect 6557 37328 6591 37362
rect 6629 37328 6663 37362
rect 6701 37328 6735 37362
rect 6557 37253 6591 37287
rect 6629 37253 6663 37287
rect 6701 37253 6735 37287
rect 6557 37178 6591 37212
rect 6629 37178 6663 37212
rect 6701 37178 6735 37212
rect 6557 37103 6591 37137
rect 6629 37103 6663 37137
rect 6701 37103 6735 37137
rect 7477 38972 7511 39006
rect 7549 38972 7583 39006
rect 7621 38972 7655 39006
rect 7477 38898 7511 38932
rect 7549 38898 7583 38932
rect 7621 38898 7655 38932
rect 7477 38824 7511 38858
rect 7549 38824 7583 38858
rect 7621 38824 7655 38858
rect 7477 38750 7511 38784
rect 7549 38750 7583 38784
rect 7621 38750 7655 38784
rect 7477 38676 7511 38710
rect 7549 38676 7583 38710
rect 7621 38676 7655 38710
rect 7477 38602 7511 38636
rect 7549 38602 7583 38636
rect 7621 38602 7655 38636
rect 7477 38528 7511 38562
rect 7549 38528 7583 38562
rect 7621 38528 7655 38562
rect 7477 38453 7511 38487
rect 7549 38453 7583 38487
rect 7621 38453 7655 38487
rect 7477 38378 7511 38412
rect 7549 38378 7583 38412
rect 7621 38378 7655 38412
rect 7477 38303 7511 38337
rect 7549 38303 7583 38337
rect 7621 38303 7655 38337
rect 7477 38228 7511 38262
rect 7549 38228 7583 38262
rect 7621 38228 7655 38262
rect 7477 38153 7511 38187
rect 7549 38153 7583 38187
rect 7621 38153 7655 38187
rect 7477 38078 7511 38112
rect 7549 38078 7583 38112
rect 7621 38078 7655 38112
rect 7477 38003 7511 38037
rect 7549 38003 7583 38037
rect 7621 38003 7655 38037
rect 7477 37928 7511 37962
rect 7549 37928 7583 37962
rect 7621 37928 7655 37962
rect 7477 37853 7511 37887
rect 7549 37853 7583 37887
rect 7621 37853 7655 37887
rect 7477 37778 7511 37812
rect 7549 37778 7583 37812
rect 7621 37778 7655 37812
rect 7477 37703 7511 37737
rect 7549 37703 7583 37737
rect 7621 37703 7655 37737
rect 7477 37628 7511 37662
rect 7549 37628 7583 37662
rect 7621 37628 7655 37662
rect 7477 37553 7511 37587
rect 7549 37553 7583 37587
rect 7621 37553 7655 37587
rect 7477 37478 7511 37512
rect 7549 37478 7583 37512
rect 7621 37478 7655 37512
rect 7477 37403 7511 37437
rect 7549 37403 7583 37437
rect 7621 37403 7655 37437
rect 7477 37328 7511 37362
rect 7549 37328 7583 37362
rect 7621 37328 7655 37362
rect 7477 37253 7511 37287
rect 7549 37253 7583 37287
rect 7621 37253 7655 37287
rect 7477 37178 7511 37212
rect 7549 37178 7583 37212
rect 7621 37178 7655 37212
rect 7477 37103 7511 37137
rect 7549 37103 7583 37137
rect 7621 37103 7655 37137
rect 8397 38972 8431 39006
rect 8469 38972 8503 39006
rect 8541 38972 8575 39006
rect 8397 38898 8431 38932
rect 8469 38898 8503 38932
rect 8541 38898 8575 38932
rect 8397 38824 8431 38858
rect 8469 38824 8503 38858
rect 8541 38824 8575 38858
rect 8397 38750 8431 38784
rect 8469 38750 8503 38784
rect 8541 38750 8575 38784
rect 8397 38676 8431 38710
rect 8469 38676 8503 38710
rect 8541 38676 8575 38710
rect 8397 38602 8431 38636
rect 8469 38602 8503 38636
rect 8541 38602 8575 38636
rect 8397 38528 8431 38562
rect 8469 38528 8503 38562
rect 8541 38528 8575 38562
rect 8397 38453 8431 38487
rect 8469 38453 8503 38487
rect 8541 38453 8575 38487
rect 8397 38378 8431 38412
rect 8469 38378 8503 38412
rect 8541 38378 8575 38412
rect 8397 38303 8431 38337
rect 8469 38303 8503 38337
rect 8541 38303 8575 38337
rect 8397 38228 8431 38262
rect 8469 38228 8503 38262
rect 8541 38228 8575 38262
rect 8397 38153 8431 38187
rect 8469 38153 8503 38187
rect 8541 38153 8575 38187
rect 8397 38078 8431 38112
rect 8469 38078 8503 38112
rect 8541 38078 8575 38112
rect 8397 38003 8431 38037
rect 8469 38003 8503 38037
rect 8541 38003 8575 38037
rect 8397 37928 8431 37962
rect 8469 37928 8503 37962
rect 8541 37928 8575 37962
rect 8397 37853 8431 37887
rect 8469 37853 8503 37887
rect 8541 37853 8575 37887
rect 8397 37778 8431 37812
rect 8469 37778 8503 37812
rect 8541 37778 8575 37812
rect 8397 37703 8431 37737
rect 8469 37703 8503 37737
rect 8541 37703 8575 37737
rect 8397 37628 8431 37662
rect 8469 37628 8503 37662
rect 8541 37628 8575 37662
rect 8397 37553 8431 37587
rect 8469 37553 8503 37587
rect 8541 37553 8575 37587
rect 8397 37478 8431 37512
rect 8469 37478 8503 37512
rect 8541 37478 8575 37512
rect 8397 37403 8431 37437
rect 8469 37403 8503 37437
rect 8541 37403 8575 37437
rect 8397 37328 8431 37362
rect 8469 37328 8503 37362
rect 8541 37328 8575 37362
rect 8397 37253 8431 37287
rect 8469 37253 8503 37287
rect 8541 37253 8575 37287
rect 8397 37178 8431 37212
rect 8469 37178 8503 37212
rect 8541 37178 8575 37212
rect 8397 37103 8431 37137
rect 8469 37103 8503 37137
rect 8541 37103 8575 37137
rect 9317 38972 9351 39006
rect 9389 38972 9423 39006
rect 9461 38972 9495 39006
rect 9317 38898 9351 38932
rect 9389 38898 9423 38932
rect 9461 38898 9495 38932
rect 9317 38824 9351 38858
rect 9389 38824 9423 38858
rect 9461 38824 9495 38858
rect 9317 38750 9351 38784
rect 9389 38750 9423 38784
rect 9461 38750 9495 38784
rect 9317 38676 9351 38710
rect 9389 38676 9423 38710
rect 9461 38676 9495 38710
rect 9317 38602 9351 38636
rect 9389 38602 9423 38636
rect 9461 38602 9495 38636
rect 9317 38528 9351 38562
rect 9389 38528 9423 38562
rect 9461 38528 9495 38562
rect 9317 38453 9351 38487
rect 9389 38453 9423 38487
rect 9461 38453 9495 38487
rect 9317 38378 9351 38412
rect 9389 38378 9423 38412
rect 9461 38378 9495 38412
rect 9317 38303 9351 38337
rect 9389 38303 9423 38337
rect 9461 38303 9495 38337
rect 9317 38228 9351 38262
rect 9389 38228 9423 38262
rect 9461 38228 9495 38262
rect 9317 38153 9351 38187
rect 9389 38153 9423 38187
rect 9461 38153 9495 38187
rect 9317 38078 9351 38112
rect 9389 38078 9423 38112
rect 9461 38078 9495 38112
rect 9317 38003 9351 38037
rect 9389 38003 9423 38037
rect 9461 38003 9495 38037
rect 9317 37928 9351 37962
rect 9389 37928 9423 37962
rect 9461 37928 9495 37962
rect 9317 37853 9351 37887
rect 9389 37853 9423 37887
rect 9461 37853 9495 37887
rect 9317 37778 9351 37812
rect 9389 37778 9423 37812
rect 9461 37778 9495 37812
rect 9317 37703 9351 37737
rect 9389 37703 9423 37737
rect 9461 37703 9495 37737
rect 9317 37628 9351 37662
rect 9389 37628 9423 37662
rect 9461 37628 9495 37662
rect 9317 37553 9351 37587
rect 9389 37553 9423 37587
rect 9461 37553 9495 37587
rect 9317 37478 9351 37512
rect 9389 37478 9423 37512
rect 9461 37478 9495 37512
rect 9317 37403 9351 37437
rect 9389 37403 9423 37437
rect 9461 37403 9495 37437
rect 9317 37328 9351 37362
rect 9389 37328 9423 37362
rect 9461 37328 9495 37362
rect 9317 37253 9351 37287
rect 9389 37253 9423 37287
rect 9461 37253 9495 37287
rect 9317 37178 9351 37212
rect 9389 37178 9423 37212
rect 9461 37178 9495 37212
rect 9317 37103 9351 37137
rect 9389 37103 9423 37137
rect 9461 37103 9495 37137
rect 10237 38972 10271 39006
rect 10309 38972 10343 39006
rect 10381 38972 10415 39006
rect 10237 38898 10271 38932
rect 10309 38898 10343 38932
rect 10381 38898 10415 38932
rect 10237 38824 10271 38858
rect 10309 38824 10343 38858
rect 10381 38824 10415 38858
rect 10237 38750 10271 38784
rect 10309 38750 10343 38784
rect 10381 38750 10415 38784
rect 10237 38676 10271 38710
rect 10309 38676 10343 38710
rect 10381 38676 10415 38710
rect 10237 38602 10271 38636
rect 10309 38602 10343 38636
rect 10381 38602 10415 38636
rect 10237 38528 10271 38562
rect 10309 38528 10343 38562
rect 10381 38528 10415 38562
rect 10237 38453 10271 38487
rect 10309 38453 10343 38487
rect 10381 38453 10415 38487
rect 10237 38378 10271 38412
rect 10309 38378 10343 38412
rect 10381 38378 10415 38412
rect 10237 38303 10271 38337
rect 10309 38303 10343 38337
rect 10381 38303 10415 38337
rect 10237 38228 10271 38262
rect 10309 38228 10343 38262
rect 10381 38228 10415 38262
rect 10237 38153 10271 38187
rect 10309 38153 10343 38187
rect 10381 38153 10415 38187
rect 10237 38078 10271 38112
rect 10309 38078 10343 38112
rect 10381 38078 10415 38112
rect 10237 38003 10271 38037
rect 10309 38003 10343 38037
rect 10381 38003 10415 38037
rect 10237 37928 10271 37962
rect 10309 37928 10343 37962
rect 10381 37928 10415 37962
rect 10237 37853 10271 37887
rect 10309 37853 10343 37887
rect 10381 37853 10415 37887
rect 10237 37778 10271 37812
rect 10309 37778 10343 37812
rect 10381 37778 10415 37812
rect 10237 37703 10271 37737
rect 10309 37703 10343 37737
rect 10381 37703 10415 37737
rect 10237 37628 10271 37662
rect 10309 37628 10343 37662
rect 10381 37628 10415 37662
rect 10237 37553 10271 37587
rect 10309 37553 10343 37587
rect 10381 37553 10415 37587
rect 10237 37478 10271 37512
rect 10309 37478 10343 37512
rect 10381 37478 10415 37512
rect 10237 37403 10271 37437
rect 10309 37403 10343 37437
rect 10381 37403 10415 37437
rect 10237 37328 10271 37362
rect 10309 37328 10343 37362
rect 10381 37328 10415 37362
rect 10237 37253 10271 37287
rect 10309 37253 10343 37287
rect 10381 37253 10415 37287
rect 10237 37178 10271 37212
rect 10309 37178 10343 37212
rect 10381 37178 10415 37212
rect 10237 37103 10271 37137
rect 10309 37103 10343 37137
rect 10381 37103 10415 37137
rect 11157 38490 11335 39028
rect 11157 38417 11191 38451
rect 11229 38417 11263 38451
rect 11301 38417 11335 38451
rect 11157 38344 11191 38378
rect 11229 38344 11263 38378
rect 11301 38344 11335 38378
rect 11157 38271 11191 38305
rect 11229 38271 11263 38305
rect 11301 38271 11335 38305
rect 11157 38198 11191 38232
rect 11229 38198 11263 38232
rect 11301 38198 11335 38232
rect 11157 38125 11191 38159
rect 11229 38125 11263 38159
rect 11301 38125 11335 38159
rect 11157 38052 11191 38086
rect 11229 38052 11263 38086
rect 11301 38052 11335 38086
rect 11157 37979 11191 38013
rect 11229 37979 11263 38013
rect 11301 37979 11335 38013
rect 11157 37906 11191 37940
rect 11229 37906 11263 37940
rect 11301 37906 11335 37940
rect 11157 37833 11191 37867
rect 11229 37833 11263 37867
rect 11301 37833 11335 37867
rect 11157 37760 11191 37794
rect 11229 37760 11263 37794
rect 11301 37760 11335 37794
rect 11157 37687 11191 37721
rect 11229 37687 11263 37721
rect 11301 37687 11335 37721
rect 11157 37614 11191 37648
rect 11229 37614 11263 37648
rect 11301 37614 11335 37648
rect 11157 37541 11191 37575
rect 11229 37541 11263 37575
rect 11301 37541 11335 37575
rect 11157 37468 11191 37502
rect 11229 37468 11263 37502
rect 11301 37468 11335 37502
rect 11157 37395 11191 37429
rect 11229 37395 11263 37429
rect 11301 37395 11335 37429
rect 11157 37322 11191 37356
rect 11229 37322 11263 37356
rect 11301 37322 11335 37356
rect 11157 37249 11191 37283
rect 11229 37249 11263 37283
rect 11301 37249 11335 37283
rect 11157 37176 11191 37210
rect 11229 37176 11263 37210
rect 11301 37176 11335 37210
rect 11157 37103 11191 37137
rect 11229 37103 11263 37137
rect 11301 37103 11335 37137
rect 12077 38490 12255 39028
rect 12077 38417 12111 38451
rect 12149 38417 12183 38451
rect 12221 38417 12255 38451
rect 12077 38344 12111 38378
rect 12149 38344 12183 38378
rect 12221 38344 12255 38378
rect 12077 38271 12111 38305
rect 12149 38271 12183 38305
rect 12221 38271 12255 38305
rect 12077 38198 12111 38232
rect 12149 38198 12183 38232
rect 12221 38198 12255 38232
rect 12077 38125 12111 38159
rect 12149 38125 12183 38159
rect 12221 38125 12255 38159
rect 12077 38052 12111 38086
rect 12149 38052 12183 38086
rect 12221 38052 12255 38086
rect 12077 37979 12111 38013
rect 12149 37979 12183 38013
rect 12221 37979 12255 38013
rect 12077 37906 12111 37940
rect 12149 37906 12183 37940
rect 12221 37906 12255 37940
rect 12077 37833 12111 37867
rect 12149 37833 12183 37867
rect 12221 37833 12255 37867
rect 12077 37760 12111 37794
rect 12149 37760 12183 37794
rect 12221 37760 12255 37794
rect 12077 37687 12111 37721
rect 12149 37687 12183 37721
rect 12221 37687 12255 37721
rect 12077 37614 12111 37648
rect 12149 37614 12183 37648
rect 12221 37614 12255 37648
rect 12077 37541 12111 37575
rect 12149 37541 12183 37575
rect 12221 37541 12255 37575
rect 12077 37468 12111 37502
rect 12149 37468 12183 37502
rect 12221 37468 12255 37502
rect 12077 37395 12111 37429
rect 12149 37395 12183 37429
rect 12221 37395 12255 37429
rect 12077 37322 12111 37356
rect 12149 37322 12183 37356
rect 12221 37322 12255 37356
rect 12077 37249 12111 37283
rect 12149 37249 12183 37283
rect 12221 37249 12255 37283
rect 12077 37176 12111 37210
rect 12149 37176 12183 37210
rect 12221 37176 12255 37210
rect 12077 37103 12111 37137
rect 12149 37103 12183 37137
rect 12221 37103 12255 37137
rect 12997 38490 13175 39028
rect 12997 38417 13031 38451
rect 13069 38417 13103 38451
rect 13141 38417 13175 38451
rect 12997 38344 13031 38378
rect 13069 38344 13103 38378
rect 13141 38344 13175 38378
rect 12997 38271 13031 38305
rect 13069 38271 13103 38305
rect 13141 38271 13175 38305
rect 12997 38198 13031 38232
rect 13069 38198 13103 38232
rect 13141 38198 13175 38232
rect 12997 38125 13031 38159
rect 13069 38125 13103 38159
rect 13141 38125 13175 38159
rect 12997 38052 13031 38086
rect 13069 38052 13103 38086
rect 13141 38052 13175 38086
rect 12997 37979 13031 38013
rect 13069 37979 13103 38013
rect 13141 37979 13175 38013
rect 12997 37906 13031 37940
rect 13069 37906 13103 37940
rect 13141 37906 13175 37940
rect 12997 37833 13031 37867
rect 13069 37833 13103 37867
rect 13141 37833 13175 37867
rect 12997 37760 13031 37794
rect 13069 37760 13103 37794
rect 13141 37760 13175 37794
rect 12997 37687 13031 37721
rect 13069 37687 13103 37721
rect 13141 37687 13175 37721
rect 12997 37614 13031 37648
rect 13069 37614 13103 37648
rect 13141 37614 13175 37648
rect 12997 37541 13031 37575
rect 13069 37541 13103 37575
rect 13141 37541 13175 37575
rect 12997 37468 13031 37502
rect 13069 37468 13103 37502
rect 13141 37468 13175 37502
rect 12997 37395 13031 37429
rect 13069 37395 13103 37429
rect 13141 37395 13175 37429
rect 12997 37322 13031 37356
rect 13069 37322 13103 37356
rect 13141 37322 13175 37356
rect 12997 37249 13031 37283
rect 13069 37249 13103 37283
rect 13141 37249 13175 37283
rect 12997 37176 13031 37210
rect 13069 37176 13103 37210
rect 13141 37176 13175 37210
rect 12997 37103 13031 37137
rect 13069 37103 13103 37137
rect 13141 37103 13175 37137
rect 13453 39002 13458 39036
rect 13458 39002 13487 39036
rect 13525 39001 13559 39035
rect 13597 39001 13628 39035
rect 13628 39001 13631 39035
rect 13453 38929 13458 38963
rect 13458 38929 13487 38963
rect 13525 38928 13559 38962
rect 13597 38928 13628 38962
rect 13628 38928 13631 38962
rect 13453 38856 13458 38890
rect 13458 38856 13487 38890
rect 13525 38855 13559 38889
rect 13597 38855 13628 38889
rect 13628 38855 13631 38889
rect 13453 38783 13458 38817
rect 13458 38783 13487 38817
rect 13525 38782 13559 38816
rect 13597 38782 13628 38816
rect 13628 38782 13631 38816
rect 13453 38710 13458 38744
rect 13458 38710 13487 38744
rect 13525 38709 13559 38743
rect 13597 38709 13628 38743
rect 13628 38709 13631 38743
rect 13453 38637 13458 38671
rect 13458 38637 13487 38671
rect 13525 38636 13559 38670
rect 13597 38636 13628 38670
rect 13628 38636 13631 38670
rect 13453 38564 13458 38598
rect 13458 38564 13487 38598
rect 13525 38563 13559 38597
rect 13597 38563 13628 38597
rect 13628 38563 13631 38597
rect 13453 38491 13458 38525
rect 13458 38491 13487 38525
rect 13525 38490 13559 38524
rect 13597 38490 13628 38524
rect 13628 38490 13631 38524
rect 13453 38418 13458 38452
rect 13458 38418 13487 38452
rect 13525 38417 13559 38451
rect 13597 38417 13628 38451
rect 13628 38417 13631 38451
rect 13453 38345 13458 38379
rect 13458 38345 13487 38379
rect 13525 38344 13559 38378
rect 13597 38344 13628 38378
rect 13628 38344 13631 38378
rect 13453 38272 13458 38306
rect 13458 38272 13487 38306
rect 13525 38271 13559 38305
rect 13597 38271 13628 38305
rect 13628 38271 13631 38305
rect 13453 38199 13458 38233
rect 13458 38199 13487 38233
rect 13525 38198 13559 38232
rect 13597 38198 13628 38232
rect 13628 38198 13631 38232
rect 13453 38126 13458 38160
rect 13458 38126 13487 38160
rect 13525 38125 13559 38159
rect 13597 38125 13628 38159
rect 13628 38125 13631 38159
rect 13453 38053 13458 38087
rect 13458 38053 13487 38087
rect 13525 38052 13559 38086
rect 13597 38052 13628 38086
rect 13628 38052 13631 38086
rect 13453 37980 13458 38014
rect 13458 37980 13487 38014
rect 13525 37979 13559 38013
rect 13597 37979 13628 38013
rect 13628 37979 13631 38013
rect 13453 37907 13458 37941
rect 13458 37907 13487 37941
rect 13525 37906 13559 37940
rect 13597 37906 13628 37940
rect 13628 37906 13631 37940
rect 13453 37834 13458 37868
rect 13458 37834 13487 37868
rect 13525 37833 13559 37867
rect 13597 37833 13628 37867
rect 13628 37833 13631 37867
rect 13453 37761 13458 37795
rect 13458 37761 13487 37795
rect 13525 37760 13559 37794
rect 13597 37760 13628 37794
rect 13628 37760 13631 37794
rect 13453 37688 13458 37722
rect 13458 37688 13487 37722
rect 13525 37687 13559 37721
rect 13597 37687 13628 37721
rect 13628 37687 13631 37721
rect 13453 37615 13458 37649
rect 13458 37615 13487 37649
rect 13525 37614 13559 37648
rect 13597 37614 13628 37648
rect 13628 37614 13631 37648
rect 13453 37542 13458 37576
rect 13458 37542 13487 37576
rect 13525 37541 13559 37575
rect 13597 37541 13628 37575
rect 13628 37541 13631 37575
rect 13453 37469 13458 37503
rect 13458 37469 13487 37503
rect 13525 37468 13559 37502
rect 13597 37468 13628 37502
rect 13628 37468 13631 37502
rect 13453 37396 13458 37430
rect 13458 37396 13487 37430
rect 13525 37395 13559 37429
rect 13597 37395 13628 37429
rect 13628 37395 13631 37429
rect 13453 37323 13458 37357
rect 13458 37323 13487 37357
rect 13525 37322 13559 37356
rect 13597 37322 13628 37356
rect 13628 37322 13631 37356
rect 13453 37250 13458 37284
rect 13458 37250 13487 37284
rect 13525 37249 13559 37283
rect 13597 37249 13628 37283
rect 13628 37249 13631 37283
rect 13453 37177 13458 37211
rect 13458 37177 13487 37211
rect 13525 37176 13559 37210
rect 13597 37176 13628 37210
rect 13628 37176 13631 37210
rect 13453 37104 13458 37138
rect 13458 37104 13487 37138
rect 13525 37103 13559 37137
rect 13597 37103 13628 37137
rect 13628 37103 13631 37137
rect 2220 36979 2225 37013
rect 2225 36979 2254 37013
rect 2292 36979 2326 37013
rect 2364 36979 2395 37013
rect 2395 36979 2398 37013
rect 13453 37031 13458 37065
rect 13458 37031 13487 37065
rect 2220 36906 2225 36940
rect 2225 36906 2254 36940
rect 2292 36906 2326 36940
rect 2364 36906 2395 36940
rect 2395 36906 2398 36940
rect 2220 36833 2225 36867
rect 2225 36833 2254 36867
rect 2292 36833 2326 36867
rect 2364 36833 2395 36867
rect 2395 36833 2398 36867
rect 2220 36760 2225 36794
rect 2225 36760 2254 36794
rect 2292 36760 2326 36794
rect 2364 36760 2395 36794
rect 2395 36760 2398 36794
rect 2220 36687 2225 36721
rect 2225 36687 2254 36721
rect 2292 36687 2326 36721
rect 2364 36687 2395 36721
rect 2395 36687 2398 36721
rect 2220 36614 2225 36648
rect 2225 36614 2254 36648
rect 2292 36614 2326 36648
rect 2364 36614 2395 36648
rect 2395 36614 2398 36648
rect 2220 36541 2225 36575
rect 2225 36541 2254 36575
rect 2292 36541 2326 36575
rect 2364 36541 2395 36575
rect 2395 36541 2398 36575
rect 2583 36952 2617 36986
rect 2583 36867 2617 36901
rect 2583 36782 2617 36816
rect 2583 36697 2617 36731
rect 2583 36612 2617 36646
rect 2583 36526 2617 36560
rect 2220 36468 2225 36502
rect 2225 36468 2254 36502
rect 2292 36468 2326 36502
rect 2364 36468 2395 36502
rect 2395 36468 2398 36502
rect 13525 37030 13559 37064
rect 13597 37030 13628 37064
rect 13628 37030 13631 37064
rect 13453 36958 13458 36992
rect 13458 36958 13487 36992
rect 13525 36957 13559 36991
rect 13597 36957 13628 36991
rect 13628 36957 13631 36991
rect 13453 36885 13458 36919
rect 13458 36885 13487 36919
rect 13525 36884 13559 36918
rect 13597 36884 13628 36918
rect 13628 36884 13631 36918
rect 13453 36812 13458 36846
rect 13458 36812 13487 36846
rect 13525 36811 13559 36845
rect 13597 36811 13628 36845
rect 13628 36811 13631 36845
rect 13453 36739 13458 36773
rect 13458 36739 13487 36773
rect 13525 36738 13559 36772
rect 13597 36738 13628 36772
rect 13628 36738 13631 36772
rect 13453 36666 13458 36700
rect 13458 36666 13487 36700
rect 13525 36665 13559 36699
rect 13597 36665 13628 36699
rect 13628 36665 13631 36699
rect 13453 36593 13458 36627
rect 13458 36593 13487 36627
rect 13525 36592 13559 36626
rect 13597 36592 13628 36626
rect 13628 36592 13631 36626
rect 13453 36520 13458 36554
rect 13458 36520 13487 36554
rect 13525 36519 13559 36553
rect 13597 36519 13628 36553
rect 13628 36519 13631 36553
rect 2220 36395 2225 36429
rect 2225 36395 2254 36429
rect 2292 36395 2326 36429
rect 2364 36395 2395 36429
rect 2395 36395 2398 36429
rect 13453 36447 13458 36481
rect 13458 36447 13487 36481
rect 13525 36446 13559 36480
rect 13597 36446 13628 36480
rect 13628 36446 13631 36480
rect 2220 36322 2225 36356
rect 2225 36322 2254 36356
rect 2292 36322 2326 36356
rect 2364 36322 2395 36356
rect 2395 36322 2398 36356
rect 2220 36249 2225 36283
rect 2225 36249 2254 36283
rect 2292 36249 2326 36283
rect 2364 36249 2395 36283
rect 2395 36249 2398 36283
rect 2220 36176 2225 36210
rect 2225 36176 2254 36210
rect 2292 36176 2326 36210
rect 2364 36176 2395 36210
rect 2395 36176 2398 36210
rect 2220 36103 2225 36137
rect 2225 36103 2254 36137
rect 2292 36103 2326 36137
rect 2364 36103 2395 36137
rect 2395 36103 2398 36137
rect 2220 36030 2225 36064
rect 2225 36030 2254 36064
rect 2292 36030 2326 36064
rect 2364 36030 2395 36064
rect 2395 36030 2398 36064
rect 2220 35957 2225 35991
rect 2225 35957 2254 35991
rect 2292 35957 2326 35991
rect 2364 35957 2395 35991
rect 2395 35957 2398 35991
rect 2220 35884 2225 35918
rect 2225 35884 2254 35918
rect 2292 35884 2326 35918
rect 2364 35884 2395 35918
rect 2395 35884 2398 35918
rect 2220 35811 2225 35845
rect 2225 35811 2254 35845
rect 2292 35811 2326 35845
rect 2364 35811 2395 35845
rect 2395 35811 2398 35845
rect 2220 35738 2225 35772
rect 2225 35738 2254 35772
rect 2292 35738 2326 35772
rect 2364 35738 2395 35772
rect 2395 35738 2398 35772
rect 2220 35665 2225 35699
rect 2225 35665 2254 35699
rect 2292 35665 2326 35699
rect 2364 35665 2395 35699
rect 2395 35665 2398 35699
rect 2220 35592 2225 35626
rect 2225 35592 2254 35626
rect 2292 35592 2326 35626
rect 2364 35592 2395 35626
rect 2395 35592 2398 35626
rect 2220 35519 2225 35553
rect 2225 35519 2254 35553
rect 2292 35519 2326 35553
rect 2364 35519 2395 35553
rect 2395 35519 2398 35553
rect 2220 35446 2225 35480
rect 2225 35446 2254 35480
rect 2292 35446 2326 35480
rect 2364 35446 2395 35480
rect 2395 35446 2398 35480
rect 2220 35373 2225 35407
rect 2225 35373 2254 35407
rect 2292 35373 2326 35407
rect 2364 35373 2395 35407
rect 2395 35373 2398 35407
rect 2220 35300 2225 35334
rect 2225 35300 2254 35334
rect 2292 35300 2326 35334
rect 2364 35300 2395 35334
rect 2395 35300 2398 35334
rect 2220 35227 2225 35261
rect 2225 35227 2254 35261
rect 2292 35227 2326 35261
rect 2364 35227 2395 35261
rect 2395 35227 2398 35261
rect 2220 35154 2225 35188
rect 2225 35154 2254 35188
rect 2292 35154 2326 35188
rect 2364 35154 2395 35188
rect 2395 35154 2398 35188
rect 2220 35081 2225 35115
rect 2225 35081 2254 35115
rect 2292 35081 2326 35115
rect 2364 35081 2395 35115
rect 2395 35081 2398 35115
rect 2220 35008 2225 35042
rect 2225 35008 2254 35042
rect 2292 35008 2326 35042
rect 2364 35008 2395 35042
rect 2395 35008 2398 35042
rect 2220 34935 2225 34969
rect 2225 34935 2254 34969
rect 2292 34935 2326 34969
rect 2364 34935 2395 34969
rect 2395 34935 2398 34969
rect 2220 34862 2225 34896
rect 2225 34862 2254 34896
rect 2292 34862 2326 34896
rect 2364 34862 2395 34896
rect 2395 34862 2398 34896
rect 2220 34789 2225 34823
rect 2225 34789 2254 34823
rect 2292 34789 2326 34823
rect 2364 34789 2395 34823
rect 2395 34789 2398 34823
rect 2220 34716 2225 34750
rect 2225 34716 2254 34750
rect 2292 34716 2326 34750
rect 2364 34716 2395 34750
rect 2395 34716 2398 34750
rect 2220 34643 2225 34677
rect 2225 34643 2254 34677
rect 2292 34643 2326 34677
rect 2364 34643 2395 34677
rect 2395 34643 2398 34677
rect 2220 34570 2225 34604
rect 2225 34570 2254 34604
rect 2292 34570 2326 34604
rect 2364 34570 2395 34604
rect 2395 34570 2398 34604
rect 2220 34497 2225 34531
rect 2225 34497 2254 34531
rect 2292 34497 2326 34531
rect 2364 34497 2395 34531
rect 2395 34497 2398 34531
rect 2220 34424 2225 34458
rect 2225 34424 2254 34458
rect 2292 34424 2326 34458
rect 2364 34424 2395 34458
rect 2395 34424 2398 34458
rect 2220 34351 2225 34385
rect 2225 34351 2254 34385
rect 2292 34351 2326 34385
rect 2364 34351 2395 34385
rect 2395 34351 2398 34385
rect 2220 34278 2225 34312
rect 2225 34278 2254 34312
rect 2292 34278 2326 34312
rect 2364 34278 2395 34312
rect 2395 34278 2398 34312
rect 2220 34205 2225 34239
rect 2225 34205 2254 34239
rect 2292 34205 2326 34239
rect 2364 34205 2395 34239
rect 2395 34205 2398 34239
rect 2943 36328 2977 36362
rect 3021 36328 3055 36362
rect 2943 36256 2977 36290
rect 3021 36256 3055 36290
rect 2943 36184 2977 36218
rect 3021 36184 3055 36218
rect 2943 36112 2977 36146
rect 3021 36112 3055 36146
rect 2943 36040 2977 36074
rect 3021 36040 3055 36074
rect 2943 35968 2977 36002
rect 3021 35968 3055 36002
rect 2943 35896 2977 35930
rect 3021 35896 3055 35930
rect 2943 35824 2977 35858
rect 3021 35824 3055 35858
rect 2943 35752 2977 35786
rect 3021 35752 3055 35786
rect 2943 35680 2977 35714
rect 3021 35680 3055 35714
rect 2943 35608 2977 35642
rect 3021 35608 3055 35642
rect 2943 35536 2977 35570
rect 3021 35536 3055 35570
rect 2943 35464 2977 35498
rect 3021 35464 3055 35498
rect 2943 35392 2977 35426
rect 3021 35392 3055 35426
rect 2943 35320 2977 35354
rect 3021 35320 3055 35354
rect 2943 35248 2977 35282
rect 3021 35248 3055 35282
rect 2943 35176 2977 35210
rect 3021 35176 3055 35210
rect 2943 35104 2977 35138
rect 3021 35104 3055 35138
rect 2943 35032 2977 35066
rect 3021 35032 3055 35066
rect 2943 34960 2977 34994
rect 3021 34960 3055 34994
rect 2943 34888 2977 34922
rect 3021 34888 3055 34922
rect 2943 34816 2977 34850
rect 3021 34816 3055 34850
rect 2943 34744 2977 34778
rect 3021 34744 3055 34778
rect 2943 34672 2977 34706
rect 3021 34672 3055 34706
rect 2943 34600 2977 34634
rect 3021 34600 3055 34634
rect 2943 34528 2977 34562
rect 3021 34528 3055 34562
rect 2943 34456 2977 34490
rect 3021 34456 3055 34490
rect 2943 34384 2977 34418
rect 3021 34384 3055 34418
rect 2943 34312 2977 34346
rect 3021 34312 3055 34346
rect 2943 34240 2977 34274
rect 3021 34240 3055 34274
rect 1702 34110 1736 34144
rect 1808 34110 1834 34144
rect 1834 34110 1842 34144
rect 1702 34035 1736 34069
rect 1808 34035 1834 34069
rect 1834 34035 1842 34069
rect 1702 33960 1736 33994
rect 1808 33960 1834 33994
rect 1834 33960 1842 33994
rect 1702 33885 1736 33919
rect 1808 33885 1834 33919
rect 1834 33885 1842 33919
rect 1702 33810 1736 33844
rect 1808 33810 1834 33844
rect 1834 33810 1842 33844
rect 1702 33735 1736 33769
rect 1808 33735 1834 33769
rect 1834 33735 1842 33769
rect 1702 33660 1736 33694
rect 1808 33660 1834 33694
rect 1834 33660 1842 33694
rect 1702 33585 1736 33619
rect 1808 33585 1834 33619
rect 1834 33585 1842 33619
rect 1702 33510 1736 33544
rect 1808 33510 1834 33544
rect 1834 33510 1842 33544
rect 1702 33435 1736 33469
rect 1808 33435 1834 33469
rect 1834 33435 1842 33469
rect 1702 33360 1736 33394
rect 1808 33360 1834 33394
rect 1834 33360 1842 33394
rect 1702 33285 1736 33319
rect 1808 33285 1834 33319
rect 1834 33285 1842 33319
rect 1702 33210 1736 33244
rect 1808 33210 1834 33244
rect 1834 33210 1842 33244
rect 1702 33135 1736 33169
rect 1808 33135 1834 33169
rect 1834 33135 1842 33169
rect 1702 33060 1736 33094
rect 1808 33060 1834 33094
rect 1834 33060 1842 33094
rect 1702 32985 1736 33019
rect 1808 32985 1834 33019
rect 1834 32985 1842 33019
rect 1702 32910 1736 32944
rect 1808 32910 1834 32944
rect 1834 32910 1842 32944
rect 1702 32835 1736 32869
rect 1808 32835 1834 32869
rect 1834 32835 1842 32869
rect 1702 32759 1736 32793
rect 1808 32759 1834 32793
rect 1834 32759 1842 32793
rect 1702 32683 1736 32717
rect 1808 32683 1834 32717
rect 1834 32683 1842 32717
rect 1702 32607 1736 32641
rect 1808 32607 1834 32641
rect 1834 32607 1842 32641
rect 1702 32531 1736 32565
rect 1808 32531 1834 32565
rect 1834 32531 1842 32565
rect 2154 34069 2188 34103
rect 2226 34069 2260 34103
rect 2154 33996 2188 34030
rect 2226 33996 2260 34030
rect 2154 33923 2188 33957
rect 2226 33923 2260 33957
rect 2154 33850 2188 33884
rect 2226 33850 2260 33884
rect 2154 33777 2188 33811
rect 2226 33777 2260 33811
rect 2154 33704 2188 33738
rect 2226 33704 2260 33738
rect 2154 33631 2188 33665
rect 2226 33631 2260 33665
rect 2154 33558 2188 33592
rect 2226 33558 2260 33592
rect 2154 33485 2188 33519
rect 2226 33485 2260 33519
rect 2154 33412 2188 33446
rect 2226 33412 2260 33446
rect 2154 33339 2188 33373
rect 2226 33339 2260 33373
rect 2154 33266 2188 33300
rect 2226 33266 2260 33300
rect 2154 33193 2188 33227
rect 2226 33193 2260 33227
rect 2154 33120 2188 33154
rect 2226 33120 2260 33154
rect 2154 33047 2188 33081
rect 2226 33047 2260 33081
rect 2154 32974 2188 33008
rect 2226 32974 2260 33008
rect 2154 32901 2188 32935
rect 2226 32901 2260 32935
rect 2154 32827 2188 32861
rect 2226 32827 2260 32861
rect 2154 32753 2188 32787
rect 2226 32753 2260 32787
rect 2154 32679 2188 32713
rect 2226 32679 2260 32713
rect 2154 32605 2188 32639
rect 2226 32605 2260 32639
rect 2154 32531 2188 32565
rect 2226 32531 2260 32565
rect 1840 31749 1874 31783
rect 1946 31749 1980 31783
rect 1840 31677 1874 31711
rect 1946 31677 1980 31711
rect 1840 31604 1874 31638
rect 1946 31605 1980 31639
rect 1840 31531 1874 31565
rect 1946 31533 1980 31567
rect 1840 31458 1874 31492
rect 1946 31461 1980 31495
rect 1840 31385 1874 31419
rect 1946 31389 1980 31423
rect 1840 31312 1874 31346
rect 1946 31317 1980 31351
rect 1840 31239 1874 31273
rect 1946 31245 1980 31279
rect 1840 31166 1874 31200
rect 1946 31173 1980 31207
rect 1840 31093 1874 31127
rect 1946 31101 1980 31135
rect 1840 31020 1874 31054
rect 1946 31029 1980 31063
rect 1840 30947 1874 30981
rect 1946 30957 1980 30991
rect 1840 30874 1874 30908
rect 1946 30885 1980 30919
rect 1840 30801 1874 30835
rect 1946 30813 1980 30847
rect 1840 30728 1874 30762
rect 1946 30741 1980 30775
rect 1840 30655 1874 30689
rect 1946 30669 1980 30703
rect 1840 30582 1874 30616
rect 1946 30597 1980 30631
rect 1840 30509 1874 30543
rect 1946 30525 1980 30559
rect 1840 30436 1874 30470
rect 1946 30453 1980 30487
rect 1840 30363 1874 30397
rect 1946 30381 1980 30415
rect 1840 30290 1874 30324
rect 1946 30309 1980 30343
rect 1840 30217 1874 30251
rect 1946 30237 1980 30271
rect 1840 30144 1874 30178
rect 1946 30165 1980 30199
rect 1840 30071 1874 30105
rect 1946 30093 1980 30127
rect 1840 29998 1874 30032
rect 1946 30021 1980 30055
rect 1840 29925 1874 29959
rect 1946 29949 1980 29983
rect 1840 29852 1874 29886
rect 1946 29877 1980 29911
rect 1840 29779 1874 29813
rect 1946 29805 1980 29839
rect 1840 29706 1874 29740
rect 1946 29733 1980 29767
rect 1840 29633 1874 29667
rect 1946 29661 1980 29695
rect 1840 29560 1874 29594
rect 1946 29589 1980 29623
rect 1840 29487 1874 29521
rect 1946 29517 1980 29551
rect 1840 29414 1874 29448
rect 1946 29445 1980 29479
rect 1840 29341 1874 29375
rect 1946 29373 1980 29407
rect 1840 29268 1874 29302
rect 1946 29301 1980 29335
rect 1946 29229 1980 29263
rect 1840 29195 1874 29229
rect 1946 29156 1980 29190
rect 1840 29122 1874 29156
rect 1946 29083 1980 29117
rect 1840 29049 1874 29083
rect 1946 29010 1980 29044
rect 1840 28976 1874 29010
rect 1946 28937 1980 28971
rect 1840 28903 1874 28937
rect 1946 28864 1980 28898
rect 1840 28830 1874 28864
rect 1946 28791 1980 28825
rect 1840 28757 1874 28791
rect 1946 28718 1980 28752
rect 1840 28684 1874 28718
rect 1946 28645 1980 28679
rect 1840 28611 1874 28645
rect 1946 28572 1980 28606
rect 1840 28538 1874 28572
rect 1946 28499 1980 28533
rect 1840 28465 1874 28499
rect 1946 28426 1980 28460
rect 1840 28392 1874 28426
rect 1946 28353 1980 28387
rect 1840 28319 1874 28353
rect 1946 28280 1980 28314
rect 1840 28246 1874 28280
rect 1946 28207 1980 28241
rect 1840 28173 1874 28207
rect 1946 28134 1980 28168
rect 1840 28100 1874 28134
rect 1946 28061 1980 28095
rect 1840 28027 1874 28061
rect 1946 27988 1980 28022
rect 1840 27954 1874 27988
rect 1946 27915 1980 27949
rect 1840 27881 1874 27915
rect 1946 27842 1980 27876
rect 1840 27808 1874 27842
rect 1946 27769 1980 27803
rect 1840 27735 1874 27769
rect 1946 27696 1980 27730
rect 1840 27662 1874 27696
rect 1946 27623 1980 27657
rect 1840 27589 1874 27623
rect 1946 27550 1980 27584
rect 1840 27516 1874 27550
rect 1946 27477 1980 27511
rect 1840 27443 1874 27477
rect 1946 27404 1980 27438
rect 1840 27370 1874 27404
rect 1946 27331 1980 27365
rect 1840 27297 1874 27331
rect 1946 27258 1980 27292
rect 1840 27224 1874 27258
rect 1946 27185 1980 27219
rect 1840 27151 1874 27185
rect 1946 27112 1980 27146
rect 1840 27078 1874 27112
rect 1946 27039 1980 27073
rect 2943 34168 2977 34202
rect 3021 34168 3055 34202
rect 2943 34096 2977 34130
rect 3021 34096 3055 34130
rect 2943 34024 2977 34058
rect 3021 34024 3055 34058
rect 2943 33952 2977 33986
rect 3021 33952 3055 33986
rect 2943 33880 2977 33914
rect 3021 33880 3055 33914
rect 2943 33808 2977 33842
rect 3021 33808 3055 33842
rect 2943 33736 2977 33770
rect 3021 33736 3055 33770
rect 2943 33664 2977 33698
rect 3021 33664 3055 33698
rect 2943 33592 2977 33626
rect 3021 33592 3055 33626
rect 2943 33520 2977 33554
rect 3021 33520 3055 33554
rect 2943 33448 2977 33482
rect 3021 33448 3055 33482
rect 2943 33376 2977 33410
rect 3021 33376 3055 33410
rect 2943 33304 2977 33338
rect 3021 33304 3055 33338
rect 2943 33232 2977 33266
rect 3021 33232 3055 33266
rect 2943 33160 2977 33194
rect 3021 33160 3055 33194
rect 2943 33087 2977 33121
rect 3021 33087 3055 33121
rect 2943 33014 2977 33048
rect 3021 33014 3055 33048
rect 2943 32941 2977 32975
rect 3021 32941 3055 32975
rect 2943 32868 2977 32902
rect 3021 32868 3055 32902
rect 2943 32795 2977 32829
rect 3021 32795 3055 32829
rect 2943 32722 2977 32756
rect 3021 32722 3055 32756
rect 2943 32649 2977 32683
rect 3021 32649 3055 32683
rect 2943 32576 2977 32610
rect 3021 32576 3055 32610
rect 2943 32503 2977 32537
rect 3021 32503 3055 32537
rect 3797 33160 3975 36362
rect 3797 33087 3831 33121
rect 3869 33087 3903 33121
rect 3941 33087 3975 33121
rect 3797 33014 3831 33048
rect 3869 33014 3903 33048
rect 3941 33014 3975 33048
rect 3797 32941 3831 32975
rect 3869 32941 3903 32975
rect 3941 32941 3975 32975
rect 3797 32868 3831 32902
rect 3869 32868 3903 32902
rect 3941 32868 3975 32902
rect 3797 32795 3831 32829
rect 3869 32795 3903 32829
rect 3941 32795 3975 32829
rect 3797 32722 3831 32756
rect 3869 32722 3903 32756
rect 3941 32722 3975 32756
rect 3797 32649 3831 32683
rect 3869 32649 3903 32683
rect 3941 32649 3975 32683
rect 3797 32576 3831 32610
rect 3869 32576 3903 32610
rect 3941 32576 3975 32610
rect 3797 32503 3831 32537
rect 3869 32503 3903 32537
rect 3941 32503 3975 32537
rect 4717 32503 4895 36353
rect 5637 32503 5815 36353
rect 6557 32503 6735 36353
rect 7477 32503 7655 36353
rect 8397 32503 8575 36353
rect 9317 32503 9495 36353
rect 10237 32503 10415 36353
rect 11157 32503 11335 36353
rect 12077 32503 12255 36353
rect 12997 32503 13175 36353
rect 13453 36374 13458 36408
rect 13458 36374 13487 36408
rect 13525 36373 13559 36407
rect 13597 36373 13628 36407
rect 13628 36373 13631 36407
rect 13453 36301 13458 36335
rect 13458 36301 13487 36335
rect 13525 36300 13559 36334
rect 13597 36300 13628 36334
rect 13628 36300 13631 36334
rect 13453 36228 13458 36262
rect 13458 36228 13487 36262
rect 13525 36227 13559 36261
rect 13597 36227 13628 36261
rect 13628 36227 13631 36261
rect 13453 36155 13458 36189
rect 13458 36155 13487 36189
rect 13525 36154 13559 36188
rect 13597 36154 13628 36188
rect 13628 36154 13631 36188
rect 13453 36082 13458 36116
rect 13458 36082 13487 36116
rect 13525 36081 13559 36115
rect 13597 36081 13628 36115
rect 13628 36081 13631 36115
rect 13453 36009 13458 36043
rect 13458 36009 13487 36043
rect 13525 36008 13559 36042
rect 13597 36008 13628 36042
rect 13628 36008 13631 36042
rect 13453 35936 13458 35970
rect 13458 35936 13487 35970
rect 13525 35935 13559 35969
rect 13597 35935 13628 35969
rect 13628 35935 13631 35969
rect 13453 35863 13458 35897
rect 13458 35863 13487 35897
rect 13525 35824 13628 35896
rect 13453 33198 13458 35824
rect 13458 33198 13628 35824
rect 13628 33198 13631 35896
rect 13775 39543 13781 39577
rect 13781 39543 13809 39577
rect 13847 39542 13881 39576
rect 13919 39541 13953 39575
rect 13991 39541 14019 39575
rect 14019 39541 14025 39575
rect 13775 39470 13781 39504
rect 13781 39470 13809 39504
rect 13847 39469 13881 39503
rect 13919 39468 13953 39502
rect 13991 39468 14019 39502
rect 14019 39468 14025 39502
rect 13775 39397 13781 39431
rect 13781 39397 13809 39431
rect 13847 39396 13881 39430
rect 13919 39395 13953 39429
rect 13991 39395 14019 39429
rect 14019 39395 14025 39429
rect 13775 39324 13781 39358
rect 13781 39324 13809 39358
rect 13847 39323 13881 39357
rect 13919 39322 13953 39356
rect 13991 39322 14019 39356
rect 14019 39322 14025 39356
rect 13775 39251 13781 39285
rect 13781 39251 13809 39285
rect 13847 39250 13881 39284
rect 13919 39249 13953 39283
rect 13991 39249 14019 39283
rect 14019 39249 14025 39283
rect 13775 39178 13781 39212
rect 13781 39178 13809 39212
rect 13847 39177 13881 39211
rect 13919 39176 13953 39210
rect 13991 39176 14019 39210
rect 14019 39176 14025 39210
rect 13775 39105 13781 39139
rect 13781 39105 13809 39139
rect 13847 39104 13881 39138
rect 13919 39103 13953 39137
rect 13991 39103 14019 39137
rect 14019 39103 14025 39137
rect 13775 39032 13781 39066
rect 13781 39032 13809 39066
rect 13847 39031 13881 39065
rect 13919 39030 13953 39064
rect 13991 39030 14019 39064
rect 14019 39030 14025 39064
rect 13775 38959 13781 38993
rect 13781 38959 13809 38993
rect 13847 38958 13881 38992
rect 13919 38957 13953 38991
rect 13991 38957 14019 38991
rect 14019 38957 14025 38991
rect 13775 38886 13781 38920
rect 13781 38886 13809 38920
rect 13847 38885 13881 38919
rect 13919 38884 13953 38918
rect 13991 38884 14019 38918
rect 14019 38884 14025 38918
rect 13775 38813 13781 38847
rect 13781 38813 13809 38847
rect 13847 38812 13881 38846
rect 13919 38811 13953 38845
rect 13991 38811 14019 38845
rect 14019 38811 14025 38845
rect 13775 38740 13781 38774
rect 13781 38740 13809 38774
rect 13847 38739 13881 38773
rect 13919 38738 13953 38772
rect 13991 38738 14019 38772
rect 14019 38738 14025 38772
rect 13775 38667 13781 38701
rect 13781 38667 13809 38701
rect 13847 38666 13881 38700
rect 13919 38665 13953 38699
rect 13991 38665 14019 38699
rect 14019 38665 14025 38699
rect 13775 38594 13781 38628
rect 13781 38594 13809 38628
rect 13847 38593 13881 38627
rect 13919 38592 13953 38626
rect 13991 38592 14019 38626
rect 14019 38592 14025 38626
rect 13775 38521 13781 38555
rect 13781 38521 13809 38555
rect 13847 38520 13881 38554
rect 13919 38519 13953 38553
rect 13991 38519 14019 38553
rect 14019 38519 14025 38553
rect 13775 38448 13781 38482
rect 13781 38448 13809 38482
rect 13847 38447 13881 38481
rect 13919 38446 13953 38480
rect 13991 38446 14019 38480
rect 14019 38446 14025 38480
rect 13775 38375 13781 38409
rect 13781 38375 13809 38409
rect 13847 38374 13881 38408
rect 13919 38373 13953 38407
rect 13991 38373 14019 38407
rect 14019 38373 14025 38407
rect 13775 38302 13781 38336
rect 13781 38302 13809 38336
rect 13847 38301 13881 38335
rect 13919 38300 13953 38334
rect 13991 38300 14019 38334
rect 14019 38300 14025 38334
rect 13775 38229 13781 38263
rect 13781 38229 13809 38263
rect 13847 38228 13881 38262
rect 13919 38227 13953 38261
rect 13991 38227 14019 38261
rect 14019 38227 14025 38261
rect 13775 38156 13781 38190
rect 13781 38156 13809 38190
rect 13847 38155 13881 38189
rect 13919 38154 13953 38188
rect 13991 38154 14019 38188
rect 14019 38154 14025 38188
rect 13775 38083 13781 38117
rect 13781 38083 13809 38117
rect 13847 38082 13881 38116
rect 13919 38081 13953 38115
rect 13991 38081 14019 38115
rect 14019 38081 14025 38115
rect 13775 38010 13781 38044
rect 13781 38010 13809 38044
rect 13847 38009 13881 38043
rect 13919 38008 13953 38042
rect 13991 38008 14019 38042
rect 14019 38008 14025 38042
rect 13775 37937 13781 37971
rect 13781 37937 13809 37971
rect 13847 37936 13881 37970
rect 13919 37935 13953 37969
rect 13991 37935 14019 37969
rect 14019 37935 14025 37969
rect 13775 37864 13781 37898
rect 13781 37864 13809 37898
rect 13847 37863 13881 37897
rect 13919 37862 13953 37896
rect 13991 37862 14019 37896
rect 14019 37862 14025 37896
rect 13775 37791 13781 37825
rect 13781 37791 13809 37825
rect 13847 37790 13881 37824
rect 13919 37789 13953 37823
rect 13991 37789 14019 37823
rect 14019 37789 14025 37823
rect 13775 37718 13781 37752
rect 13781 37718 13809 37752
rect 13847 37717 13881 37751
rect 13919 37716 13953 37750
rect 13991 37716 14019 37750
rect 14019 37716 14025 37750
rect 13775 37645 13781 37679
rect 13781 37645 13809 37679
rect 13847 37644 13881 37678
rect 13919 37643 13953 37677
rect 13991 37643 14019 37677
rect 14019 37643 14025 37677
rect 13775 37572 13781 37606
rect 13781 37572 13809 37606
rect 13847 37571 13881 37605
rect 13919 37570 13953 37604
rect 13991 37570 14019 37604
rect 14019 37570 14025 37604
rect 13775 37499 13781 37533
rect 13781 37499 13809 37533
rect 13847 37498 13881 37532
rect 13919 37497 13953 37531
rect 13991 37497 14019 37531
rect 14019 37497 14025 37531
rect 13775 37426 13781 37460
rect 13781 37426 13809 37460
rect 13847 37425 13881 37459
rect 13919 37424 13953 37458
rect 13991 37424 14019 37458
rect 14019 37424 14025 37458
rect 13775 37353 13781 37387
rect 13781 37353 13809 37387
rect 13847 37352 13881 37386
rect 13919 37351 13953 37385
rect 13991 37351 14019 37385
rect 14019 37351 14025 37385
rect 13775 37280 13781 37314
rect 13781 37280 13809 37314
rect 13847 37279 13881 37313
rect 13919 37278 13953 37312
rect 13991 37278 14019 37312
rect 14019 37278 14025 37312
rect 13775 37207 13781 37241
rect 13781 37207 13809 37241
rect 13847 37206 13881 37240
rect 13919 37205 13953 37239
rect 13991 37205 14019 37239
rect 14019 37205 14025 37239
rect 13775 37134 13781 37168
rect 13781 37134 13809 37168
rect 13847 37133 13881 37167
rect 13919 37132 13953 37166
rect 13991 37132 14019 37166
rect 14019 37132 14025 37166
rect 13775 37061 13781 37095
rect 13781 37061 13809 37095
rect 13847 37060 13881 37094
rect 13919 37059 13953 37093
rect 13991 37059 14019 37093
rect 14019 37059 14025 37093
rect 13775 36988 13781 37022
rect 13781 36988 13809 37022
rect 13847 36987 13881 37021
rect 13919 36986 13953 37020
rect 13991 36986 14019 37020
rect 14019 36986 14025 37020
rect 13775 36915 13781 36949
rect 13781 36915 13809 36949
rect 13847 36914 13881 36948
rect 13919 36913 13953 36947
rect 13991 36913 14019 36947
rect 14019 36913 14025 36947
rect 13775 36842 13781 36876
rect 13781 36842 13809 36876
rect 13847 36841 13881 36875
rect 13919 36840 13953 36874
rect 13991 36840 14019 36874
rect 14019 36840 14025 36874
rect 13775 36769 13781 36803
rect 13781 36769 13809 36803
rect 13847 36768 13881 36802
rect 13919 36767 13953 36801
rect 13991 36767 14019 36801
rect 14019 36767 14025 36801
rect 13775 36696 13781 36730
rect 13781 36696 13809 36730
rect 13847 36695 13881 36729
rect 13919 36694 13953 36728
rect 13991 36694 14019 36728
rect 14019 36694 14025 36728
rect 13775 36623 13781 36657
rect 13781 36623 13809 36657
rect 13847 36622 13881 36656
rect 13919 36621 13953 36655
rect 13991 36621 14019 36655
rect 14019 36621 14025 36655
rect 13775 36550 13781 36584
rect 13781 36550 13809 36584
rect 13847 36549 13881 36583
rect 13919 36548 13953 36582
rect 13991 36548 14019 36582
rect 14019 36548 14025 36582
rect 13775 36477 13781 36511
rect 13781 36477 13809 36511
rect 13847 36476 13881 36510
rect 13919 36475 13953 36509
rect 13991 36475 14019 36509
rect 14019 36475 14025 36509
rect 13775 36404 13781 36438
rect 13781 36404 13809 36438
rect 13847 36403 13881 36437
rect 13919 36402 13953 36436
rect 13991 36402 14019 36436
rect 14019 36402 14025 36436
rect 13775 36331 13781 36365
rect 13781 36331 13809 36365
rect 13847 36330 13881 36364
rect 13919 36329 13953 36363
rect 13991 36329 14019 36363
rect 14019 36329 14025 36363
rect 13775 36258 13781 36292
rect 13781 36258 13809 36292
rect 13847 36257 13881 36291
rect 13919 36256 13953 36290
rect 13991 36256 14019 36290
rect 14019 36256 14025 36290
rect 13775 36185 13781 36219
rect 13781 36185 13809 36219
rect 13847 36184 13881 36218
rect 13919 36183 13953 36217
rect 13991 36183 14019 36217
rect 14019 36183 14025 36217
rect 13775 36112 13781 36146
rect 13781 36112 13809 36146
rect 13847 36111 13881 36145
rect 13919 36110 13953 36144
rect 13991 36110 14019 36144
rect 14019 36110 14025 36144
rect 13775 36039 13781 36073
rect 13781 36039 13809 36073
rect 13847 36038 13881 36072
rect 13919 36037 13953 36071
rect 13991 36037 14019 36071
rect 14019 36037 14025 36071
rect 13775 35966 13781 36000
rect 13781 35966 13809 36000
rect 13847 35965 13881 35999
rect 13919 35964 13953 35998
rect 13991 35964 14019 35998
rect 14019 35964 14025 35998
rect 13775 35893 13781 35927
rect 13781 35893 13809 35927
rect 13847 35892 13881 35926
rect 13919 35891 13953 35925
rect 13991 35891 14019 35925
rect 14019 35891 14025 35925
rect 13775 35820 13781 35854
rect 13781 35820 13809 35854
rect 13847 35819 13881 35853
rect 13919 35818 13953 35852
rect 13991 35818 14019 35852
rect 14019 35818 14025 35852
rect 13775 35747 13781 35781
rect 13781 35747 13809 35781
rect 13847 35746 13881 35780
rect 13919 35745 13953 35779
rect 13991 35745 14019 35779
rect 14019 35745 14025 35779
rect 13775 35674 13781 35708
rect 13781 35674 13809 35708
rect 13847 35673 13881 35707
rect 13919 35672 13953 35706
rect 13991 35672 14019 35706
rect 14019 35672 14025 35706
rect 13775 35601 13781 35635
rect 13781 35601 13809 35635
rect 13847 35600 13881 35634
rect 13919 35599 13953 35633
rect 13991 35599 14019 35633
rect 14019 35599 14025 35633
rect 13775 35528 13781 35562
rect 13781 35528 13809 35562
rect 13847 35527 13881 35561
rect 13919 35526 13953 35560
rect 13991 35526 14019 35560
rect 14019 35526 14025 35560
rect 13775 35455 13781 35489
rect 13781 35455 13809 35489
rect 13847 35454 13881 35488
rect 13919 35453 13953 35487
rect 13991 35453 14019 35487
rect 14019 35453 14025 35487
rect 13775 35382 13781 35416
rect 13781 35382 13809 35416
rect 13847 35381 13881 35415
rect 13919 35380 13953 35414
rect 13991 35380 14019 35414
rect 14019 35380 14025 35414
rect 13775 35309 13781 35343
rect 13781 35309 13809 35343
rect 13847 35308 13881 35342
rect 13919 35307 13953 35341
rect 13991 35307 14019 35341
rect 14019 35307 14025 35341
rect 13775 35236 13781 35270
rect 13781 35236 13809 35270
rect 13847 35235 13881 35269
rect 13919 35234 13953 35268
rect 13991 35234 14019 35268
rect 14019 35234 14025 35268
rect 13775 35163 13781 35197
rect 13781 35163 13809 35197
rect 13847 35162 13881 35196
rect 13919 35161 13953 35195
rect 13991 35161 14019 35195
rect 14019 35161 14025 35195
rect 13775 35090 13781 35124
rect 13781 35090 13809 35124
rect 13847 35089 13881 35123
rect 13775 35017 13781 35051
rect 13781 35017 13809 35051
rect 13919 35050 14019 35122
rect 13847 34978 14019 35050
rect 13507 33084 13541 33118
rect 13597 33084 13628 33118
rect 13628 33084 13631 33118
rect 13507 33012 13541 33046
rect 13597 33012 13628 33046
rect 13628 33012 13631 33046
rect 13507 32940 13541 32974
rect 13597 32940 13628 32974
rect 13628 32940 13631 32974
rect 13507 32868 13541 32902
rect 13597 32868 13628 32902
rect 13628 32868 13631 32902
rect 13507 32796 13541 32830
rect 13597 32796 13628 32830
rect 13628 32796 13631 32830
rect 13507 32724 13541 32758
rect 13597 32724 13628 32758
rect 13628 32724 13631 32758
rect 13507 32652 13541 32686
rect 13597 32652 13628 32686
rect 13628 32652 13631 32686
rect 13507 32580 13541 32614
rect 13597 32580 13628 32614
rect 13628 32580 13631 32614
rect 13507 32508 13541 32542
rect 13597 32508 13628 32542
rect 13628 32508 13631 32542
rect 13507 32436 13541 32470
rect 13597 32436 13628 32470
rect 13628 32436 13631 32470
rect 2494 32176 2528 32210
rect 2579 32176 2613 32210
rect 2664 32176 2698 32210
rect 2494 32104 2528 32138
rect 2579 32104 2613 32138
rect 2664 32104 2698 32138
rect 13507 32364 13541 32398
rect 13597 32364 13628 32398
rect 13628 32364 13631 32398
rect 13507 32292 13541 32326
rect 13597 32292 13628 32326
rect 13628 32292 13631 32326
rect 13507 32220 13541 32254
rect 13597 32220 13628 32254
rect 13628 32220 13631 32254
rect 13507 32148 13541 32182
rect 13597 32148 13628 32182
rect 13628 32148 13631 32182
rect 13507 32076 13541 32110
rect 13597 32076 13628 32110
rect 13628 32076 13631 32110
rect 13507 32004 13541 32038
rect 13597 32004 13628 32038
rect 13628 32004 13631 32038
rect 13507 31932 13541 31966
rect 13597 31932 13628 31966
rect 13628 31932 13631 31966
rect 13507 31860 13541 31894
rect 13597 31860 13628 31894
rect 13628 31860 13631 31894
rect 13507 31788 13541 31822
rect 13597 31788 13628 31822
rect 13628 31788 13631 31822
rect 2314 30381 2395 31783
rect 2395 30381 2420 31783
rect 2314 30308 2348 30342
rect 2386 30308 2395 30342
rect 2395 30308 2420 30342
rect 2314 30235 2348 30269
rect 2386 30235 2395 30269
rect 2395 30235 2420 30269
rect 2314 30162 2348 30196
rect 2386 30162 2395 30196
rect 2395 30162 2420 30196
rect 2314 30089 2348 30123
rect 2386 30089 2395 30123
rect 2395 30089 2420 30123
rect 2314 30016 2348 30050
rect 2386 30016 2395 30050
rect 2395 30016 2420 30050
rect 2314 29943 2348 29977
rect 2386 29943 2395 29977
rect 2395 29943 2420 29977
rect 2314 29870 2348 29904
rect 2386 29870 2395 29904
rect 2395 29870 2420 29904
rect 2314 29797 2348 29831
rect 2386 29797 2395 29831
rect 2395 29797 2420 29831
rect 2314 29724 2348 29758
rect 2386 29724 2395 29758
rect 2395 29724 2420 29758
rect 2314 29651 2348 29685
rect 2386 29651 2395 29685
rect 2395 29651 2420 29685
rect 2314 29578 2348 29612
rect 2386 29578 2395 29612
rect 2395 29578 2420 29612
rect 2314 29505 2348 29539
rect 2386 29505 2395 29539
rect 2395 29505 2420 29539
rect 2314 29432 2348 29466
rect 2386 29432 2395 29466
rect 2395 29432 2420 29466
rect 2314 29359 2348 29393
rect 2386 29359 2395 29393
rect 2395 29359 2420 29393
rect 2314 29286 2348 29320
rect 2386 29286 2395 29320
rect 2395 29286 2420 29320
rect 2314 29213 2348 29247
rect 2386 29213 2395 29247
rect 2395 29213 2420 29247
rect 2314 29140 2348 29174
rect 2386 29140 2395 29174
rect 2395 29140 2420 29174
rect 2314 29067 2348 29101
rect 2386 29067 2395 29101
rect 2395 29067 2420 29101
rect 2314 28994 2348 29028
rect 2386 28994 2395 29028
rect 2395 28994 2420 29028
rect 2314 28921 2348 28955
rect 2386 28921 2395 28955
rect 2395 28921 2420 28955
rect 2314 28848 2348 28882
rect 2386 28848 2395 28882
rect 2395 28848 2420 28882
rect 2314 28775 2348 28809
rect 2386 28775 2395 28809
rect 2395 28775 2420 28809
rect 2314 28702 2348 28736
rect 2386 28702 2395 28736
rect 2395 28702 2420 28736
rect 2314 28629 2348 28663
rect 2386 28629 2395 28663
rect 2395 28629 2420 28663
rect 2314 28556 2348 28590
rect 2386 28556 2395 28590
rect 2395 28556 2420 28590
rect 2314 28483 2348 28517
rect 2386 28483 2395 28517
rect 2395 28483 2420 28517
rect 2314 28410 2348 28444
rect 2386 28410 2395 28444
rect 2395 28410 2420 28444
rect 2314 28337 2348 28371
rect 2386 28337 2395 28371
rect 2395 28337 2420 28371
rect 2314 28264 2348 28298
rect 2386 28264 2395 28298
rect 2395 28264 2420 28298
rect 2314 28191 2348 28225
rect 2386 28191 2395 28225
rect 2395 28191 2420 28225
rect 2314 28118 2348 28152
rect 2386 28118 2395 28152
rect 2395 28118 2420 28152
rect 2314 28045 2348 28079
rect 2386 28045 2395 28079
rect 2395 28045 2420 28079
rect 2314 27972 2348 28006
rect 2386 27972 2395 28006
rect 2395 27972 2420 28006
rect 2314 27899 2348 27933
rect 2386 27899 2395 27933
rect 2395 27899 2420 27933
rect 2314 27826 2348 27860
rect 2386 27826 2395 27860
rect 2395 27826 2420 27860
rect 2877 28560 3055 31762
rect 2877 28487 2911 28521
rect 2949 28487 2983 28521
rect 3021 28487 3055 28521
rect 2877 28414 2911 28448
rect 2949 28414 2983 28448
rect 3021 28414 3055 28448
rect 2877 28341 2911 28375
rect 2949 28341 2983 28375
rect 3021 28341 3055 28375
rect 2877 28268 2911 28302
rect 2949 28268 2983 28302
rect 3021 28268 3055 28302
rect 2877 28195 2911 28229
rect 2949 28195 2983 28229
rect 3021 28195 3055 28229
rect 2877 28122 2911 28156
rect 2949 28122 2983 28156
rect 3021 28122 3055 28156
rect 2877 28049 2911 28083
rect 2949 28049 2983 28083
rect 3021 28049 3055 28083
rect 2877 27976 2911 28010
rect 2949 27976 2983 28010
rect 3021 27976 3055 28010
rect 2877 27903 2911 27937
rect 2949 27903 2983 27937
rect 3021 27903 3055 27937
rect 3797 28560 3975 31762
rect 3797 28487 3831 28521
rect 3869 28487 3903 28521
rect 3941 28487 3975 28521
rect 3797 28414 3831 28448
rect 3869 28414 3903 28448
rect 3941 28414 3975 28448
rect 3797 28341 3831 28375
rect 3869 28341 3903 28375
rect 3941 28341 3975 28375
rect 3797 28268 3831 28302
rect 3869 28268 3903 28302
rect 3941 28268 3975 28302
rect 3797 28195 3831 28229
rect 3869 28195 3903 28229
rect 3941 28195 3975 28229
rect 3797 28122 3831 28156
rect 3869 28122 3903 28156
rect 3941 28122 3975 28156
rect 3797 28049 3831 28083
rect 3869 28049 3903 28083
rect 3941 28049 3975 28083
rect 3797 27976 3831 28010
rect 3869 27976 3903 28010
rect 3941 27976 3975 28010
rect 3797 27903 3831 27937
rect 3869 27903 3903 27937
rect 3941 27903 3975 27937
rect 4717 27903 4895 31753
rect 5637 27903 5815 31753
rect 6557 27903 6735 31753
rect 7477 27903 7655 31753
rect 8397 27903 8575 31753
rect 9317 27903 9495 31753
rect 10237 27903 10415 31753
rect 11157 27903 11335 31753
rect 12077 27903 12255 31753
rect 12997 27903 13175 31753
rect 13507 31716 13541 31750
rect 13597 31716 13628 31750
rect 13628 31716 13631 31750
rect 13507 31644 13541 31678
rect 13597 31644 13628 31678
rect 13628 31644 13631 31678
rect 13507 31572 13541 31606
rect 13597 31572 13628 31606
rect 13628 31572 13631 31606
rect 13507 31500 13541 31534
rect 13597 31500 13628 31534
rect 13628 31500 13631 31534
rect 13507 31428 13541 31462
rect 13597 31428 13628 31462
rect 13628 31428 13631 31462
rect 13507 31356 13541 31390
rect 13597 31356 13628 31390
rect 13628 31356 13631 31390
rect 13507 31284 13541 31318
rect 13597 31284 13628 31318
rect 13628 31284 13631 31318
rect 13507 31212 13541 31246
rect 13597 31212 13628 31246
rect 13628 31212 13631 31246
rect 13507 31140 13541 31174
rect 13597 31140 13628 31174
rect 13628 31140 13631 31174
rect 13507 31068 13541 31102
rect 13597 31068 13628 31102
rect 13628 31068 13631 31102
rect 13507 30996 13541 31030
rect 13597 30996 13628 31030
rect 13628 30996 13631 31030
rect 13507 30924 13541 30958
rect 13597 30924 13628 30958
rect 13628 30924 13631 30958
rect 13507 30852 13541 30886
rect 13597 30852 13628 30886
rect 13628 30852 13631 30886
rect 13507 30780 13541 30814
rect 13597 30780 13628 30814
rect 13628 30780 13631 30814
rect 13507 30708 13541 30742
rect 13597 30708 13628 30742
rect 13628 30708 13631 30742
rect 13507 30636 13541 30670
rect 13597 30636 13628 30670
rect 13628 30636 13631 30670
rect 13507 30564 13541 30598
rect 13597 30564 13628 30598
rect 13628 30564 13631 30598
rect 13507 30492 13541 30526
rect 13597 30492 13628 30526
rect 13628 30492 13631 30526
rect 13507 30420 13541 30454
rect 13597 30420 13628 30454
rect 13628 30420 13631 30454
rect 13507 30348 13541 30382
rect 13597 30348 13628 30382
rect 13628 30348 13631 30382
rect 13507 30276 13541 30310
rect 13597 30276 13628 30310
rect 13628 30276 13631 30310
rect 13507 30204 13541 30238
rect 13597 30204 13628 30238
rect 13628 30204 13631 30238
rect 13507 30132 13541 30166
rect 13597 30132 13628 30166
rect 13628 30132 13631 30166
rect 13507 30060 13541 30094
rect 13597 30060 13628 30094
rect 13628 30060 13631 30094
rect 13507 29988 13541 30022
rect 13597 29988 13628 30022
rect 13628 29988 13631 30022
rect 13507 29916 13541 29950
rect 13597 29916 13628 29950
rect 13628 29916 13631 29950
rect 13507 29844 13541 29878
rect 13597 29844 13628 29878
rect 13628 29844 13631 29878
rect 13507 29772 13541 29806
rect 13597 29772 13628 29806
rect 13628 29772 13631 29806
rect 13507 29700 13541 29734
rect 13597 29700 13628 29734
rect 13628 29700 13631 29734
rect 13507 29628 13541 29662
rect 13597 29628 13628 29662
rect 13628 29628 13631 29662
rect 13507 29556 13541 29590
rect 13597 29556 13628 29590
rect 13628 29556 13631 29590
rect 13507 29484 13541 29518
rect 13597 29484 13628 29518
rect 13628 29484 13631 29518
rect 13507 29412 13541 29446
rect 13597 29412 13628 29446
rect 13628 29412 13631 29446
rect 13507 29340 13541 29374
rect 13597 29340 13628 29374
rect 13628 29340 13631 29374
rect 13507 29268 13541 29302
rect 13597 29268 13628 29302
rect 13628 29268 13631 29302
rect 13507 29196 13541 29230
rect 13597 29196 13628 29230
rect 13628 29196 13631 29230
rect 13507 29124 13541 29158
rect 13597 29124 13628 29158
rect 13628 29124 13631 29158
rect 13507 29052 13541 29086
rect 13597 29052 13628 29086
rect 13628 29052 13631 29086
rect 13507 28980 13541 29014
rect 13597 28980 13628 29014
rect 13628 28980 13631 29014
rect 13507 28908 13541 28942
rect 13597 28908 13628 28942
rect 13628 28908 13631 28942
rect 13507 28836 13541 28870
rect 13597 28836 13628 28870
rect 13628 28836 13631 28870
rect 13507 28764 13541 28798
rect 13597 28764 13628 28798
rect 13628 28764 13631 28798
rect 13507 28692 13541 28726
rect 13597 28692 13628 28726
rect 13628 28692 13631 28726
rect 13507 28620 13541 28654
rect 13597 28620 13628 28654
rect 13628 28620 13631 28654
rect 13507 28548 13541 28582
rect 13597 28548 13628 28582
rect 13628 28548 13631 28582
rect 13507 28476 13541 28510
rect 13597 28476 13628 28510
rect 13628 28476 13631 28510
rect 13507 28404 13541 28438
rect 13597 28404 13628 28438
rect 13628 28404 13631 28438
rect 13507 28332 13541 28366
rect 13597 28332 13628 28366
rect 13628 28332 13631 28366
rect 13507 28260 13541 28294
rect 13597 28260 13628 28294
rect 13628 28260 13631 28294
rect 13507 28188 13541 28222
rect 13597 28188 13628 28222
rect 13628 28188 13631 28222
rect 13507 28116 13541 28150
rect 13597 28116 13628 28150
rect 13628 28116 13631 28150
rect 13507 28044 13541 28078
rect 13597 28044 13628 28078
rect 13628 28044 13631 28078
rect 13507 27972 13541 28006
rect 13597 27972 13628 28006
rect 13628 27972 13631 28006
rect 13507 27900 13541 27934
rect 13597 27900 13628 27934
rect 13628 27900 13631 27934
rect 13507 27828 13541 27862
rect 13597 27828 13628 27862
rect 13628 27828 13631 27862
rect 2314 27753 2348 27787
rect 2386 27753 2395 27787
rect 2395 27753 2420 27787
rect 2314 27680 2348 27714
rect 2386 27680 2395 27714
rect 2395 27680 2420 27714
rect 2314 27607 2348 27641
rect 2386 27607 2395 27641
rect 2395 27607 2420 27641
rect 2314 27534 2348 27568
rect 2386 27534 2395 27568
rect 2395 27534 2420 27568
rect 2314 27461 2348 27495
rect 2386 27461 2395 27495
rect 2395 27461 2420 27495
rect 2314 27388 2348 27422
rect 2386 27388 2395 27422
rect 2395 27388 2420 27422
rect 2314 27315 2348 27349
rect 2386 27315 2395 27349
rect 2395 27315 2420 27349
rect 3170 27540 3204 27574
rect 3245 27540 3279 27574
rect 3320 27540 3354 27574
rect 2314 27268 2348 27276
rect 2386 27268 2395 27276
rect 2395 27268 2420 27276
rect 13507 27756 13541 27790
rect 13597 27756 13628 27790
rect 13628 27756 13631 27790
rect 13507 27684 13541 27718
rect 13597 27684 13628 27718
rect 13628 27684 13631 27718
rect 13507 27612 13541 27646
rect 13597 27612 13628 27646
rect 13628 27612 13631 27646
rect 13507 27540 13541 27574
rect 13597 27540 13628 27574
rect 13628 27540 13631 27574
rect 13507 27468 13541 27502
rect 13597 27468 13628 27502
rect 13628 27468 13631 27502
rect 13507 27396 13541 27430
rect 13597 27396 13628 27430
rect 13628 27396 13631 27430
rect 13507 27324 13541 27358
rect 13597 27324 13628 27358
rect 13628 27324 13631 27358
rect 2314 27242 2327 27268
rect 2327 27242 2348 27268
rect 2386 27242 2420 27268
rect 13507 27252 13541 27286
rect 13597 27252 13628 27286
rect 13628 27252 13631 27286
rect 2314 27200 2327 27203
rect 2327 27200 2348 27203
rect 2314 27169 2348 27200
rect 2386 27169 2420 27203
rect 2471 27169 2505 27203
rect 2550 27169 2584 27203
rect 2629 27169 2663 27203
rect 2708 27169 2742 27203
rect 2787 27169 2821 27203
rect 3584 27197 3618 27231
rect 3662 27197 3696 27231
rect 3740 27197 3774 27231
rect 3818 27197 3852 27231
rect 3896 27197 3930 27231
rect 3974 27197 4008 27231
rect 4052 27197 4086 27231
rect 4130 27197 4164 27231
rect 4208 27197 4242 27231
rect 4286 27197 4320 27231
rect 4363 27197 4367 27231
rect 4367 27197 4397 27231
rect 2392 27097 2426 27131
rect 2471 27097 2505 27131
rect 2550 27097 2584 27131
rect 2629 27097 2663 27131
rect 2708 27097 2742 27131
rect 2787 27097 2821 27131
rect 3584 27089 3618 27123
rect 3662 27089 3696 27123
rect 3740 27089 3774 27123
rect 3818 27089 3852 27123
rect 3896 27089 3930 27123
rect 3974 27089 4008 27123
rect 4052 27089 4086 27123
rect 4130 27089 4164 27123
rect 4208 27089 4242 27123
rect 4286 27089 4299 27123
rect 4299 27089 4320 27123
rect 4363 27097 4397 27123
rect 4363 27089 4397 27097
rect 1840 27005 1874 27039
rect 1946 26966 1980 27000
rect 1840 26932 1874 26966
rect 1946 26911 1980 26927
rect 1946 26893 1980 26911
rect 1840 26859 1874 26893
rect 1946 26840 1980 26854
rect 1946 26820 1970 26840
rect 1970 26820 1980 26840
rect 1840 26809 1874 26820
rect 1840 26786 1868 26809
rect 1868 26786 1874 26809
rect 1946 26772 1970 26781
rect 1970 26772 1980 26781
rect 1946 26747 1980 26772
rect 2024 26747 2058 26781
rect 2102 26747 2136 26781
rect 2180 26747 2214 26781
rect 2258 26747 2292 26781
rect 2336 26747 2370 26781
rect 2414 26747 2448 26781
rect 2492 26747 2526 26781
rect 2570 26747 2604 26781
rect 2648 26747 2682 26781
rect 2726 26747 2760 26781
rect 2804 26747 2838 26781
rect 1840 26713 1874 26747
rect 3567 26735 3601 26769
rect 3643 26735 3677 26769
rect 3719 26735 3753 26769
rect 3795 26735 3829 26769
rect 3871 26735 3905 26769
rect 3947 26738 3976 26769
rect 3976 26738 3981 26769
rect 3947 26735 3981 26738
rect 1914 26670 1948 26675
rect 1988 26670 2022 26675
rect 2062 26670 2096 26675
rect 2136 26670 2170 26675
rect 2210 26670 2244 26675
rect 2284 26670 2318 26675
rect 2358 26670 2392 26675
rect 2432 26670 2466 26675
rect 2506 26670 2540 26675
rect 2580 26670 2614 26675
rect 2654 26670 2688 26675
rect 2729 26670 2763 26675
rect 2804 26670 2838 26675
rect 1914 26641 1948 26670
rect 1988 26641 2022 26670
rect 2062 26641 2096 26670
rect 2136 26641 2170 26670
rect 2210 26641 2244 26670
rect 2284 26641 2318 26670
rect 2358 26641 2392 26670
rect 2432 26641 2466 26670
rect 2506 26641 2540 26670
rect 2580 26641 2614 26670
rect 2654 26641 2688 26670
rect 2729 26641 2763 26670
rect 2804 26641 2838 26670
rect 4019 26663 4053 26697
rect 3567 26629 3601 26663
rect 3653 26629 3687 26663
rect 3739 26629 3773 26663
rect 3826 26629 3860 26663
rect 3913 26629 3947 26663
rect 4019 26591 4053 26625
rect 3913 26557 3947 26591
rect 4019 26519 4053 26553
rect 3913 26485 3947 26519
rect 4019 26447 4053 26481
rect 3913 26413 3947 26447
rect 4019 26375 4053 26409
rect 3913 26341 3947 26375
rect 4019 26303 4053 26337
rect 3913 26269 3947 26303
rect 4019 26231 4053 26265
rect 3913 26197 3947 26231
rect 4019 26159 4053 26193
rect 3913 26125 3947 26159
rect 4019 26087 4053 26121
rect 3913 26053 3947 26087
rect 4019 26015 4053 26049
rect 3913 25981 3947 26015
rect 4019 25943 4053 25977
rect 3913 25909 3947 25943
rect 4019 25871 4053 25905
rect 3913 25837 3947 25871
rect 4019 25799 4053 25833
rect 3913 25765 3947 25799
rect 4019 25727 4053 25761
rect 3913 25693 3947 25727
rect 4019 25655 4053 25689
rect 3913 25621 3947 25655
rect 4019 25583 4053 25617
rect 3913 25549 3947 25583
rect 4019 25511 4053 25545
rect 3913 25477 3947 25511
rect 4019 25439 4053 25473
rect 3913 25405 3947 25439
rect 4019 25367 4053 25401
rect 3913 25333 3947 25367
rect 4019 25295 4053 25329
rect 3913 25261 3947 25295
rect 4019 25223 4053 25257
rect 3913 25189 3947 25223
rect 4019 25151 4053 25185
rect 3913 25117 3947 25151
rect 4019 25079 4053 25113
rect 3913 25045 3947 25079
rect 4019 25007 4053 25041
rect 3913 24973 3947 25007
rect 4019 24935 4053 24969
rect 3913 24901 3947 24935
rect 4019 24863 4053 24897
rect 3913 24829 3947 24863
rect 4019 24791 4053 24825
rect 3913 24757 3947 24791
rect 4019 24719 4053 24753
rect 3913 24685 3947 24719
rect 4019 24647 4053 24681
rect 3913 24613 3947 24647
rect 4019 24575 4053 24609
rect 3913 24541 3947 24575
rect 4019 24503 4053 24537
rect 3913 24469 3947 24503
rect 4019 24431 4053 24465
rect 3913 24397 3947 24431
rect 4019 24359 4053 24393
rect 3913 24325 3947 24359
rect 4019 24287 4053 24321
rect 3913 24253 3947 24287
rect 4019 24215 4053 24249
rect 3913 24181 3947 24215
rect 4019 24143 4053 24177
rect 3913 24109 3947 24143
rect 4019 24071 4053 24105
rect 3913 24037 3947 24071
rect 4019 23999 4053 24033
rect 3913 23965 3947 23999
rect 4019 23927 4053 23961
rect 3913 23893 3947 23927
rect 4019 23855 4053 23889
rect 3913 23821 3947 23855
rect 4019 23783 4053 23817
rect 3913 23749 3947 23783
rect 4019 23711 4053 23745
rect 3913 23677 3947 23711
rect 4019 23639 4053 23673
rect 3913 23605 3947 23639
rect 4019 23567 4053 23601
rect 3913 23533 3947 23567
rect 4019 23495 4053 23529
rect 3913 23461 3947 23495
rect 4019 23423 4053 23457
rect 3913 23389 3947 23423
rect 4019 23351 4053 23385
rect 3913 23317 3947 23351
rect 4019 23279 4053 23313
rect 3913 23245 3947 23279
rect 4019 23207 4053 23241
rect 3913 23173 3947 23207
rect 4019 23135 4053 23169
rect 3913 23101 3947 23135
rect 4019 23063 4053 23097
rect 3913 23029 3947 23063
rect 4019 22991 4053 23025
rect 3913 22957 3947 22991
rect 4019 22919 4053 22953
rect 3913 22885 3947 22919
rect 4019 22847 4053 22881
rect 3913 22813 3947 22847
rect 4019 22775 4053 22809
rect 3913 22741 3947 22775
rect 4019 22703 4053 22737
rect 3913 22669 3947 22703
rect 4019 22631 4053 22665
rect 3913 22597 3947 22631
rect 4019 22559 4053 22593
rect 3913 22525 3947 22559
rect 4019 22487 4053 22521
rect 3913 22453 3947 22487
rect 4019 22415 4053 22449
rect 3913 22381 3947 22415
rect 4019 22343 4053 22377
rect 3913 22309 3947 22343
rect 4019 22271 4053 22305
rect 3913 22237 3947 22271
rect 4019 22199 4053 22233
rect 3913 22165 3947 22199
rect 4019 22127 4053 22161
rect 3913 22093 3947 22127
rect 4019 22055 4053 22089
rect 3913 22021 3947 22055
rect 3913 21949 3947 21983
rect 4019 21982 4053 22016
rect 3913 21877 3947 21911
rect 4019 21909 4053 21943
rect 3913 21805 3947 21839
rect 4019 21836 4053 21870
rect 3913 21733 3947 21767
rect 4019 21763 4053 21797
rect 3913 21661 3947 21695
rect 4019 21690 4053 21724
rect 3913 21589 3947 21623
rect 4019 21617 4053 21651
rect 3913 21517 3947 21551
rect 4019 21544 4053 21578
rect 3913 21445 3947 21479
rect 4019 21471 4053 21505
rect 3913 21373 3947 21407
rect 4019 21398 4053 21432
rect 3913 21301 3947 21335
rect 4019 21325 4053 21359
rect 3913 21229 3947 21263
rect 4019 21252 4053 21286
rect 3913 21157 3947 21191
rect 4019 21179 4053 21213
rect 3913 21085 3947 21119
rect 4019 21106 4053 21140
rect 3913 21013 3947 21047
rect 4019 21033 4053 21067
rect 3913 20941 3947 20975
rect 4019 20960 4053 20994
rect 3913 20869 3947 20903
rect 4019 20887 4053 20921
rect 3913 20797 3947 20831
rect 4019 20814 4053 20848
rect 3913 20725 3947 20759
rect 4019 20741 4053 20775
rect 3913 20653 3947 20687
rect 4019 20668 4053 20702
rect 3913 20581 3947 20615
rect 4019 20595 4053 20629
rect 3913 20509 3947 20543
rect 4019 20522 4053 20556
rect 3913 20437 3947 20471
rect 4019 20449 4053 20483
rect 3913 20365 3947 20399
rect 4019 20376 4053 20410
rect 3913 20293 3947 20327
rect 4019 20303 4053 20337
rect 3913 20221 3947 20255
rect 4019 20230 4053 20264
rect 3913 20149 3947 20183
rect 4019 20157 4053 20191
rect 3913 20077 3947 20111
rect 4019 20084 4053 20118
rect 3913 20005 3947 20039
rect 4019 20011 4053 20045
rect 3913 19933 3947 19967
rect 4019 19938 4053 19972
rect 3913 19861 3947 19895
rect 4019 19865 4053 19899
rect 3913 19789 3947 19823
rect 4019 19792 4053 19826
rect 3913 19717 3947 19751
rect 4019 19719 4053 19753
rect 3913 19645 3947 19679
rect 4019 19646 4053 19680
rect 3913 19573 3947 19607
rect 4019 19573 4053 19607
rect 3913 19500 3947 19534
rect 4019 19500 4053 19534
rect 4365 23557 4471 27047
rect 4365 23484 4399 23518
rect 4437 23484 4471 23518
rect 4365 23411 4399 23445
rect 4437 23411 4471 23445
rect 4365 23338 4399 23372
rect 4437 23338 4471 23372
rect 4365 23265 4399 23299
rect 4437 23265 4471 23299
rect 4783 27128 4817 27162
rect 4861 27128 4895 27162
rect 4783 27055 4817 27089
rect 4861 27055 4895 27089
rect 4783 26982 4817 27016
rect 4861 26982 4895 27016
rect 4783 26909 4817 26943
rect 4861 26909 4895 26943
rect 4783 26836 4817 26870
rect 4861 26836 4895 26870
rect 4783 26763 4817 26797
rect 4861 26763 4895 26797
rect 4783 26690 4817 26724
rect 4861 26690 4895 26724
rect 4783 26617 4817 26651
rect 4861 26617 4895 26651
rect 4783 26544 4817 26578
rect 4861 26544 4895 26578
rect 4783 26471 4817 26505
rect 4861 26471 4895 26505
rect 4783 26398 4817 26432
rect 4861 26398 4895 26432
rect 4783 26325 4817 26359
rect 4861 26325 4895 26359
rect 4783 26252 4817 26286
rect 4861 26252 4895 26286
rect 4783 26179 4817 26213
rect 4861 26179 4895 26213
rect 4783 26106 4817 26140
rect 4861 26106 4895 26140
rect 4783 26033 4817 26067
rect 4861 26033 4895 26067
rect 4783 25960 4817 25994
rect 4861 25960 4895 25994
rect 4783 25887 4817 25921
rect 4861 25887 4895 25921
rect 4783 25814 4817 25848
rect 4861 25814 4895 25848
rect 4783 25741 4817 25775
rect 4861 25741 4895 25775
rect 4783 25668 4817 25702
rect 4861 25668 4895 25702
rect 4783 25595 4817 25629
rect 4861 25595 4895 25629
rect 4783 25522 4817 25556
rect 4861 25522 4895 25556
rect 4783 25449 4817 25483
rect 4861 25449 4895 25483
rect 4783 25376 4817 25410
rect 4861 25376 4895 25410
rect 4783 25303 4817 25337
rect 4861 25303 4895 25337
rect 4783 25230 4817 25264
rect 4861 25230 4895 25264
rect 4783 25157 4817 25191
rect 4861 25157 4895 25191
rect 4783 25084 4817 25118
rect 4861 25084 4895 25118
rect 4783 25011 4817 25045
rect 4861 25011 4895 25045
rect 4783 24938 4817 24972
rect 4861 24938 4895 24972
rect 4783 24865 4817 24899
rect 4861 24865 4895 24899
rect 4783 24792 4817 24826
rect 4861 24792 4895 24826
rect 4783 24719 4817 24753
rect 4861 24719 4895 24753
rect 4783 24646 4817 24680
rect 4861 24646 4895 24680
rect 4783 24572 4817 24606
rect 4861 24572 4895 24606
rect 4783 24498 4817 24532
rect 4861 24498 4895 24532
rect 4783 24424 4817 24458
rect 4861 24424 4895 24458
rect 4783 24350 4817 24384
rect 4861 24350 4895 24384
rect 4783 24276 4817 24310
rect 4861 24276 4895 24310
rect 4783 24202 4817 24236
rect 4861 24202 4895 24236
rect 4783 24128 4817 24162
rect 4861 24128 4895 24162
rect 4783 24054 4817 24088
rect 4861 24054 4895 24088
rect 4783 23980 4817 24014
rect 4861 23980 4895 24014
rect 4783 23906 4817 23940
rect 4861 23906 4895 23940
rect 4783 23832 4817 23866
rect 4861 23832 4895 23866
rect 4783 23758 4817 23792
rect 4861 23758 4895 23792
rect 4783 23684 4817 23718
rect 4861 23684 4895 23718
rect 4783 23610 4817 23644
rect 4861 23610 4895 23644
rect 4783 23536 4817 23570
rect 4861 23536 4895 23570
rect 4783 23462 4817 23496
rect 4861 23462 4895 23496
rect 4783 23388 4817 23422
rect 4861 23388 4895 23422
rect 4783 23314 4817 23348
rect 4861 23314 4895 23348
rect 5637 23960 5815 27162
rect 5637 23887 5671 23921
rect 5709 23887 5743 23921
rect 5781 23887 5815 23921
rect 5637 23814 5671 23848
rect 5709 23814 5743 23848
rect 5781 23814 5815 23848
rect 5637 23741 5671 23775
rect 5709 23741 5743 23775
rect 5781 23741 5815 23775
rect 5637 23668 5671 23702
rect 5709 23668 5743 23702
rect 5781 23668 5815 23702
rect 5637 23595 5671 23629
rect 5709 23595 5743 23629
rect 5781 23595 5815 23629
rect 5637 23522 5671 23556
rect 5709 23522 5743 23556
rect 5781 23522 5815 23556
rect 5637 23449 5671 23483
rect 5709 23449 5743 23483
rect 5781 23449 5815 23483
rect 5637 23376 5671 23410
rect 5709 23376 5743 23410
rect 5781 23376 5815 23410
rect 5637 23303 5671 23337
rect 5709 23303 5743 23337
rect 5781 23303 5815 23337
rect 6557 23303 6735 27153
rect 7477 23303 7655 27153
rect 8397 23303 8575 27153
rect 9317 23303 9495 27153
rect 10237 23303 10415 27153
rect 11157 23303 11335 27153
rect 12077 23303 12255 27153
rect 12997 23303 13175 27153
rect 13507 27180 13541 27214
rect 13597 27180 13628 27214
rect 13628 27180 13631 27214
rect 13507 27108 13541 27142
rect 13597 27108 13628 27142
rect 13628 27108 13631 27142
rect 13507 27036 13541 27070
rect 13597 27036 13628 27070
rect 13628 27036 13631 27070
rect 13507 26964 13541 26998
rect 13597 26964 13628 26998
rect 13628 26964 13631 26998
rect 13507 26892 13541 26926
rect 13597 26892 13628 26926
rect 13628 26892 13631 26926
rect 13507 26820 13541 26854
rect 13597 26820 13628 26854
rect 13628 26820 13631 26854
rect 13507 26748 13541 26782
rect 13597 26748 13628 26782
rect 13628 26748 13631 26782
rect 13507 26676 13541 26710
rect 13597 26676 13628 26710
rect 13628 26676 13631 26710
rect 13507 26604 13541 26638
rect 13597 26604 13628 26638
rect 13628 26604 13631 26638
rect 13507 26532 13541 26566
rect 13597 26532 13628 26566
rect 13628 26532 13631 26566
rect 13507 26460 13541 26494
rect 13597 26460 13628 26494
rect 13628 26460 13631 26494
rect 13507 26388 13541 26422
rect 13597 26388 13628 26422
rect 13628 26388 13631 26422
rect 13507 26316 13541 26350
rect 13597 26316 13628 26350
rect 13628 26316 13631 26350
rect 13507 26244 13541 26278
rect 13597 26244 13628 26278
rect 13628 26244 13631 26278
rect 13507 26172 13541 26206
rect 13597 26172 13628 26206
rect 13628 26172 13631 26206
rect 13507 26100 13541 26134
rect 13597 26100 13628 26134
rect 13628 26100 13631 26134
rect 13507 26028 13541 26062
rect 13597 26028 13628 26062
rect 13628 26028 13631 26062
rect 13507 25956 13541 25990
rect 13597 25956 13628 25990
rect 13628 25956 13631 25990
rect 13507 25884 13541 25918
rect 13597 25884 13628 25918
rect 13628 25884 13631 25918
rect 13507 25812 13541 25846
rect 13597 25812 13628 25846
rect 13628 25812 13631 25846
rect 13507 25740 13541 25774
rect 13597 25740 13628 25774
rect 13628 25740 13631 25774
rect 13507 25668 13541 25702
rect 13597 25668 13628 25702
rect 13628 25668 13631 25702
rect 13507 25596 13541 25630
rect 13597 25596 13628 25630
rect 13628 25596 13631 25630
rect 13507 25524 13541 25558
rect 13597 25524 13628 25558
rect 13628 25524 13631 25558
rect 13507 25452 13541 25486
rect 13597 25452 13628 25486
rect 13628 25452 13631 25486
rect 13507 25379 13541 25413
rect 13597 25379 13628 25413
rect 13628 25379 13631 25413
rect 13507 25306 13541 25340
rect 13597 25306 13628 25340
rect 13628 25306 13631 25340
rect 13507 25233 13541 25267
rect 13597 25233 13628 25267
rect 13628 25233 13631 25267
rect 13507 25160 13541 25194
rect 13597 25160 13628 25194
rect 13628 25160 13631 25194
rect 13507 25087 13541 25121
rect 13597 25087 13628 25121
rect 13628 25087 13631 25121
rect 13507 25014 13541 25048
rect 13597 25014 13628 25048
rect 13628 25014 13631 25048
rect 13507 24941 13541 24975
rect 13597 24941 13628 24975
rect 13628 24941 13631 24975
rect 13507 24868 13541 24902
rect 13597 24868 13628 24902
rect 13628 24868 13631 24902
rect 13507 24795 13541 24829
rect 13597 24795 13628 24829
rect 13628 24795 13631 24829
rect 13507 24722 13541 24756
rect 13597 24722 13628 24756
rect 13628 24722 13631 24756
rect 13507 24649 13541 24683
rect 13597 24649 13628 24683
rect 13628 24649 13631 24683
rect 13507 24576 13541 24610
rect 13597 24576 13628 24610
rect 13628 24576 13631 24610
rect 13507 24503 13541 24537
rect 13597 24503 13628 24537
rect 13628 24503 13631 24537
rect 13507 24430 13541 24464
rect 13597 24430 13628 24464
rect 13628 24430 13631 24464
rect 13507 24357 13541 24391
rect 13597 24357 13628 24391
rect 13628 24357 13631 24391
rect 13507 24284 13541 24318
rect 13597 24284 13628 24318
rect 13628 24284 13631 24318
rect 13507 24211 13541 24245
rect 13597 24211 13628 24245
rect 13628 24211 13631 24245
rect 13507 24138 13541 24172
rect 13597 24138 13628 24172
rect 13628 24138 13631 24172
rect 13507 24065 13541 24099
rect 13597 24065 13628 24099
rect 13628 24065 13631 24099
rect 13507 23992 13541 24026
rect 13597 23992 13628 24026
rect 13628 23992 13631 24026
rect 13507 23919 13541 23953
rect 13597 23919 13628 23953
rect 13628 23919 13631 23953
rect 13507 23846 13541 23880
rect 13597 23846 13628 23880
rect 13628 23846 13631 23880
rect 13507 23773 13541 23807
rect 13597 23773 13628 23807
rect 13628 23773 13631 23807
rect 13507 23700 13541 23734
rect 13597 23700 13628 23734
rect 13628 23700 13631 23734
rect 13507 23627 13541 23661
rect 13597 23627 13628 23661
rect 13628 23627 13631 23661
rect 13507 23554 13541 23588
rect 13597 23554 13628 23588
rect 13628 23554 13631 23588
rect 13507 23481 13541 23515
rect 13597 23481 13628 23515
rect 13628 23481 13631 23515
rect 13507 23408 13541 23442
rect 13597 23408 13628 23442
rect 13628 23408 13631 23442
rect 13507 23335 13541 23369
rect 13597 23335 13628 23369
rect 13628 23335 13631 23369
rect 13507 23262 13541 23296
rect 13597 23262 13628 23296
rect 13628 23262 13631 23296
rect 4365 23192 4399 23226
rect 4437 23192 4471 23226
rect 4365 23119 4399 23153
rect 4437 23119 4471 23153
rect 4365 23046 4399 23080
rect 4437 23046 4471 23080
rect 4365 22973 4399 23007
rect 4437 22973 4471 23007
rect 4365 22900 4399 22934
rect 4437 22900 4471 22934
rect 4365 22827 4399 22861
rect 4437 22827 4471 22861
rect 4365 22754 4399 22788
rect 4437 22754 4471 22788
rect 4365 22681 4399 22715
rect 4437 22681 4471 22715
rect 4789 22959 4823 22993
rect 4789 22887 4823 22921
rect 13507 23189 13541 23223
rect 13597 23189 13628 23223
rect 13628 23189 13631 23223
rect 13507 23116 13541 23150
rect 13597 23116 13628 23150
rect 13628 23116 13631 23150
rect 13507 23043 13541 23077
rect 13597 23043 13628 23077
rect 13628 23043 13631 23077
rect 13507 22970 13541 23004
rect 13597 22970 13628 23004
rect 13628 22970 13631 23004
rect 13507 22897 13541 22931
rect 13597 22897 13628 22931
rect 13628 22897 13631 22931
rect 13507 22824 13541 22858
rect 13597 22824 13628 22858
rect 13628 22824 13631 22858
rect 13507 22751 13541 22785
rect 13597 22751 13628 22785
rect 13628 22751 13631 22785
rect 13507 22678 13541 22712
rect 13597 22678 13628 22712
rect 13628 22678 13631 22712
rect 4365 22608 4399 22642
rect 4437 22608 4471 22642
rect 13507 22605 13541 22639
rect 13597 22605 13628 22639
rect 13628 22605 13631 22639
rect 4365 22535 4399 22569
rect 4437 22535 4471 22569
rect 4365 22462 4399 22496
rect 4437 22462 4471 22496
rect 4365 22389 4399 22423
rect 4437 22389 4471 22423
rect 4365 22316 4399 22350
rect 4437 22316 4471 22350
rect 4365 22243 4399 22277
rect 4437 22243 4471 22277
rect 4365 22170 4399 22204
rect 4437 22170 4471 22204
rect 4365 22097 4399 22131
rect 4437 22097 4471 22131
rect 4365 22024 4399 22058
rect 4437 22024 4471 22058
rect 4365 21951 4399 21985
rect 4437 21951 4471 21985
rect 4365 21878 4399 21912
rect 4437 21878 4471 21912
rect 4365 21805 4399 21839
rect 4437 21805 4471 21839
rect 4365 21732 4399 21766
rect 4437 21732 4471 21766
rect 4365 21659 4399 21693
rect 4437 21659 4471 21693
rect 4365 21586 4399 21620
rect 4437 21586 4471 21620
rect 4365 21513 4399 21547
rect 4437 21513 4471 21547
rect 4365 21440 4399 21474
rect 4437 21440 4471 21474
rect 4365 21367 4399 21401
rect 4437 21367 4471 21401
rect 4365 21294 4399 21328
rect 4437 21294 4471 21328
rect 4365 21221 4399 21255
rect 4437 21221 4471 21255
rect 4365 21148 4399 21182
rect 4437 21148 4471 21182
rect 4365 21075 4399 21109
rect 4437 21075 4471 21109
rect 4365 21002 4399 21036
rect 4437 21002 4471 21036
rect 4365 20929 4399 20963
rect 4437 20929 4471 20963
rect 4365 20856 4399 20890
rect 4437 20856 4471 20890
rect 4365 20783 4399 20817
rect 4437 20783 4471 20817
rect 4365 20710 4399 20744
rect 4437 20710 4471 20744
rect 4365 20637 4399 20671
rect 4437 20637 4471 20671
rect 4365 20564 4399 20598
rect 4437 20564 4471 20598
rect 4365 20491 4399 20525
rect 4437 20491 4471 20525
rect 4365 20418 4399 20452
rect 4437 20418 4471 20452
rect 4365 20345 4399 20379
rect 4437 20345 4471 20379
rect 4365 20272 4399 20306
rect 4437 20272 4471 20306
rect 4365 20199 4399 20233
rect 4437 20199 4471 20233
rect 4365 20126 4399 20160
rect 4437 20126 4471 20160
rect 4365 20053 4399 20087
rect 4437 20053 4471 20087
rect 4365 19980 4399 20014
rect 4437 19980 4471 20014
rect 4365 19907 4399 19941
rect 4437 19907 4471 19941
rect 4365 19834 4399 19868
rect 4437 19834 4471 19868
rect 4365 19761 4399 19795
rect 4437 19761 4471 19795
rect 4365 19688 4399 19722
rect 4437 19688 4471 19722
rect 4365 19615 4399 19649
rect 4437 19615 4471 19649
rect 4365 19542 4399 19576
rect 4437 19542 4471 19576
rect 3967 19129 4198 19379
rect 3967 19056 4001 19090
rect 4039 19057 4198 19129
rect 3967 18983 4001 19017
rect 4039 18984 4073 19018
rect 4111 18985 4198 19057
rect 4198 18985 4217 19379
rect 3967 18910 4001 18944
rect 4039 18911 4073 18945
rect 4111 18912 4145 18946
rect 4183 18912 4198 18946
rect 4198 18912 4217 18946
rect 3967 18837 4001 18871
rect 4039 18838 4073 18872
rect 4111 18839 4145 18873
rect 4183 18839 4198 18873
rect 4198 18839 4217 18873
rect 3967 18764 4001 18798
rect 4039 18765 4073 18799
rect 4111 18766 4145 18800
rect 4183 18766 4198 18800
rect 4198 18766 4217 18800
rect 3967 18691 4001 18725
rect 4039 18692 4073 18726
rect 4111 18693 4145 18727
rect 4183 18693 4198 18727
rect 4198 18693 4217 18727
rect 3967 18618 4001 18652
rect 4039 18619 4073 18653
rect 4111 18620 4145 18654
rect 4183 18620 4198 18654
rect 4198 18620 4217 18654
rect 3967 18545 4001 18579
rect 4039 18546 4073 18580
rect 4111 18547 4145 18581
rect 4183 18547 4198 18581
rect 4198 18547 4217 18581
rect 3967 18472 4001 18506
rect 4039 18473 4073 18507
rect 4111 18474 4145 18508
rect 4183 18474 4198 18508
rect 4198 18474 4217 18508
rect 3967 18399 4001 18433
rect 4039 18400 4073 18434
rect 4111 18401 4145 18435
rect 4183 18401 4198 18435
rect 4198 18401 4217 18435
rect 3967 18326 4001 18360
rect 4039 18327 4073 18361
rect 4111 18328 4145 18362
rect 4183 18328 4198 18362
rect 4198 18328 4217 18362
rect 3967 18253 4001 18287
rect 4039 18254 4073 18288
rect 4111 18255 4145 18289
rect 4183 18255 4198 18289
rect 4198 18255 4217 18289
rect 3967 18180 4001 18214
rect 4039 18181 4073 18215
rect 4111 18182 4145 18216
rect 4183 18182 4198 18216
rect 4198 18182 4217 18216
rect 3967 18107 4001 18141
rect 4039 18108 4073 18142
rect 4111 18109 4145 18143
rect 4183 18109 4198 18143
rect 4198 18109 4217 18143
rect 3967 18034 4001 18068
rect 4039 18035 4073 18069
rect 4111 18036 4145 18070
rect 4183 18036 4198 18070
rect 4198 18036 4217 18070
rect 3967 17961 4001 17995
rect 4039 17962 4073 17996
rect 4111 17963 4145 17997
rect 4183 17963 4198 17997
rect 4198 17963 4217 17997
rect 3967 17888 4001 17922
rect 4039 17889 4073 17923
rect 4111 17890 4145 17924
rect 4183 17890 4198 17924
rect 4198 17890 4217 17924
rect 3967 17815 4001 17849
rect 4039 17816 4073 17850
rect 4111 17817 4145 17851
rect 4183 17817 4198 17851
rect 4198 17817 4217 17851
rect 3967 17742 4001 17776
rect 4039 17743 4073 17777
rect 4111 17744 4145 17778
rect 4183 17744 4198 17778
rect 4198 17744 4217 17778
rect 3967 17669 4001 17703
rect 4039 17670 4073 17704
rect 4111 17671 4145 17705
rect 4183 17671 4198 17705
rect 4198 17671 4217 17705
rect 3967 17596 4001 17630
rect 4039 17597 4073 17631
rect 4111 17598 4145 17632
rect 4183 17598 4198 17632
rect 4198 17598 4217 17632
rect 3967 17523 4001 17557
rect 4039 17524 4073 17558
rect 4111 17525 4145 17559
rect 4183 17525 4198 17559
rect 4198 17525 4217 17559
rect 3967 17450 4001 17484
rect 4039 17451 4073 17485
rect 4111 17452 4145 17486
rect 4183 17452 4198 17486
rect 4198 17452 4217 17486
rect 3967 17377 4001 17411
rect 4039 17378 4073 17412
rect 4111 17379 4145 17413
rect 4183 17379 4198 17413
rect 4198 17379 4217 17413
rect 3967 17304 4001 17338
rect 4039 17305 4073 17339
rect 4111 17306 4145 17340
rect 4183 17306 4198 17340
rect 4198 17306 4217 17340
rect 3967 17231 4001 17265
rect 4039 17232 4073 17266
rect 4111 17233 4145 17267
rect 4183 17233 4198 17267
rect 4198 17233 4217 17267
rect 3967 17158 4001 17192
rect 4039 17159 4073 17193
rect 4111 17160 4145 17194
rect 4183 17160 4198 17194
rect 4198 17160 4217 17194
rect 3967 17085 4001 17119
rect 4039 17086 4073 17120
rect 4111 17087 4145 17121
rect 4183 17087 4198 17121
rect 4198 17087 4217 17121
rect 3967 17012 4001 17046
rect 4039 17013 4073 17047
rect 4111 17014 4145 17048
rect 4183 17014 4198 17048
rect 4198 17014 4217 17048
rect 3967 16939 4001 16973
rect 4039 16940 4073 16974
rect 4111 16941 4145 16975
rect 4183 16941 4198 16975
rect 4198 16941 4217 16975
rect 3967 16866 4001 16900
rect 4039 16867 4073 16901
rect 4111 16868 4145 16902
rect 4183 16868 4198 16902
rect 4198 16868 4217 16902
rect 3967 16793 4001 16827
rect 4039 16794 4073 16828
rect 4111 16795 4145 16829
rect 4183 16795 4198 16829
rect 4198 16795 4217 16829
rect 3967 16720 4001 16754
rect 4039 16721 4073 16755
rect 4111 16722 4145 16756
rect 4183 16722 4198 16756
rect 4198 16722 4217 16756
rect 3967 16647 4001 16681
rect 4039 16648 4073 16682
rect 4111 16649 4145 16683
rect 4183 16649 4198 16683
rect 4198 16649 4217 16683
rect 3967 16574 4001 16608
rect 4039 16575 4073 16609
rect 4111 16576 4145 16610
rect 4183 16576 4198 16610
rect 4198 16576 4217 16610
rect 3967 16501 4001 16535
rect 4039 16502 4073 16536
rect 4111 16503 4145 16537
rect 4183 16503 4198 16537
rect 4198 16503 4217 16537
rect 3967 16428 4001 16462
rect 4039 16429 4073 16463
rect 4111 16430 4145 16464
rect 4183 16430 4198 16464
rect 4198 16430 4217 16464
rect 3967 16355 4001 16389
rect 4039 16356 4073 16390
rect 4111 16357 4145 16391
rect 4183 16357 4198 16391
rect 4198 16357 4217 16391
rect 3967 16282 4001 16316
rect 4039 16283 4073 16317
rect 4111 16284 4145 16318
rect 4183 16284 4198 16318
rect 4198 16284 4217 16318
rect 3967 16209 4001 16243
rect 4039 16210 4073 16244
rect 4111 16211 4145 16245
rect 4183 16211 4198 16245
rect 4198 16211 4217 16245
rect 3967 16136 4001 16170
rect 4039 16137 4073 16171
rect 4111 16138 4145 16172
rect 4183 16138 4198 16172
rect 4198 16138 4217 16172
rect 3967 16063 4001 16097
rect 4039 16064 4073 16098
rect 4111 16065 4145 16099
rect 4183 16065 4198 16099
rect 4198 16065 4217 16099
rect 3967 15990 4001 16024
rect 4039 15991 4073 16025
rect 4111 15992 4145 16026
rect 4183 15992 4198 16026
rect 4198 15992 4217 16026
rect 3967 15917 4001 15951
rect 4039 15918 4073 15952
rect 4111 15919 4145 15953
rect 4183 15919 4198 15953
rect 4198 15919 4217 15953
rect 3967 15844 4001 15878
rect 4039 15845 4073 15879
rect 4111 15846 4145 15880
rect 4183 15846 4198 15880
rect 4198 15846 4217 15880
rect 3967 15771 4001 15805
rect 4039 15772 4073 15806
rect 4111 15773 4145 15807
rect 4183 15773 4198 15807
rect 4198 15773 4217 15807
rect 3967 15698 4001 15732
rect 4039 15699 4073 15733
rect 4111 15700 4145 15734
rect 4183 15700 4198 15734
rect 4198 15700 4217 15734
rect 3967 15625 4001 15659
rect 4039 15626 4073 15660
rect 4111 15627 4145 15661
rect 4183 15627 4198 15661
rect 4198 15627 4217 15661
rect 3967 15552 4001 15586
rect 4039 15553 4073 15587
rect 4111 15554 4145 15588
rect 4183 15554 4198 15588
rect 4198 15554 4217 15588
rect 3967 15479 4001 15513
rect 4039 15480 4073 15514
rect 4111 15481 4145 15515
rect 4183 15481 4198 15515
rect 4198 15481 4217 15515
rect 3967 15406 4001 15440
rect 4039 15407 4073 15441
rect 4111 15408 4145 15442
rect 4183 15408 4198 15442
rect 4198 15408 4217 15442
rect 3967 15333 4001 15367
rect 4039 15334 4073 15368
rect 4111 15335 4145 15369
rect 4183 15335 4198 15369
rect 4198 15335 4217 15369
rect 3967 15260 4001 15294
rect 4039 15261 4073 15295
rect 4111 15262 4145 15296
rect 4183 15262 4198 15296
rect 4198 15262 4217 15296
rect 3967 15187 4001 15221
rect 4039 15188 4073 15222
rect 4111 15189 4145 15223
rect 4183 15189 4198 15223
rect 4198 15189 4217 15223
rect 3967 15114 4001 15148
rect 4039 15115 4073 15149
rect 4111 15116 4145 15150
rect 4183 15116 4198 15150
rect 4198 15116 4217 15150
rect 3967 15041 4001 15075
rect 4039 15042 4073 15076
rect 4111 15043 4145 15077
rect 4183 15043 4198 15077
rect 4198 15043 4217 15077
rect 3967 14968 4001 15002
rect 4039 14969 4073 15003
rect 4111 14970 4145 15004
rect 4183 14970 4198 15004
rect 4198 14970 4217 15004
rect 3967 14895 4001 14929
rect 4039 14896 4073 14930
rect 4111 14897 4145 14931
rect 4183 14897 4198 14931
rect 4198 14897 4217 14931
rect 1881 14836 1915 14870
rect 1953 14836 1987 14870
rect 3694 14840 3728 14874
rect 3766 14840 3800 14874
rect 3967 14822 4001 14856
rect 4039 14823 4073 14857
rect 4111 14824 4145 14858
rect 4183 14824 4198 14858
rect 4198 14824 4217 14858
rect 3967 14749 4001 14783
rect 4039 14750 4073 14784
rect 4111 14751 4145 14785
rect 4183 14751 4198 14785
rect 4198 14751 4217 14785
rect 3967 14676 4001 14710
rect 4039 14677 4073 14711
rect 4111 14678 4145 14712
rect 4183 14678 4198 14712
rect 4198 14678 4217 14712
rect 3967 14634 4001 14637
rect 3967 14603 4001 14634
rect 4039 14604 4073 14638
rect 4111 14605 4145 14639
rect 4183 14605 4198 14639
rect 4198 14605 4217 14639
rect 1899 14562 1933 14564
rect 1973 14562 2007 14564
rect 2047 14562 2081 14564
rect 2121 14562 2155 14564
rect 2195 14562 2229 14564
rect 2269 14562 2303 14564
rect 2343 14562 2377 14564
rect 2417 14562 2451 14564
rect 2491 14562 2525 14564
rect 2565 14562 2599 14564
rect 2639 14562 2673 14564
rect 2713 14562 2747 14564
rect 2787 14562 2821 14564
rect 2861 14562 2895 14564
rect 2935 14562 2969 14564
rect 3009 14562 3043 14564
rect 3083 14562 3117 14564
rect 3157 14562 3191 14564
rect 3231 14562 3265 14564
rect 3305 14562 3339 14564
rect 3379 14562 3413 14564
rect 3453 14562 3487 14564
rect 3527 14562 3561 14564
rect 3601 14562 3635 14564
rect 3675 14562 3709 14564
rect 3748 14562 3782 14564
rect 3821 14562 3855 14564
rect 3894 14562 3928 14564
rect 3967 14562 4001 14564
rect 1899 14530 1920 14562
rect 1920 14530 1933 14562
rect 1973 14530 1988 14562
rect 1988 14530 2007 14562
rect 2047 14530 2081 14562
rect 2121 14530 2155 14562
rect 2195 14530 2229 14562
rect 2269 14530 2303 14562
rect 2343 14530 2377 14562
rect 2417 14530 2451 14562
rect 2491 14530 2525 14562
rect 2565 14530 2599 14562
rect 2639 14530 2673 14562
rect 2713 14530 2747 14562
rect 2787 14530 2821 14562
rect 2861 14530 2895 14562
rect 2935 14530 2969 14562
rect 3009 14530 3043 14562
rect 3083 14530 3117 14562
rect 3157 14530 3191 14562
rect 3231 14530 3265 14562
rect 3305 14530 3339 14562
rect 3379 14530 3413 14562
rect 3453 14530 3487 14562
rect 3527 14530 3561 14562
rect 3601 14530 3635 14562
rect 3675 14530 3709 14562
rect 3748 14530 3782 14562
rect 3821 14530 3855 14562
rect 3894 14530 3928 14562
rect 3967 14530 3994 14562
rect 3994 14530 4001 14562
rect 4039 14531 4073 14565
rect 4111 14532 4145 14566
rect 4183 14532 4198 14566
rect 4198 14532 4217 14566
rect 1827 13882 1834 14492
rect 1834 14420 1933 14492
rect 1973 14460 1988 14492
rect 1988 14460 2007 14492
rect 2047 14460 2081 14492
rect 1973 14458 2007 14460
rect 2047 14458 2056 14460
rect 2056 14458 2081 14460
rect 2121 14458 2155 14492
rect 2195 14458 2229 14492
rect 2269 14458 2303 14492
rect 2343 14458 2377 14492
rect 2417 14458 2451 14492
rect 2491 14458 2525 14492
rect 2565 14458 2599 14492
rect 2639 14458 2673 14492
rect 2713 14458 2747 14492
rect 2787 14458 2821 14492
rect 2861 14458 2895 14492
rect 2935 14458 2969 14492
rect 3009 14458 3043 14492
rect 3083 14458 3117 14492
rect 3157 14458 3191 14492
rect 3231 14458 3265 14492
rect 3305 14458 3339 14492
rect 3379 14458 3413 14492
rect 3453 14458 3487 14492
rect 3527 14458 3561 14492
rect 3601 14458 3635 14492
rect 3674 14458 3708 14492
rect 3747 14458 3781 14492
rect 3820 14458 3854 14492
rect 3893 14458 3927 14492
rect 3966 14458 4000 14492
rect 4039 14458 4062 14492
rect 4062 14458 4073 14492
rect 4111 14459 4145 14493
rect 4183 14464 4217 14493
rect 4183 14459 4198 14464
rect 4198 14459 4217 14464
rect 1834 14358 2004 14420
rect 2004 14358 2005 14420
rect 2045 14392 2056 14420
rect 2056 14392 2079 14420
rect 2119 14392 2153 14420
rect 2045 14386 2079 14392
rect 2119 14386 2124 14392
rect 2124 14386 2153 14392
rect 2193 14386 2227 14420
rect 2267 14386 2301 14420
rect 2341 14386 2375 14420
rect 2415 14386 2449 14420
rect 2489 14386 2523 14420
rect 2563 14386 2597 14420
rect 2637 14386 2671 14420
rect 2711 14386 2745 14420
rect 2785 14386 2819 14420
rect 2859 14386 2893 14420
rect 2933 14386 2967 14420
rect 3007 14386 3041 14420
rect 3081 14386 3115 14420
rect 3155 14386 3189 14420
rect 3229 14386 3263 14420
rect 3303 14386 3337 14420
rect 3377 14386 3411 14420
rect 3451 14386 3485 14420
rect 3525 14386 3559 14420
rect 3599 14386 3633 14420
rect 3672 14386 3706 14420
rect 3745 14386 3779 14420
rect 3818 14386 3852 14420
rect 3891 14386 3925 14420
rect 3964 14386 3998 14420
rect 4037 14386 4071 14420
rect 4111 14386 4130 14420
rect 4130 14386 4145 14420
rect 4183 14386 4217 14420
rect 1834 14348 2005 14358
rect 1834 13882 2072 14348
rect 2072 13882 2077 14348
rect 2117 14324 2124 14348
rect 2124 14324 2151 14348
rect 2191 14324 2225 14348
rect 2265 14324 2299 14348
rect 2339 14324 2373 14348
rect 2413 14324 2447 14348
rect 2487 14324 2521 14348
rect 2561 14324 2595 14348
rect 2635 14324 2669 14348
rect 2709 14324 2743 14348
rect 2783 14324 2817 14348
rect 2857 14324 2891 14348
rect 2931 14324 2965 14348
rect 3005 14324 3039 14348
rect 3079 14324 3113 14348
rect 3153 14324 3187 14348
rect 3227 14324 3261 14348
rect 3301 14324 3335 14348
rect 3375 14324 3409 14348
rect 3449 14324 3483 14348
rect 3523 14324 3557 14348
rect 3597 14324 3631 14348
rect 3671 14324 3705 14348
rect 3745 14324 3779 14348
rect 3818 14324 3852 14348
rect 3891 14324 3925 14348
rect 3964 14324 3998 14348
rect 4037 14324 4071 14348
rect 4110 14324 4130 14348
rect 4130 14324 4144 14348
rect 2117 14314 2151 14324
rect 2191 14314 2225 14324
rect 2265 14314 2299 14324
rect 2339 14314 2373 14324
rect 2413 14314 2447 14324
rect 2487 14314 2521 14324
rect 2561 14314 2595 14324
rect 2635 14314 2669 14324
rect 2709 14314 2743 14324
rect 2783 14314 2817 14324
rect 2857 14314 2891 14324
rect 2931 14314 2965 14324
rect 3005 14314 3039 14324
rect 3079 14314 3113 14324
rect 3153 14314 3187 14324
rect 3227 14314 3261 14324
rect 3301 14314 3335 14324
rect 3375 14314 3409 14324
rect 3449 14314 3483 14324
rect 3523 14314 3557 14324
rect 3597 14314 3631 14324
rect 3671 14314 3705 14324
rect 3745 14314 3779 14324
rect 3818 14314 3852 14324
rect 3891 14314 3925 14324
rect 3964 14314 3998 14324
rect 4037 14314 4071 14324
rect 4110 14314 4144 14324
rect 4358 18592 4362 19490
rect 4362 18592 4532 19490
rect 4358 18519 4362 18553
rect 4362 18519 4392 18553
rect 4430 18520 4532 18592
rect 4532 18520 4536 19490
rect 4784 18922 4890 22484
rect 4784 18849 4818 18883
rect 4856 18849 4890 18883
rect 4784 18776 4818 18810
rect 4856 18776 4890 18810
rect 4784 18703 4818 18737
rect 4856 18703 4890 18737
rect 5637 20017 5815 22571
rect 5637 19944 5671 19978
rect 5709 19944 5743 19978
rect 5781 19944 5815 19978
rect 5637 19871 5671 19905
rect 5709 19871 5743 19905
rect 5781 19871 5815 19905
rect 5637 19798 5671 19832
rect 5709 19798 5743 19832
rect 5781 19798 5815 19832
rect 5637 19725 5671 19759
rect 5709 19725 5743 19759
rect 5781 19725 5815 19759
rect 5637 19652 5671 19686
rect 5709 19652 5743 19686
rect 5781 19652 5815 19686
rect 5637 19579 5671 19613
rect 5709 19579 5743 19613
rect 5781 19579 5815 19613
rect 5637 19506 5671 19540
rect 5709 19506 5743 19540
rect 5781 19506 5815 19540
rect 5637 19433 5671 19467
rect 5709 19433 5743 19467
rect 5781 19433 5815 19467
rect 5637 19360 5671 19394
rect 5709 19360 5743 19394
rect 5781 19360 5815 19394
rect 5637 19287 5671 19321
rect 5709 19287 5743 19321
rect 5781 19287 5815 19321
rect 5637 19214 5671 19248
rect 5709 19214 5743 19248
rect 5781 19214 5815 19248
rect 5637 19141 5671 19175
rect 5709 19141 5743 19175
rect 5781 19141 5815 19175
rect 5637 19068 5671 19102
rect 5709 19068 5743 19102
rect 5781 19068 5815 19102
rect 5637 18995 5671 19029
rect 5709 18995 5743 19029
rect 5781 18995 5815 19029
rect 5637 18922 5671 18956
rect 5709 18922 5743 18956
rect 5781 18922 5815 18956
rect 5637 18849 5671 18883
rect 5709 18849 5743 18883
rect 5781 18849 5815 18883
rect 5637 18776 5671 18810
rect 5709 18776 5743 18810
rect 5781 18776 5815 18810
rect 5637 18703 5671 18737
rect 5709 18703 5743 18737
rect 5781 18703 5815 18737
rect 6557 19360 6735 22562
rect 6557 19287 6591 19321
rect 6629 19287 6663 19321
rect 6701 19287 6735 19321
rect 6557 19214 6591 19248
rect 6629 19214 6663 19248
rect 6701 19214 6735 19248
rect 6557 19141 6591 19175
rect 6629 19141 6663 19175
rect 6701 19141 6735 19175
rect 6557 19068 6591 19102
rect 6629 19068 6663 19102
rect 6701 19068 6735 19102
rect 6557 18995 6591 19029
rect 6629 18995 6663 19029
rect 6701 18995 6735 19029
rect 6557 18922 6591 18956
rect 6629 18922 6663 18956
rect 6701 18922 6735 18956
rect 6557 18849 6591 18883
rect 6629 18849 6663 18883
rect 6701 18849 6735 18883
rect 6557 18776 6591 18810
rect 6629 18776 6663 18810
rect 6701 18776 6735 18810
rect 6557 18703 6591 18737
rect 6629 18703 6663 18737
rect 6701 18703 6735 18737
rect 7477 19360 7655 22562
rect 7477 19287 7511 19321
rect 7549 19287 7583 19321
rect 7621 19287 7655 19321
rect 7477 19214 7511 19248
rect 7549 19214 7583 19248
rect 7621 19214 7655 19248
rect 7477 19141 7511 19175
rect 7549 19141 7583 19175
rect 7621 19141 7655 19175
rect 7477 19068 7511 19102
rect 7549 19068 7583 19102
rect 7621 19068 7655 19102
rect 7477 18995 7511 19029
rect 7549 18995 7583 19029
rect 7621 18995 7655 19029
rect 7477 18922 7511 18956
rect 7549 18922 7583 18956
rect 7621 18922 7655 18956
rect 7477 18849 7511 18883
rect 7549 18849 7583 18883
rect 7621 18849 7655 18883
rect 7477 18776 7511 18810
rect 7549 18776 7583 18810
rect 7621 18776 7655 18810
rect 7477 18703 7511 18737
rect 7549 18703 7583 18737
rect 7621 18703 7655 18737
rect 8397 19360 8575 22562
rect 8397 19287 8431 19321
rect 8469 19287 8503 19321
rect 8541 19287 8575 19321
rect 8397 19214 8431 19248
rect 8469 19214 8503 19248
rect 8541 19214 8575 19248
rect 8397 19141 8431 19175
rect 8469 19141 8503 19175
rect 8541 19141 8575 19175
rect 8397 19068 8431 19102
rect 8469 19068 8503 19102
rect 8541 19068 8575 19102
rect 8397 18995 8431 19029
rect 8469 18995 8503 19029
rect 8541 18995 8575 19029
rect 8397 18922 8431 18956
rect 8469 18922 8503 18956
rect 8541 18922 8575 18956
rect 8397 18849 8431 18883
rect 8469 18849 8503 18883
rect 8541 18849 8575 18883
rect 8397 18776 8431 18810
rect 8469 18776 8503 18810
rect 8541 18776 8575 18810
rect 8397 18703 8431 18737
rect 8469 18703 8503 18737
rect 8541 18703 8575 18737
rect 9317 19360 9495 22562
rect 9317 19287 9351 19321
rect 9389 19287 9423 19321
rect 9461 19287 9495 19321
rect 9317 19214 9351 19248
rect 9389 19214 9423 19248
rect 9461 19214 9495 19248
rect 9317 19141 9351 19175
rect 9389 19141 9423 19175
rect 9461 19141 9495 19175
rect 9317 19068 9351 19102
rect 9389 19068 9423 19102
rect 9461 19068 9495 19102
rect 9317 18995 9351 19029
rect 9389 18995 9423 19029
rect 9461 18995 9495 19029
rect 9317 18922 9351 18956
rect 9389 18922 9423 18956
rect 9461 18922 9495 18956
rect 9317 18849 9351 18883
rect 9389 18849 9423 18883
rect 9461 18849 9495 18883
rect 9317 18776 9351 18810
rect 9389 18776 9423 18810
rect 9461 18776 9495 18810
rect 9317 18703 9351 18737
rect 9389 18703 9423 18737
rect 9461 18703 9495 18737
rect 10237 19360 10415 22562
rect 10237 19287 10271 19321
rect 10309 19287 10343 19321
rect 10381 19287 10415 19321
rect 10237 19214 10271 19248
rect 10309 19214 10343 19248
rect 10381 19214 10415 19248
rect 10237 19141 10271 19175
rect 10309 19141 10343 19175
rect 10381 19141 10415 19175
rect 10237 19068 10271 19102
rect 10309 19068 10343 19102
rect 10381 19068 10415 19102
rect 10237 18995 10271 19029
rect 10309 18995 10343 19029
rect 10381 18995 10415 19029
rect 10237 18922 10271 18956
rect 10309 18922 10343 18956
rect 10381 18922 10415 18956
rect 10237 18849 10271 18883
rect 10309 18849 10343 18883
rect 10381 18849 10415 18883
rect 10237 18776 10271 18810
rect 10309 18776 10343 18810
rect 10381 18776 10415 18810
rect 10237 18703 10271 18737
rect 10309 18703 10343 18737
rect 10381 18703 10415 18737
rect 11157 19360 11335 22562
rect 11157 19287 11191 19321
rect 11229 19287 11263 19321
rect 11301 19287 11335 19321
rect 11157 19214 11191 19248
rect 11229 19214 11263 19248
rect 11301 19214 11335 19248
rect 11157 19141 11191 19175
rect 11229 19141 11263 19175
rect 11301 19141 11335 19175
rect 11157 19068 11191 19102
rect 11229 19068 11263 19102
rect 11301 19068 11335 19102
rect 11157 18995 11191 19029
rect 11229 18995 11263 19029
rect 11301 18995 11335 19029
rect 11157 18922 11191 18956
rect 11229 18922 11263 18956
rect 11301 18922 11335 18956
rect 11157 18849 11191 18883
rect 11229 18849 11263 18883
rect 11301 18849 11335 18883
rect 11157 18776 11191 18810
rect 11229 18776 11263 18810
rect 11301 18776 11335 18810
rect 11157 18703 11191 18737
rect 11229 18703 11263 18737
rect 11301 18703 11335 18737
rect 12077 19360 12255 22562
rect 12077 19287 12111 19321
rect 12149 19287 12183 19321
rect 12221 19287 12255 19321
rect 12077 19214 12111 19248
rect 12149 19214 12183 19248
rect 12221 19214 12255 19248
rect 12997 19360 13175 22562
rect 13507 22532 13541 22566
rect 13597 22532 13628 22566
rect 13628 22532 13631 22566
rect 13507 22459 13541 22493
rect 13597 22459 13628 22493
rect 13628 22459 13631 22493
rect 13507 22386 13541 22420
rect 13597 22386 13628 22420
rect 13628 22386 13631 22420
rect 13507 22313 13541 22347
rect 13597 22313 13628 22347
rect 13628 22313 13631 22347
rect 13507 22240 13541 22274
rect 13597 22240 13628 22274
rect 13628 22240 13631 22274
rect 13507 22167 13541 22201
rect 13597 22167 13628 22201
rect 13628 22167 13631 22201
rect 13507 22094 13541 22128
rect 13597 22094 13628 22128
rect 13628 22094 13631 22128
rect 13507 22021 13541 22055
rect 13597 22021 13628 22055
rect 13628 22021 13631 22055
rect 13507 21948 13541 21982
rect 13597 21948 13628 21982
rect 13628 21948 13631 21982
rect 13507 21875 13541 21909
rect 13597 21875 13628 21909
rect 13628 21875 13631 21909
rect 13507 21802 13541 21836
rect 13597 21802 13628 21836
rect 13628 21802 13631 21836
rect 13507 21729 13541 21763
rect 13597 21729 13628 21763
rect 13628 21729 13631 21763
rect 13507 21656 13541 21690
rect 13597 21656 13628 21690
rect 13628 21656 13631 21690
rect 13507 21583 13541 21617
rect 13597 21583 13628 21617
rect 13628 21583 13631 21617
rect 13507 21510 13541 21544
rect 13597 21510 13628 21544
rect 13628 21510 13631 21544
rect 13507 21437 13541 21471
rect 13597 21437 13628 21471
rect 13628 21437 13631 21471
rect 13507 21364 13541 21398
rect 13597 21364 13628 21398
rect 13628 21364 13631 21398
rect 13507 21291 13541 21325
rect 13597 21291 13628 21325
rect 13628 21291 13631 21325
rect 13507 21218 13541 21252
rect 13597 21218 13628 21252
rect 13628 21218 13631 21252
rect 13507 21145 13541 21179
rect 13597 21145 13628 21179
rect 13628 21145 13631 21179
rect 13507 21072 13541 21106
rect 13597 21072 13628 21106
rect 13628 21072 13631 21106
rect 13507 20999 13541 21033
rect 13597 20999 13628 21033
rect 13628 20999 13631 21033
rect 13507 20926 13541 20960
rect 13597 20926 13628 20960
rect 13628 20926 13631 20960
rect 13507 20853 13541 20887
rect 13597 20853 13628 20887
rect 13628 20853 13631 20887
rect 13507 20780 13541 20814
rect 13597 20780 13628 20814
rect 13628 20780 13631 20814
rect 13507 20707 13541 20741
rect 13597 20707 13628 20741
rect 13628 20707 13631 20741
rect 13507 20634 13541 20668
rect 13597 20634 13628 20668
rect 13628 20634 13631 20668
rect 13507 20561 13541 20595
rect 13597 20561 13628 20595
rect 13628 20561 13631 20595
rect 13507 20488 13541 20522
rect 13597 20488 13628 20522
rect 13628 20488 13631 20522
rect 13507 20415 13541 20449
rect 13597 20415 13628 20449
rect 13628 20415 13631 20449
rect 13507 20342 13541 20376
rect 13597 20342 13628 20376
rect 13628 20342 13631 20376
rect 13775 32712 13781 34978
rect 13781 32712 14019 34978
rect 14019 32712 14025 35122
rect 13775 32623 13781 32657
rect 13781 32623 13809 32657
rect 13847 32623 13881 32657
rect 13919 32623 13953 32657
rect 13991 32623 14019 32657
rect 14019 32623 14025 32657
rect 13775 32550 13781 32584
rect 13781 32550 13809 32584
rect 13847 32550 13881 32584
rect 13919 32550 13953 32584
rect 13991 32550 14019 32584
rect 14019 32550 14025 32584
rect 13775 32477 13781 32511
rect 13781 32477 13809 32511
rect 13847 32477 13881 32511
rect 13919 32477 13953 32511
rect 13991 32477 14019 32511
rect 14019 32477 14025 32511
rect 13775 32404 13781 32438
rect 13781 32404 13809 32438
rect 13847 32404 13881 32438
rect 13919 32404 13953 32438
rect 13991 32404 14019 32438
rect 14019 32404 14025 32438
rect 13775 32331 13781 32365
rect 13781 32331 13809 32365
rect 13847 32331 13881 32365
rect 13919 32331 13953 32365
rect 13991 32331 14019 32365
rect 14019 32331 14025 32365
rect 13775 32258 13781 32292
rect 13781 32258 13809 32292
rect 13847 32258 13881 32292
rect 13919 32258 13953 32292
rect 13991 32258 14019 32292
rect 14019 32258 14025 32292
rect 13775 32185 13781 32219
rect 13781 32185 13809 32219
rect 13847 32185 13881 32219
rect 13919 32185 13953 32219
rect 13991 32185 14019 32219
rect 14019 32185 14025 32219
rect 13775 32112 13781 32146
rect 13781 32112 13809 32146
rect 13847 32112 13881 32146
rect 13919 32112 13953 32146
rect 13991 32112 14019 32146
rect 14019 32112 14025 32146
rect 13775 32039 13781 32073
rect 13781 32039 13809 32073
rect 13847 32039 13881 32073
rect 13919 32039 13953 32073
rect 13991 32039 14019 32073
rect 14019 32039 14025 32073
rect 13775 31966 13781 32000
rect 13781 31966 13809 32000
rect 13847 31966 13881 32000
rect 13919 31966 13953 32000
rect 13991 31966 14019 32000
rect 14019 31966 14025 32000
rect 13775 31893 13781 31927
rect 13781 31893 13809 31927
rect 13847 31893 13881 31927
rect 13919 31893 13953 31927
rect 13991 31893 14019 31927
rect 14019 31893 14025 31927
rect 13775 31820 13781 31854
rect 13781 31820 13809 31854
rect 13847 31820 13881 31854
rect 13919 31820 13953 31854
rect 13991 31820 14019 31854
rect 14019 31820 14025 31854
rect 13775 31747 13781 31781
rect 13781 31747 13809 31781
rect 13847 31747 13881 31781
rect 13919 31747 13953 31781
rect 13991 31747 14019 31781
rect 14019 31747 14025 31781
rect 13775 31674 13781 31708
rect 13781 31674 13809 31708
rect 13847 31674 13881 31708
rect 13919 31674 13953 31708
rect 13991 31674 14019 31708
rect 14019 31674 14025 31708
rect 13775 31601 13781 31635
rect 13781 31601 13809 31635
rect 13847 31601 13881 31635
rect 13919 31601 13953 31635
rect 13991 31601 14019 31635
rect 14019 31601 14025 31635
rect 13775 31528 13781 31562
rect 13781 31528 13809 31562
rect 13847 31528 13881 31562
rect 13919 31528 13953 31562
rect 13991 31528 14019 31562
rect 14019 31528 14025 31562
rect 13775 31455 13781 31489
rect 13781 31455 13809 31489
rect 13847 31455 13881 31489
rect 13919 31455 13953 31489
rect 13991 31455 14019 31489
rect 14019 31455 14025 31489
rect 13775 31382 13781 31416
rect 13781 31382 13809 31416
rect 13847 31382 13881 31416
rect 13919 31382 13953 31416
rect 13991 31382 14019 31416
rect 14019 31382 14025 31416
rect 13775 31309 13781 31343
rect 13781 31309 13809 31343
rect 13847 31309 13881 31343
rect 13919 31309 13953 31343
rect 13991 31309 14019 31343
rect 14019 31309 14025 31343
rect 13775 31236 13781 31270
rect 13781 31236 13809 31270
rect 13847 31236 13881 31270
rect 13919 31236 13953 31270
rect 13991 31236 14019 31270
rect 14019 31236 14025 31270
rect 13775 31163 13781 31197
rect 13781 31163 13809 31197
rect 13847 31163 13881 31197
rect 13919 31163 13953 31197
rect 13991 31163 14019 31197
rect 14019 31163 14025 31197
rect 13775 31090 13781 31124
rect 13781 31090 13809 31124
rect 13847 31090 13881 31124
rect 13919 31090 13953 31124
rect 13991 31090 14019 31124
rect 14019 31090 14025 31124
rect 13775 31017 13781 31051
rect 13781 31017 13809 31051
rect 13847 31017 13881 31051
rect 13919 31017 13953 31051
rect 13991 31017 14019 31051
rect 14019 31017 14025 31051
rect 13775 30944 13781 30978
rect 13781 30944 13809 30978
rect 13847 30944 13881 30978
rect 13919 30944 13953 30978
rect 13991 30944 14019 30978
rect 14019 30944 14025 30978
rect 13775 30871 13781 30905
rect 13781 30871 13809 30905
rect 13847 30871 13881 30905
rect 13919 30871 13953 30905
rect 13991 30871 14019 30905
rect 14019 30871 14025 30905
rect 13775 30798 13781 30832
rect 13781 30798 13809 30832
rect 13847 30798 13881 30832
rect 13919 30798 13953 30832
rect 13991 30798 14019 30832
rect 14019 30798 14025 30832
rect 13775 30725 13781 30759
rect 13781 30725 13809 30759
rect 13847 30725 13881 30759
rect 13919 30725 13953 30759
rect 13991 30725 14019 30759
rect 14019 30725 14025 30759
rect 13775 30652 13781 30686
rect 13781 30652 13809 30686
rect 13847 30652 13881 30686
rect 13919 30652 13953 30686
rect 13991 30652 14019 30686
rect 14019 30652 14025 30686
rect 13775 30579 13781 30613
rect 13781 30579 13809 30613
rect 13847 30579 13881 30613
rect 13919 30579 13953 30613
rect 13991 30579 14019 30613
rect 14019 30579 14025 30613
rect 13775 30506 13781 30540
rect 13781 30506 13809 30540
rect 13847 30506 13881 30540
rect 13919 30506 13953 30540
rect 13991 30506 14019 30540
rect 14019 30506 14025 30540
rect 13775 30433 13781 30467
rect 13781 30433 13809 30467
rect 13847 30433 13881 30467
rect 13919 30433 13953 30467
rect 13991 30433 14019 30467
rect 14019 30433 14025 30467
rect 13775 30360 13781 30394
rect 13781 30360 13809 30394
rect 13847 30360 13881 30394
rect 13919 30360 13953 30394
rect 13991 30360 14019 30394
rect 14019 30360 14025 30394
rect 13775 30287 13781 30321
rect 13781 30287 13809 30321
rect 13847 30287 13881 30321
rect 13919 30287 13953 30321
rect 13991 30287 14019 30321
rect 14019 30287 14025 30321
rect 13775 30214 13781 30248
rect 13781 30214 13809 30248
rect 13847 30214 13881 30248
rect 13919 30214 13953 30248
rect 13991 30214 14019 30248
rect 14019 30214 14025 30248
rect 13775 30141 13781 30175
rect 13781 30141 13809 30175
rect 13847 30141 13881 30175
rect 13919 30141 13953 30175
rect 13991 30141 14019 30175
rect 14019 30141 14025 30175
rect 13775 30068 13781 30102
rect 13781 30068 13809 30102
rect 13847 30068 13881 30102
rect 13919 30068 13953 30102
rect 13991 30068 14019 30102
rect 14019 30068 14025 30102
rect 13775 29995 13781 30029
rect 13781 29995 13809 30029
rect 13847 29995 13881 30029
rect 13919 29995 13953 30029
rect 13991 29995 14019 30029
rect 14019 29995 14025 30029
rect 13775 29922 13781 29956
rect 13781 29922 13809 29956
rect 13847 29922 13881 29956
rect 13919 29922 13953 29956
rect 13991 29922 14019 29956
rect 14019 29922 14025 29956
rect 13775 29849 13781 29883
rect 13781 29849 13809 29883
rect 13847 29849 13881 29883
rect 13919 29849 13953 29883
rect 13991 29849 14019 29883
rect 14019 29849 14025 29883
rect 13775 29776 13781 29810
rect 13781 29776 13809 29810
rect 13847 29776 13881 29810
rect 13919 29776 13953 29810
rect 13991 29776 14019 29810
rect 14019 29776 14025 29810
rect 13775 29703 13781 29737
rect 13781 29703 13809 29737
rect 13847 29703 13881 29737
rect 13919 29703 13953 29737
rect 13991 29703 14019 29737
rect 14019 29703 14025 29737
rect 13775 29630 13781 29664
rect 13781 29630 13809 29664
rect 13847 29630 13881 29664
rect 13919 29630 13953 29664
rect 13991 29630 14019 29664
rect 14019 29630 14025 29664
rect 13775 29557 13781 29591
rect 13781 29557 13809 29591
rect 13847 29557 13881 29591
rect 13919 29557 13953 29591
rect 13991 29557 14019 29591
rect 14019 29557 14025 29591
rect 13775 29484 13781 29518
rect 13781 29484 13809 29518
rect 13847 29484 13881 29518
rect 13919 29484 13953 29518
rect 13991 29484 14019 29518
rect 14019 29484 14025 29518
rect 13775 29411 13781 29445
rect 13781 29411 13809 29445
rect 13847 29411 13881 29445
rect 13919 29411 13953 29445
rect 13991 29411 14019 29445
rect 14019 29411 14025 29445
rect 13775 29338 13781 29372
rect 13781 29338 13809 29372
rect 13847 29338 13881 29372
rect 13919 29338 13953 29372
rect 13991 29338 14019 29372
rect 14019 29338 14025 29372
rect 13775 29265 13781 29299
rect 13781 29265 13809 29299
rect 13847 29265 13881 29299
rect 13919 29265 13953 29299
rect 13991 29265 14019 29299
rect 14019 29265 14025 29299
rect 13775 29192 13781 29226
rect 13781 29192 13809 29226
rect 13847 29192 13881 29226
rect 13919 29192 13953 29226
rect 13991 29192 14019 29226
rect 14019 29192 14025 29226
rect 13775 29119 13781 29153
rect 13781 29119 13809 29153
rect 13847 29119 13881 29153
rect 13919 29119 13953 29153
rect 13991 29119 14019 29153
rect 14019 29119 14025 29153
rect 13775 29046 13781 29080
rect 13781 29046 13809 29080
rect 13847 29046 13881 29080
rect 13919 29046 13953 29080
rect 13991 29046 14019 29080
rect 14019 29046 14025 29080
rect 13775 28973 13781 29007
rect 13781 28973 13809 29007
rect 13847 28973 13881 29007
rect 13919 28973 13953 29007
rect 13991 28973 14019 29007
rect 14019 28973 14025 29007
rect 13775 28900 13781 28934
rect 13781 28900 13809 28934
rect 13847 28900 13881 28934
rect 13919 28900 13953 28934
rect 13991 28900 14019 28934
rect 14019 28900 14025 28934
rect 13775 28827 13781 28861
rect 13781 28827 13809 28861
rect 13847 28827 13881 28861
rect 13919 28827 13953 28861
rect 13991 28827 14019 28861
rect 14019 28827 14025 28861
rect 13775 28754 13781 28788
rect 13781 28754 13809 28788
rect 13847 28754 13881 28788
rect 13919 28754 13953 28788
rect 13991 28754 14019 28788
rect 14019 28754 14025 28788
rect 13775 28681 13781 28715
rect 13781 28681 13809 28715
rect 13847 28681 13881 28715
rect 13919 28681 13953 28715
rect 13991 28681 14019 28715
rect 14019 28681 14025 28715
rect 13775 28608 13781 28642
rect 13781 28608 13809 28642
rect 13847 28608 13881 28642
rect 13919 28608 13953 28642
rect 13991 28608 14019 28642
rect 14019 28608 14025 28642
rect 13775 28535 13781 28569
rect 13781 28535 13809 28569
rect 13847 28535 13881 28569
rect 13919 28535 13953 28569
rect 13991 28535 14019 28569
rect 14019 28535 14025 28569
rect 13775 28462 13781 28496
rect 13781 28462 13809 28496
rect 13847 28462 13881 28496
rect 13919 28462 13953 28496
rect 13991 28462 14019 28496
rect 14019 28462 14025 28496
rect 12997 19287 13031 19321
rect 13069 19287 13103 19321
rect 13141 19287 13175 19321
rect 12997 19214 13031 19248
rect 13069 19214 13103 19248
rect 13141 19214 13175 19248
rect 12077 19141 12111 19175
rect 12149 19141 12183 19175
rect 12221 19141 12255 19175
rect 12077 19068 12111 19102
rect 12149 19068 12183 19102
rect 12221 19068 12255 19102
rect 12077 18995 12111 19029
rect 12149 18995 12183 19029
rect 12221 18995 12255 19029
rect 12077 18922 12111 18956
rect 12149 18922 12183 18956
rect 12221 18922 12255 18956
rect 12077 18849 12111 18883
rect 12149 18849 12183 18883
rect 12221 18849 12255 18883
rect 12077 18776 12111 18810
rect 12149 18776 12183 18810
rect 12221 18776 12255 18810
rect 12077 18703 12111 18737
rect 12149 18703 12183 18737
rect 12221 18703 12255 18737
rect 12997 19141 13031 19175
rect 13069 19141 13103 19175
rect 13141 19141 13175 19175
rect 12997 19068 13031 19102
rect 13069 19068 13103 19102
rect 13141 19068 13175 19102
rect 12997 18995 13031 19029
rect 13069 18995 13103 19029
rect 13141 18995 13175 19029
rect 12997 18922 13031 18956
rect 13069 18922 13103 18956
rect 13141 18922 13175 18956
rect 12997 18849 13031 18883
rect 13069 18849 13103 18883
rect 13141 18849 13175 18883
rect 12997 18776 13031 18810
rect 13069 18776 13103 18810
rect 13141 18776 13175 18810
rect 12997 18703 13031 18737
rect 13069 18703 13103 18737
rect 13141 18703 13175 18737
rect 13453 20229 13458 20263
rect 13458 20229 13487 20263
rect 13525 20229 13559 20263
rect 13597 20229 13628 20263
rect 13628 20229 13631 20263
rect 13453 20156 13458 20190
rect 13458 20156 13487 20190
rect 13525 20156 13559 20190
rect 13597 20156 13628 20190
rect 13628 20156 13631 20190
rect 13453 20083 13458 20117
rect 13458 20083 13487 20117
rect 13525 20083 13559 20117
rect 13597 20083 13628 20117
rect 13628 20083 13631 20117
rect 13453 20010 13458 20044
rect 13458 20010 13487 20044
rect 13525 20010 13559 20044
rect 13597 20010 13628 20044
rect 13628 20010 13631 20044
rect 13453 19937 13458 19971
rect 13458 19937 13487 19971
rect 13525 19937 13559 19971
rect 13597 19937 13628 19971
rect 13628 19937 13631 19971
rect 13453 19864 13458 19898
rect 13458 19864 13487 19898
rect 13525 19864 13559 19898
rect 13597 19864 13628 19898
rect 13628 19864 13631 19898
rect 13453 19791 13458 19825
rect 13458 19791 13487 19825
rect 13525 19791 13559 19825
rect 13597 19791 13628 19825
rect 13628 19791 13631 19825
rect 13453 19718 13458 19752
rect 13458 19718 13487 19752
rect 13525 19718 13559 19752
rect 13597 19718 13628 19752
rect 13628 19718 13631 19752
rect 13453 19645 13458 19679
rect 13458 19645 13487 19679
rect 13525 19645 13559 19679
rect 13597 19645 13628 19679
rect 13628 19645 13631 19679
rect 13453 19572 13458 19606
rect 13458 19572 13487 19606
rect 13525 19572 13559 19606
rect 13597 19572 13628 19606
rect 13628 19572 13631 19606
rect 13453 19499 13458 19533
rect 13458 19499 13487 19533
rect 13525 19499 13559 19533
rect 13597 19499 13628 19533
rect 13628 19499 13631 19533
rect 13453 19426 13458 19460
rect 13458 19426 13487 19460
rect 13525 19426 13559 19460
rect 13597 19426 13628 19460
rect 13628 19426 13631 19460
rect 13453 19353 13458 19387
rect 13458 19353 13487 19387
rect 13525 19353 13559 19387
rect 13597 19353 13628 19387
rect 13628 19353 13631 19387
rect 13453 19280 13458 19314
rect 13458 19280 13487 19314
rect 13525 19280 13559 19314
rect 13597 19280 13628 19314
rect 13628 19280 13631 19314
rect 13453 19207 13458 19241
rect 13458 19207 13487 19241
rect 13525 19207 13559 19241
rect 13597 19207 13628 19241
rect 13628 19207 13631 19241
rect 13453 19134 13458 19168
rect 13458 19134 13487 19168
rect 13525 19134 13559 19168
rect 13597 19134 13628 19168
rect 13628 19134 13631 19168
rect 13453 19061 13458 19095
rect 13458 19061 13487 19095
rect 13525 19061 13559 19095
rect 13597 19061 13628 19095
rect 13628 19061 13631 19095
rect 13453 18988 13458 19022
rect 13458 18988 13487 19022
rect 13525 18988 13559 19022
rect 13597 18988 13628 19022
rect 13628 18988 13631 19022
rect 13453 18915 13458 18949
rect 13458 18915 13487 18949
rect 13525 18915 13559 18949
rect 13597 18915 13628 18949
rect 13628 18915 13631 18949
rect 13453 18842 13458 18876
rect 13458 18842 13487 18876
rect 13525 18842 13559 18876
rect 13597 18842 13628 18876
rect 13628 18842 13631 18876
rect 13453 18769 13458 18803
rect 13458 18769 13487 18803
rect 13525 18769 13559 18803
rect 13597 18769 13628 18803
rect 13628 18769 13631 18803
rect 13453 18696 13458 18730
rect 13458 18696 13487 18730
rect 13525 18696 13559 18730
rect 13597 18696 13628 18730
rect 13628 18696 13631 18730
rect 13453 18623 13458 18657
rect 13458 18623 13487 18657
rect 13525 18623 13559 18657
rect 13597 18623 13628 18657
rect 13628 18623 13631 18657
rect 4358 18446 4362 18480
rect 4362 18446 4392 18480
rect 4430 18447 4464 18481
rect 4502 18447 4532 18481
rect 4532 18447 4536 18481
rect 4358 18373 4362 18407
rect 4362 18373 4392 18407
rect 4430 18374 4464 18408
rect 4502 18374 4532 18408
rect 4532 18374 4536 18408
rect 4358 18300 4362 18334
rect 4362 18300 4392 18334
rect 4430 18301 4464 18335
rect 4502 18301 4532 18335
rect 4532 18301 4536 18335
rect 4358 18227 4362 18261
rect 4362 18227 4392 18261
rect 4430 18228 4464 18262
rect 4502 18228 4532 18262
rect 4532 18228 4536 18262
rect 4358 18154 4362 18188
rect 4362 18154 4392 18188
rect 4430 18155 4464 18189
rect 4502 18155 4532 18189
rect 4532 18155 4536 18189
rect 4358 18081 4362 18115
rect 4362 18081 4392 18115
rect 4430 18082 4464 18116
rect 4502 18082 4532 18116
rect 4532 18082 4536 18116
rect 4611 18552 4645 18586
rect 4611 18479 4645 18513
rect 4611 18406 4645 18440
rect 4611 18333 4645 18367
rect 4611 18259 4645 18293
rect 4611 18185 4645 18219
rect 4611 18111 4645 18145
rect 13453 18550 13458 18584
rect 13458 18550 13487 18584
rect 13525 18550 13559 18584
rect 13597 18550 13628 18584
rect 13628 18550 13631 18584
rect 13453 18477 13458 18511
rect 13458 18477 13487 18511
rect 13525 18477 13559 18511
rect 13597 18477 13628 18511
rect 13628 18477 13631 18511
rect 13453 18404 13458 18438
rect 13458 18404 13487 18438
rect 13525 18404 13559 18438
rect 13597 18404 13628 18438
rect 13628 18404 13631 18438
rect 13453 18331 13458 18365
rect 13458 18331 13487 18365
rect 13525 18331 13559 18365
rect 13597 18331 13628 18365
rect 13628 18331 13631 18365
rect 13453 18258 13458 18292
rect 13458 18258 13487 18292
rect 13525 18258 13559 18292
rect 13597 18258 13628 18292
rect 13628 18258 13631 18292
rect 13453 18185 13458 18219
rect 13458 18185 13487 18219
rect 13525 18185 13559 18219
rect 13597 18185 13628 18219
rect 13628 18185 13631 18219
rect 13453 18112 13458 18146
rect 13458 18112 13487 18146
rect 13525 18112 13559 18146
rect 13597 18112 13628 18146
rect 13628 18112 13631 18146
rect 4358 18008 4362 18042
rect 4362 18008 4392 18042
rect 4430 18009 4464 18043
rect 4502 18009 4532 18043
rect 4532 18009 4536 18043
rect 13453 18039 13458 18073
rect 13458 18039 13487 18073
rect 13525 18039 13559 18073
rect 13597 18039 13628 18073
rect 13628 18039 13631 18073
rect 4358 17935 4362 17969
rect 4362 17935 4392 17969
rect 4430 17936 4464 17970
rect 4502 17936 4532 17970
rect 4532 17936 4536 17970
rect 4358 17862 4362 17896
rect 4362 17862 4392 17896
rect 4430 17863 4464 17897
rect 4502 17863 4532 17897
rect 4532 17863 4536 17897
rect 4358 17789 4362 17823
rect 4362 17789 4392 17823
rect 4430 17790 4464 17824
rect 4502 17790 4532 17824
rect 4532 17790 4536 17824
rect 4358 17716 4362 17750
rect 4362 17716 4392 17750
rect 4430 17717 4464 17751
rect 4502 17717 4532 17751
rect 4532 17717 4536 17751
rect 4358 17643 4362 17677
rect 4362 17643 4392 17677
rect 4430 17644 4464 17678
rect 4502 17644 4532 17678
rect 4532 17644 4536 17678
rect 4358 17570 4362 17604
rect 4362 17570 4392 17604
rect 4430 17571 4464 17605
rect 4502 17571 4532 17605
rect 4532 17571 4536 17605
rect 4358 17497 4362 17531
rect 4362 17497 4392 17531
rect 4430 17498 4464 17532
rect 4502 17498 4532 17532
rect 4532 17498 4536 17532
rect 4358 17424 4362 17458
rect 4362 17424 4392 17458
rect 4430 17425 4464 17459
rect 4502 17425 4532 17459
rect 4532 17425 4536 17459
rect 4358 17351 4362 17385
rect 4362 17351 4392 17385
rect 4430 17352 4464 17386
rect 4502 17352 4532 17386
rect 4532 17352 4536 17386
rect 4358 17278 4362 17312
rect 4362 17278 4392 17312
rect 4430 17279 4464 17313
rect 4502 17279 4532 17313
rect 4532 17279 4536 17313
rect 4358 17205 4362 17239
rect 4362 17205 4392 17239
rect 4430 17206 4464 17240
rect 4502 17206 4532 17240
rect 4532 17206 4536 17240
rect 4358 17132 4362 17166
rect 4362 17132 4392 17166
rect 4430 17133 4464 17167
rect 4502 17133 4532 17167
rect 4532 17133 4536 17167
rect 4358 17059 4362 17093
rect 4362 17059 4392 17093
rect 4430 17060 4464 17094
rect 4502 17060 4532 17094
rect 4532 17060 4536 17094
rect 4358 16986 4362 17020
rect 4362 16986 4392 17020
rect 4430 16987 4464 17021
rect 4502 16987 4532 17021
rect 4532 16987 4536 17021
rect 4358 16913 4362 16947
rect 4362 16913 4392 16947
rect 4430 16914 4464 16948
rect 4502 16914 4532 16948
rect 4532 16914 4536 16948
rect 4358 16840 4362 16874
rect 4362 16840 4392 16874
rect 4430 16841 4464 16875
rect 4502 16841 4532 16875
rect 4532 16841 4536 16875
rect 4358 16767 4362 16801
rect 4362 16767 4392 16801
rect 4430 16768 4464 16802
rect 4502 16768 4532 16802
rect 4532 16768 4536 16802
rect 4358 16694 4362 16728
rect 4362 16694 4392 16728
rect 4430 16695 4464 16729
rect 4502 16695 4532 16729
rect 4532 16695 4536 16729
rect 4358 16621 4362 16655
rect 4362 16621 4392 16655
rect 4430 16622 4464 16656
rect 4502 16622 4532 16656
rect 4532 16622 4536 16656
rect 4358 16548 4362 16582
rect 4362 16548 4392 16582
rect 4430 16549 4464 16583
rect 4502 16549 4532 16583
rect 4532 16549 4536 16583
rect 4358 16475 4362 16509
rect 4362 16475 4392 16509
rect 4430 16476 4464 16510
rect 4502 16476 4532 16510
rect 4532 16476 4536 16510
rect 4358 16402 4362 16436
rect 4362 16402 4392 16436
rect 4430 16403 4464 16437
rect 4502 16403 4532 16437
rect 4532 16403 4536 16437
rect 4358 16329 4362 16363
rect 4362 16329 4392 16363
rect 4430 16330 4464 16364
rect 4502 16330 4532 16364
rect 4532 16330 4536 16364
rect 4358 16256 4362 16290
rect 4362 16256 4392 16290
rect 4430 16257 4464 16291
rect 4502 16257 4532 16291
rect 4532 16257 4536 16291
rect 4358 16183 4362 16217
rect 4362 16183 4392 16217
rect 4430 16184 4464 16218
rect 4502 16184 4532 16218
rect 4532 16184 4536 16218
rect 4358 16110 4362 16144
rect 4362 16110 4392 16144
rect 4430 16111 4464 16145
rect 4502 16111 4532 16145
rect 4532 16111 4536 16145
rect 4358 16037 4362 16071
rect 4362 16037 4392 16071
rect 4430 16038 4464 16072
rect 4502 16038 4532 16072
rect 4532 16038 4536 16072
rect 4358 15964 4362 15998
rect 4362 15964 4392 15998
rect 4430 15965 4464 15999
rect 4502 15965 4532 15999
rect 4532 15965 4536 15999
rect 4358 15891 4362 15925
rect 4362 15891 4392 15925
rect 4430 15892 4464 15926
rect 4502 15892 4532 15926
rect 4532 15892 4536 15926
rect 4358 15818 4362 15852
rect 4362 15818 4392 15852
rect 4430 15819 4464 15853
rect 4502 15819 4532 15853
rect 4532 15819 4536 15853
rect 4358 15745 4362 15779
rect 4362 15745 4392 15779
rect 4430 15746 4464 15780
rect 4502 15746 4532 15780
rect 4532 15746 4536 15780
rect 4358 15672 4362 15706
rect 4362 15672 4392 15706
rect 4430 15673 4464 15707
rect 4502 15673 4532 15707
rect 4532 15673 4536 15707
rect 4358 15599 4362 15633
rect 4362 15599 4392 15633
rect 4430 15600 4464 15634
rect 4502 15600 4532 15634
rect 4532 15600 4536 15634
rect 4358 15526 4362 15560
rect 4362 15526 4392 15560
rect 4430 15527 4464 15561
rect 4502 15527 4532 15561
rect 4532 15527 4536 15561
rect 4358 15453 4362 15487
rect 4362 15453 4392 15487
rect 4430 15454 4464 15488
rect 4502 15454 4532 15488
rect 4532 15454 4536 15488
rect 4358 15380 4362 15414
rect 4362 15380 4392 15414
rect 4430 15381 4464 15415
rect 4502 15381 4532 15415
rect 4532 15381 4536 15415
rect 4358 15307 4362 15341
rect 4362 15307 4392 15341
rect 4430 15308 4464 15342
rect 4502 15308 4532 15342
rect 4532 15308 4536 15342
rect 4358 15234 4362 15268
rect 4362 15234 4392 15268
rect 4430 15235 4464 15269
rect 4502 15235 4532 15269
rect 4532 15235 4536 15269
rect 4358 15161 4362 15195
rect 4362 15161 4392 15195
rect 4430 15162 4464 15196
rect 4502 15162 4532 15196
rect 4532 15162 4536 15196
rect 4358 15088 4362 15122
rect 4362 15088 4392 15122
rect 4430 15089 4464 15123
rect 4502 15089 4532 15123
rect 4532 15089 4536 15123
rect 4358 15015 4362 15049
rect 4362 15015 4392 15049
rect 4430 15016 4464 15050
rect 4502 15016 4532 15050
rect 4532 15016 4536 15050
rect 4358 14942 4362 14976
rect 4362 14942 4392 14976
rect 4430 14943 4464 14977
rect 4502 14943 4532 14977
rect 4532 14943 4536 14977
rect 4358 14869 4362 14903
rect 4362 14869 4392 14903
rect 4430 14870 4464 14904
rect 4502 14870 4532 14904
rect 4532 14870 4536 14904
rect 4358 14796 4362 14830
rect 4362 14796 4392 14830
rect 4430 14797 4464 14831
rect 4502 14797 4532 14831
rect 4532 14797 4536 14831
rect 4358 14723 4362 14757
rect 4362 14723 4392 14757
rect 4430 14724 4464 14758
rect 4502 14724 4532 14758
rect 4532 14724 4536 14758
rect 4358 14650 4362 14684
rect 4362 14650 4392 14684
rect 4430 14651 4464 14685
rect 4502 14651 4532 14685
rect 4532 14651 4536 14685
rect 4358 14577 4362 14611
rect 4362 14577 4392 14611
rect 4430 14578 4464 14612
rect 4502 14578 4532 14612
rect 4532 14578 4536 14612
rect 4358 14504 4362 14538
rect 4362 14504 4392 14538
rect 4430 14505 4464 14539
rect 4502 14505 4532 14539
rect 4532 14505 4536 14539
rect 4358 14431 4362 14465
rect 4362 14431 4392 14465
rect 4430 14432 4464 14466
rect 4502 14432 4532 14466
rect 4532 14432 4536 14466
rect 4358 14358 4362 14392
rect 4362 14358 4392 14392
rect 4430 14359 4464 14393
rect 4502 14359 4532 14393
rect 4532 14359 4536 14393
rect 4358 14285 4362 14319
rect 4362 14285 4392 14319
rect 4430 14286 4464 14320
rect 4502 14286 4532 14320
rect 4532 14286 4536 14320
rect 4358 14212 4362 14246
rect 4362 14212 4392 14246
rect 4430 14213 4464 14247
rect 4502 14213 4532 14247
rect 4532 14213 4536 14247
rect 1827 13809 1834 13843
rect 1834 13809 1861 13843
rect 1899 13809 1933 13843
rect 1971 13809 2005 13843
rect 2043 13809 2072 13843
rect 2072 13809 2077 13843
rect 1827 13736 1834 13770
rect 1834 13736 1861 13770
rect 1899 13736 1933 13770
rect 1971 13736 2005 13770
rect 2043 13736 2072 13770
rect 2072 13736 2077 13770
rect 1827 13663 1834 13697
rect 1834 13663 1861 13697
rect 1899 13663 1933 13697
rect 1971 13663 2005 13697
rect 2043 13663 2072 13697
rect 2072 13663 2077 13697
rect 1827 13590 1834 13624
rect 1834 13590 1861 13624
rect 1899 13590 1933 13624
rect 1971 13590 2005 13624
rect 2043 13590 2072 13624
rect 2072 13590 2077 13624
rect 1827 12861 1834 13543
rect 1834 13005 2072 13543
rect 2072 13005 2077 13543
rect 1834 12933 2005 13005
rect 1834 12861 1933 12933
rect 2043 12932 2072 12966
rect 2072 12932 2077 12966
rect 1971 12860 2005 12894
rect 2043 12859 2072 12893
rect 2072 12859 2077 12893
rect 1827 12788 1834 12822
rect 1834 12788 1861 12822
rect 1899 12788 1933 12822
rect 1971 12787 2005 12821
rect 2043 12786 2072 12820
rect 2072 12786 2077 12820
rect 1827 12715 1834 12749
rect 1834 12715 1861 12749
rect 1899 12715 1933 12749
rect 1971 12714 2005 12748
rect 2043 12713 2072 12747
rect 2072 12713 2077 12747
rect 1827 12642 1834 12676
rect 1834 12642 1861 12676
rect 1899 12642 1933 12676
rect 1971 12641 2005 12675
rect 2043 12640 2072 12674
rect 2072 12640 2077 12674
rect 1827 12569 1834 12603
rect 1834 12569 1861 12603
rect 1899 12569 1933 12603
rect 1971 12568 2005 12602
rect 2043 12567 2072 12601
rect 2072 12567 2077 12601
rect 1827 12496 1834 12530
rect 1834 12496 1861 12530
rect 1899 12496 1933 12530
rect 1971 12495 2005 12529
rect 2043 12494 2072 12528
rect 2072 12494 2077 12528
rect 1827 12423 1834 12457
rect 1834 12423 1861 12457
rect 1899 12423 1933 12457
rect 1971 12422 2005 12456
rect 2043 12421 2072 12455
rect 2072 12421 2077 12455
rect 1827 12350 1834 12384
rect 1834 12350 1861 12384
rect 1899 12350 1933 12384
rect 1971 12349 2005 12383
rect 2043 12348 2072 12382
rect 2072 12348 2077 12382
rect 1827 12277 1834 12311
rect 1834 12277 1861 12311
rect 1899 12277 1933 12311
rect 1971 12276 2005 12310
rect 2043 12275 2072 12309
rect 2072 12275 2077 12309
rect 1827 12204 1834 12238
rect 1834 12204 1861 12238
rect 1899 12204 1933 12238
rect 1971 12203 2005 12237
rect 2043 12202 2072 12236
rect 2072 12202 2077 12236
rect 1827 12131 1834 12165
rect 1834 12131 1861 12165
rect 1899 12131 1933 12165
rect 1971 12130 2005 12164
rect 2043 12129 2072 12163
rect 2072 12129 2077 12163
rect 1827 12058 1834 12092
rect 1834 12058 1861 12092
rect 1899 12058 1933 12092
rect 1971 12057 2005 12091
rect 2043 12056 2072 12090
rect 2072 12056 2077 12090
rect 1827 11985 1834 12019
rect 1834 11985 1861 12019
rect 1899 11985 1933 12019
rect 1971 11984 2005 12018
rect 2043 11983 2072 12017
rect 2072 11983 2077 12017
rect 1827 11912 1834 11946
rect 1834 11912 1861 11946
rect 1899 11912 1933 11946
rect 1971 11911 2005 11945
rect 2043 11910 2072 11944
rect 2072 11910 2077 11944
rect 1827 11839 1834 11873
rect 1834 11839 1861 11873
rect 1899 11839 1933 11873
rect 1971 11838 2005 11872
rect 2043 11837 2072 11871
rect 2072 11837 2077 11871
rect 1827 11766 1834 11800
rect 1834 11766 1861 11800
rect 1899 11766 1933 11800
rect 1971 11765 2005 11799
rect 2043 11764 2072 11798
rect 2072 11764 2077 11798
rect 1827 11693 1834 11727
rect 1834 11693 1861 11727
rect 1899 11693 1933 11727
rect 1971 11692 2005 11726
rect 2043 11691 2072 11725
rect 2072 11691 2077 11725
rect 1827 11620 1834 11654
rect 1834 11620 1861 11654
rect 1899 11620 1933 11654
rect 1971 11619 2005 11653
rect 2043 11618 2072 11652
rect 2072 11618 2077 11652
rect 1827 11547 1834 11581
rect 1834 11547 1861 11581
rect 1899 11547 1933 11581
rect 1971 11546 2005 11580
rect 2043 11545 2072 11579
rect 2072 11545 2077 11579
rect 1827 11474 1834 11508
rect 1834 11474 1861 11508
rect 1899 11474 1933 11508
rect 1971 11473 2005 11507
rect 2043 11472 2072 11506
rect 2072 11472 2077 11506
rect 1827 11401 1834 11435
rect 1834 11401 1861 11435
rect 1899 11401 1933 11435
rect 1971 11400 2005 11434
rect 2043 11399 2072 11433
rect 2072 11399 2077 11433
rect 1827 11328 1834 11362
rect 1834 11328 1861 11362
rect 1899 11328 1933 11362
rect 1971 11327 2005 11361
rect 2043 11326 2072 11360
rect 2072 11326 2077 11360
rect 1827 11255 1834 11289
rect 1834 11255 1861 11289
rect 1899 11255 1933 11289
rect 1971 11254 2005 11288
rect 2043 11253 2072 11287
rect 2072 11253 2077 11287
rect 1827 11182 1834 11216
rect 1834 11182 1861 11216
rect 1899 11182 1933 11216
rect 1971 11181 2005 11215
rect 2043 11180 2072 11214
rect 2072 11180 2077 11214
rect 1827 11109 1834 11143
rect 1834 11109 1861 11143
rect 1899 11109 1933 11143
rect 1971 11108 2005 11142
rect 2043 11107 2072 11141
rect 2072 11107 2077 11141
rect 1827 11036 1834 11070
rect 1834 11036 1861 11070
rect 1899 11036 1933 11070
rect 1971 11035 2005 11069
rect 2043 11034 2072 11068
rect 2072 11034 2077 11068
rect 1827 10963 1834 10997
rect 1834 10963 1861 10997
rect 1899 10963 1933 10997
rect 1971 10962 2005 10996
rect 2043 10961 2072 10995
rect 2072 10961 2077 10995
rect 1827 10890 1834 10924
rect 1834 10890 1861 10924
rect 1899 10890 1933 10924
rect 1971 10889 2005 10923
rect 2043 10888 2072 10922
rect 2072 10888 2077 10922
rect 1827 10817 1861 10851
rect 1899 10817 1933 10851
rect 1971 10816 2005 10850
rect 2043 10815 2077 10849
rect 1827 10746 1861 10778
rect 1899 10746 1933 10778
rect 1971 10746 2005 10777
rect 2043 10746 2077 10776
rect 1827 10744 1834 10746
rect 1834 10744 1861 10746
rect 1899 10744 1933 10746
rect 1971 10743 2005 10746
rect 2043 10742 2072 10746
rect 2072 10742 2077 10746
rect 1827 10671 1834 10705
rect 1834 10671 1861 10705
rect 1899 10671 1933 10705
rect 1971 10670 2005 10704
rect 2043 10669 2072 10703
rect 2072 10669 2077 10703
rect 1827 10598 1834 10632
rect 1834 10598 1861 10632
rect 1899 10598 1933 10632
rect 1971 10597 2005 10631
rect 2043 10596 2072 10630
rect 2072 10596 2077 10630
rect 1827 10525 1834 10559
rect 1834 10525 1861 10559
rect 1899 10525 1933 10559
rect 1971 10524 2005 10558
rect 2043 10523 2072 10557
rect 2072 10523 2077 10557
rect 1827 10452 1834 10486
rect 1834 10452 1861 10486
rect 1899 10452 1933 10486
rect 1971 10451 2005 10485
rect 2043 10450 2072 10484
rect 2072 10450 2077 10484
rect 1827 10379 1834 10413
rect 1834 10379 1861 10413
rect 1899 10379 1933 10413
rect 1971 10378 2005 10412
rect 2043 10377 2072 10411
rect 2072 10377 2077 10411
rect 1827 10306 1834 10340
rect 1834 10306 1861 10340
rect 1899 10306 1933 10340
rect 1971 10305 2005 10339
rect 2043 10304 2072 10338
rect 2072 10304 2077 10338
rect 1827 10233 1834 10267
rect 1834 10233 1861 10267
rect 1899 10233 1933 10267
rect 1971 10232 2005 10266
rect 2043 10231 2072 10265
rect 2072 10231 2077 10265
rect 1827 10160 1834 10194
rect 1834 10160 1861 10194
rect 1899 10160 1933 10194
rect 1971 10159 2005 10193
rect 2043 10158 2072 10192
rect 2072 10158 2077 10192
rect 1827 10087 1834 10121
rect 1834 10087 1861 10121
rect 1899 10087 1933 10121
rect 1971 10086 2005 10120
rect 2043 10085 2072 10119
rect 2072 10085 2077 10119
rect 1827 10014 1834 10048
rect 1834 10014 1861 10048
rect 1899 10014 1933 10048
rect 1971 10013 2005 10047
rect 2043 10012 2072 10046
rect 2072 10012 2077 10046
rect 1827 9941 1834 9975
rect 1834 9941 1861 9975
rect 1899 9941 1933 9975
rect 1971 9940 2005 9974
rect 2043 9939 2072 9973
rect 2072 9939 2077 9973
rect 1827 9868 1834 9902
rect 1834 9868 1861 9902
rect 1899 9868 1933 9902
rect 1971 9867 2005 9901
rect 2043 9866 2072 9900
rect 2072 9866 2077 9900
rect 1827 9795 1834 9829
rect 1834 9795 1861 9829
rect 1899 9795 1933 9829
rect 1971 9794 2005 9828
rect 2043 9793 2072 9827
rect 2072 9793 2077 9827
rect 1827 9722 1834 9756
rect 1834 9722 1861 9756
rect 1899 9722 1933 9756
rect 1971 9721 2005 9755
rect 2043 9720 2072 9754
rect 2072 9720 2077 9754
rect 1827 9649 1834 9683
rect 1834 9649 1861 9683
rect 1899 9649 1933 9683
rect 1971 9648 2005 9682
rect 2043 9647 2072 9681
rect 2072 9647 2077 9681
rect 1827 9576 1834 9610
rect 1834 9576 1861 9610
rect 1899 9576 1933 9610
rect 1971 9575 2005 9609
rect 2043 9574 2072 9608
rect 2072 9574 2077 9608
rect 1827 9503 1834 9537
rect 1834 9503 1861 9537
rect 1899 9503 1933 9537
rect 1971 9502 2005 9536
rect 2043 9501 2072 9535
rect 2072 9501 2077 9535
rect 1827 9430 1834 9464
rect 1834 9430 1861 9464
rect 1899 9430 1933 9464
rect 1971 9429 2005 9463
rect 2043 9428 2072 9462
rect 2072 9428 2077 9462
rect 1827 9357 1834 9391
rect 1834 9357 1861 9391
rect 1899 9357 1933 9391
rect 1971 9356 2005 9390
rect 2043 9355 2072 9389
rect 2072 9355 2077 9389
rect 1827 9284 1834 9318
rect 1834 9284 1861 9318
rect 1899 9284 1933 9318
rect 1971 9283 2005 9317
rect 2043 9282 2072 9316
rect 2072 9282 2077 9316
rect 1827 9211 1834 9245
rect 1834 9211 1861 9245
rect 1899 9211 1933 9245
rect 1971 9210 2005 9244
rect 2043 9209 2072 9243
rect 2072 9209 2077 9243
rect 1827 9138 1834 9172
rect 1834 9138 1861 9172
rect 1899 9138 1933 9172
rect 1971 9137 2005 9171
rect 2043 9136 2072 9170
rect 2072 9136 2077 9170
rect 1827 9065 1834 9099
rect 1834 9065 1861 9099
rect 1899 9065 1933 9099
rect 1971 9064 2005 9098
rect 2043 9063 2072 9097
rect 2072 9063 2077 9097
rect 2293 14169 2327 14173
rect 2367 14169 2401 14173
rect 2441 14169 2475 14173
rect 2515 14169 2549 14173
rect 2589 14169 2623 14173
rect 2663 14169 2697 14173
rect 2737 14169 2771 14173
rect 2811 14169 2845 14173
rect 2885 14169 2919 14173
rect 2959 14169 2993 14173
rect 3033 14169 3067 14173
rect 3107 14169 3141 14173
rect 3181 14169 3215 14173
rect 3255 14169 3289 14173
rect 3329 14169 3363 14173
rect 3403 14169 3437 14173
rect 3477 14169 3511 14173
rect 3551 14169 3585 14173
rect 3625 14169 3659 14173
rect 3699 14169 3733 14173
rect 3773 14169 3807 14173
rect 3847 14169 3881 14173
rect 3920 14169 3954 14173
rect 3993 14169 4027 14173
rect 4066 14169 4100 14173
rect 4139 14169 4173 14173
rect 4212 14169 4246 14173
rect 4285 14169 4319 14173
rect 4358 14169 4392 14173
rect 2293 14139 2322 14169
rect 2322 14139 2327 14169
rect 2367 14139 2390 14169
rect 2390 14139 2401 14169
rect 2441 14139 2475 14169
rect 2515 14139 2549 14169
rect 2589 14139 2623 14169
rect 2663 14139 2697 14169
rect 2737 14139 2771 14169
rect 2811 14139 2845 14169
rect 2885 14139 2919 14169
rect 2959 14139 2993 14169
rect 3033 14139 3067 14169
rect 3107 14139 3141 14169
rect 3181 14139 3215 14169
rect 3255 14139 3289 14169
rect 3329 14139 3363 14169
rect 3403 14139 3437 14169
rect 3477 14139 3511 14169
rect 3551 14139 3585 14169
rect 3625 14139 3659 14169
rect 3699 14139 3733 14169
rect 3773 14139 3807 14169
rect 3847 14139 3881 14169
rect 3920 14139 3954 14169
rect 3993 14139 4027 14169
rect 4066 14139 4100 14169
rect 4139 14139 4173 14169
rect 4212 14139 4246 14169
rect 4285 14139 4319 14169
rect 4358 14139 4392 14169
rect 4430 14143 4464 14174
rect 4502 14143 4532 14174
rect 4532 14143 4536 14174
rect 4430 14140 4464 14143
rect 4502 14140 4536 14143
rect 2221 14061 2225 14095
rect 2225 14061 2255 14095
rect 2293 14067 2327 14101
rect 2367 14067 2390 14101
rect 2390 14067 2401 14101
rect 2441 14067 2475 14101
rect 2515 14067 2549 14101
rect 2589 14067 2623 14101
rect 2663 14067 2697 14101
rect 2737 14067 2771 14101
rect 2811 14067 2845 14101
rect 2885 14067 2919 14101
rect 2959 14067 2993 14101
rect 3033 14067 3067 14101
rect 3107 14067 3141 14101
rect 3181 14067 3215 14101
rect 3255 14067 3289 14101
rect 3329 14067 3363 14101
rect 3403 14067 3437 14101
rect 3477 14067 3511 14101
rect 3551 14067 3585 14101
rect 3625 14067 3659 14101
rect 3699 14067 3733 14101
rect 3772 14067 3806 14101
rect 3845 14067 3879 14101
rect 3918 14067 3952 14101
rect 3991 14067 4025 14101
rect 4064 14067 4098 14101
rect 4137 14067 4171 14101
rect 4210 14067 4244 14101
rect 4283 14067 4317 14101
rect 4356 14067 4390 14101
rect 4430 14067 4464 14101
rect 4502 14075 4532 14101
rect 4532 14075 4536 14101
rect 4502 14067 4536 14075
rect 2221 13983 2225 14017
rect 2225 13983 2255 14017
rect 2293 13983 2327 14017
rect 2365 13995 2395 14029
rect 2395 13995 2399 14029
rect 2439 13999 2458 14029
rect 2458 13999 2473 14029
rect 2513 13999 2547 14029
rect 2587 13999 2621 14029
rect 2661 13999 2695 14029
rect 2735 13999 2769 14029
rect 2809 13999 2843 14029
rect 2883 13999 2917 14029
rect 2957 13999 2991 14029
rect 3031 13999 3065 14029
rect 3105 13999 3139 14029
rect 3179 13999 3213 14029
rect 3253 13999 3287 14029
rect 3327 13999 3361 14029
rect 3401 13999 3435 14029
rect 3475 13999 3509 14029
rect 3549 13999 3583 14029
rect 3623 13999 3657 14029
rect 3697 13999 3731 14029
rect 3771 13999 3805 14029
rect 3845 13999 3879 14029
rect 3918 13999 3952 14029
rect 3991 13999 4025 14029
rect 4064 13999 4098 14029
rect 4137 13999 4171 14029
rect 4210 13999 4244 14029
rect 4283 13999 4317 14029
rect 4356 13999 4390 14029
rect 4429 13999 4463 14029
rect 4717 14760 4895 17962
rect 4717 14687 4751 14721
rect 4789 14687 4823 14721
rect 4861 14687 4895 14721
rect 4717 14614 4751 14648
rect 4789 14614 4823 14648
rect 4861 14614 4895 14648
rect 4717 14541 4751 14575
rect 4789 14541 4823 14575
rect 4861 14541 4895 14575
rect 4717 14468 4751 14502
rect 4789 14468 4823 14502
rect 4861 14468 4895 14502
rect 4717 14395 4751 14429
rect 4789 14395 4823 14429
rect 4861 14395 4895 14429
rect 4717 14322 4751 14356
rect 4789 14322 4823 14356
rect 4861 14322 4895 14356
rect 4717 14249 4751 14283
rect 4789 14249 4823 14283
rect 4861 14249 4895 14283
rect 4717 14176 4751 14210
rect 4789 14176 4823 14210
rect 4861 14176 4895 14210
rect 4717 14103 4751 14137
rect 4789 14103 4823 14137
rect 4861 14103 4895 14137
rect 5637 14760 5815 17962
rect 5637 14687 5671 14721
rect 5709 14687 5743 14721
rect 5781 14687 5815 14721
rect 5637 14614 5671 14648
rect 5709 14614 5743 14648
rect 5781 14614 5815 14648
rect 5637 14541 5671 14575
rect 5709 14541 5743 14575
rect 5781 14541 5815 14575
rect 5637 14468 5671 14502
rect 5709 14468 5743 14502
rect 5781 14468 5815 14502
rect 5637 14395 5671 14429
rect 5709 14395 5743 14429
rect 5781 14395 5815 14429
rect 5637 14322 5671 14356
rect 5709 14322 5743 14356
rect 5781 14322 5815 14356
rect 5637 14249 5671 14283
rect 5709 14249 5743 14283
rect 5781 14249 5815 14283
rect 5637 14176 5671 14210
rect 5709 14176 5743 14210
rect 5781 14176 5815 14210
rect 5637 14103 5671 14137
rect 5709 14103 5743 14137
rect 5781 14103 5815 14137
rect 6557 14103 6735 17953
rect 7477 14103 7655 17953
rect 8397 14103 8575 17953
rect 9317 14103 9495 17953
rect 10237 14103 10415 17953
rect 11157 14103 11335 17953
rect 12077 14103 12255 17953
rect 12997 14103 13175 17953
rect 13453 17966 13458 18000
rect 13458 17966 13487 18000
rect 13525 17966 13559 18000
rect 13597 17966 13628 18000
rect 13628 17966 13631 18000
rect 13453 17893 13458 17927
rect 13458 17893 13487 17927
rect 13525 17893 13559 17927
rect 13597 17893 13628 17927
rect 13628 17893 13631 17927
rect 13453 17820 13458 17854
rect 13458 17820 13487 17854
rect 13525 17820 13559 17854
rect 13597 17820 13628 17854
rect 13628 17820 13631 17854
rect 13453 17747 13458 17781
rect 13458 17747 13487 17781
rect 13525 17747 13559 17781
rect 13597 17747 13628 17781
rect 13628 17747 13631 17781
rect 13453 17674 13458 17708
rect 13458 17674 13487 17708
rect 13525 17674 13559 17708
rect 13597 17674 13628 17708
rect 13628 17674 13631 17708
rect 13453 17601 13458 17635
rect 13458 17601 13487 17635
rect 13525 17601 13559 17635
rect 13597 17601 13628 17635
rect 13628 17601 13631 17635
rect 13453 17528 13458 17562
rect 13458 17528 13487 17562
rect 13525 17528 13559 17562
rect 13597 17528 13628 17562
rect 13628 17528 13631 17562
rect 13453 17455 13458 17489
rect 13458 17455 13487 17489
rect 13525 17455 13559 17489
rect 13597 17455 13628 17489
rect 13628 17455 13631 17489
rect 13453 17382 13458 17416
rect 13458 17382 13487 17416
rect 13525 17382 13559 17416
rect 13597 17382 13628 17416
rect 13628 17382 13631 17416
rect 13453 17309 13458 17343
rect 13458 17309 13487 17343
rect 13525 17309 13559 17343
rect 13597 17309 13628 17343
rect 13628 17309 13631 17343
rect 13453 17236 13458 17270
rect 13458 17236 13487 17270
rect 13525 17236 13559 17270
rect 13597 17236 13628 17270
rect 13628 17236 13631 17270
rect 13453 17163 13458 17197
rect 13458 17163 13487 17197
rect 13525 17163 13559 17197
rect 13597 17163 13628 17197
rect 13628 17163 13631 17197
rect 13453 17090 13458 17124
rect 13458 17090 13487 17124
rect 13525 17090 13559 17124
rect 13597 17090 13628 17124
rect 13628 17090 13631 17124
rect 13453 17017 13458 17051
rect 13458 17017 13487 17051
rect 13525 17017 13559 17051
rect 13597 17017 13628 17051
rect 13628 17017 13631 17051
rect 13453 16944 13458 16978
rect 13458 16944 13487 16978
rect 13525 16944 13559 16978
rect 13597 16944 13628 16978
rect 13628 16944 13631 16978
rect 13453 16871 13458 16905
rect 13458 16871 13487 16905
rect 13525 16871 13559 16905
rect 13597 16871 13628 16905
rect 13628 16871 13631 16905
rect 13453 16798 13458 16832
rect 13458 16798 13487 16832
rect 13525 16798 13559 16832
rect 13597 16798 13628 16832
rect 13628 16798 13631 16832
rect 13453 16725 13458 16759
rect 13458 16725 13487 16759
rect 13525 16725 13559 16759
rect 13597 16725 13628 16759
rect 13628 16725 13631 16759
rect 2439 13995 2473 13999
rect 2513 13995 2547 13999
rect 2587 13995 2621 13999
rect 2661 13995 2695 13999
rect 2735 13995 2769 13999
rect 2809 13995 2843 13999
rect 2883 13995 2917 13999
rect 2957 13995 2991 13999
rect 3031 13995 3065 13999
rect 3105 13995 3139 13999
rect 3179 13995 3213 13999
rect 3253 13995 3287 13999
rect 3327 13995 3361 13999
rect 3401 13995 3435 13999
rect 3475 13995 3509 13999
rect 3549 13995 3583 13999
rect 3623 13995 3657 13999
rect 3697 13995 3731 13999
rect 3771 13995 3805 13999
rect 3845 13995 3879 13999
rect 3918 13995 3952 13999
rect 3991 13995 4025 13999
rect 4064 13995 4098 13999
rect 4137 13995 4171 13999
rect 4210 13995 4244 13999
rect 4283 13995 4317 13999
rect 4356 13995 4390 13999
rect 4429 13995 4463 13999
rect 2221 13905 2225 13939
rect 2225 13905 2255 13939
rect 2293 13905 2327 13939
rect 2365 13915 2395 13949
rect 2395 13915 2399 13949
rect 2221 13827 2225 13861
rect 2225 13827 2255 13861
rect 2293 13827 2327 13861
rect 2365 13835 2395 13869
rect 2395 13835 2399 13869
rect 2221 13749 2225 13783
rect 2225 13749 2255 13783
rect 2293 13749 2327 13783
rect 2365 13755 2395 13789
rect 2395 13755 2399 13789
rect 2221 13671 2225 13705
rect 2225 13671 2255 13705
rect 2293 13671 2327 13705
rect 2365 13674 2395 13708
rect 2395 13674 2399 13708
rect 2221 13593 2225 13627
rect 2225 13593 2255 13627
rect 2293 13593 2327 13627
rect 2365 13593 2395 13627
rect 2395 13593 2399 13627
rect 3157 13608 3191 13642
rect 3230 13608 3264 13642
rect 3303 13608 3337 13642
rect 3376 13608 3410 13642
rect 3449 13608 3483 13642
rect 3522 13608 3556 13642
rect 3595 13608 3629 13642
rect 3668 13608 3702 13642
rect 3741 13608 3775 13642
rect 3813 13608 3847 13642
rect 3885 13608 3919 13642
rect 3957 13608 3991 13642
rect 4029 13608 4063 13642
rect 4101 13608 4135 13642
rect 4173 13608 4207 13642
rect 4245 13608 4279 13642
rect 4317 13608 4351 13642
rect 4389 13608 4423 13642
rect 4461 13608 4495 13642
rect 4533 13608 4567 13642
rect 4605 13608 4639 13642
rect 2221 11755 2225 13544
rect 2225 11755 2395 13544
rect 2395 11755 2399 13544
rect 2221 11659 2399 11755
rect 2221 11062 2225 11659
rect 2225 11134 2395 11659
rect 2395 11134 2399 11659
rect 2225 11062 2327 11134
rect 2365 11061 2395 11095
rect 2395 11061 2399 11095
rect 2221 10989 2225 11023
rect 2225 10989 2255 11023
rect 2293 10989 2327 11023
rect 2365 10988 2395 11022
rect 2395 10988 2399 11022
rect 2221 10916 2225 10950
rect 2225 10916 2255 10950
rect 2293 10916 2327 10950
rect 2365 10915 2395 10949
rect 2395 10915 2399 10949
rect 2221 10843 2225 10877
rect 2225 10843 2255 10877
rect 2293 10843 2327 10877
rect 2365 10842 2395 10876
rect 2395 10842 2399 10876
rect 2221 10770 2225 10804
rect 2225 10770 2255 10804
rect 2293 10770 2327 10804
rect 2365 10769 2395 10803
rect 2395 10769 2399 10803
rect 2221 10697 2225 10731
rect 2225 10697 2255 10731
rect 2293 10697 2327 10731
rect 2365 10696 2395 10730
rect 2395 10696 2399 10730
rect 2221 10624 2225 10658
rect 2225 10624 2255 10658
rect 2293 10624 2327 10658
rect 2365 10623 2395 10657
rect 2395 10623 2399 10657
rect 2221 10551 2225 10585
rect 2225 10551 2255 10585
rect 2293 10551 2327 10585
rect 2365 10550 2395 10584
rect 2395 10550 2399 10584
rect 2221 10478 2225 10512
rect 2225 10478 2255 10512
rect 2293 10478 2327 10512
rect 2365 10477 2395 10511
rect 2395 10477 2399 10511
rect 2221 10405 2225 10439
rect 2225 10405 2255 10439
rect 2293 10405 2327 10439
rect 2365 10404 2395 10438
rect 2395 10404 2399 10438
rect 2221 10332 2225 10366
rect 2225 10332 2255 10366
rect 2293 10332 2327 10366
rect 2365 10331 2395 10365
rect 2395 10331 2399 10365
rect 2221 10259 2225 10293
rect 2225 10259 2255 10293
rect 2293 10259 2327 10293
rect 2365 10258 2395 10292
rect 2395 10258 2399 10292
rect 2221 10186 2225 10220
rect 2225 10186 2255 10220
rect 2293 10186 2327 10220
rect 2365 10185 2395 10219
rect 2395 10185 2399 10219
rect 2221 10113 2225 10147
rect 2225 10113 2255 10147
rect 2293 10113 2327 10147
rect 2365 10112 2395 10146
rect 2395 10112 2399 10146
rect 2221 10040 2225 10074
rect 2225 10040 2255 10074
rect 2293 10040 2327 10074
rect 2365 10039 2395 10073
rect 2395 10039 2399 10073
rect 2221 9967 2225 10001
rect 2225 9967 2255 10001
rect 2293 9967 2327 10001
rect 2365 9966 2395 10000
rect 2395 9966 2399 10000
rect 2221 9894 2225 9928
rect 2225 9894 2255 9928
rect 2293 9894 2327 9928
rect 2365 9893 2395 9927
rect 2395 9893 2399 9927
rect 2221 9821 2225 9855
rect 2225 9821 2255 9855
rect 2293 9821 2327 9855
rect 2365 9820 2395 9854
rect 2395 9820 2399 9854
rect 2221 9748 2225 9782
rect 2225 9748 2255 9782
rect 2293 9748 2327 9782
rect 2365 9747 2395 9781
rect 2395 9747 2399 9781
rect 2221 9675 2225 9709
rect 2225 9675 2255 9709
rect 2293 9675 2327 9709
rect 2365 9674 2395 9708
rect 2395 9674 2399 9708
rect 2221 9602 2225 9636
rect 2225 9602 2255 9636
rect 2293 9602 2327 9636
rect 2365 9601 2395 9635
rect 2395 9601 2399 9635
rect 2221 9529 2225 9563
rect 2225 9529 2255 9563
rect 2293 9529 2327 9563
rect 2365 9528 2395 9562
rect 2395 9528 2399 9562
rect 2221 9456 2225 9490
rect 2225 9456 2255 9490
rect 2293 9456 2327 9490
rect 2365 9455 2395 9489
rect 2395 9455 2399 9489
rect 2221 9383 2225 9417
rect 2225 9383 2255 9417
rect 2293 9383 2327 9417
rect 2365 9382 2395 9416
rect 2395 9382 2399 9416
rect 2221 9310 2225 9344
rect 2225 9310 2255 9344
rect 2293 9310 2327 9344
rect 2617 13559 2651 13593
rect 2617 13487 2651 13521
rect 2617 13415 2651 13449
rect 2617 13343 2651 13377
rect 2617 13271 2651 13305
rect 2617 13199 2651 13233
rect 2617 13127 2651 13161
rect 2617 13055 2651 13089
rect 2617 12983 2651 13017
rect 2617 12911 2651 12945
rect 2617 12839 2651 12873
rect 2617 12767 2651 12801
rect 2617 12695 2651 12729
rect 2617 12623 2651 12657
rect 2617 12551 2651 12585
rect 2617 12479 2651 12513
rect 2617 12407 2651 12441
rect 2617 12335 2651 12369
rect 2617 12263 2651 12297
rect 2617 12191 2651 12225
rect 2617 12119 2651 12153
rect 2617 12047 2651 12081
rect 2617 11975 2651 12009
rect 2617 11903 2651 11937
rect 2617 11831 2651 11865
rect 2617 11759 2651 11793
rect 2617 11687 2651 11721
rect 2617 11615 2651 11649
rect 2617 11543 2651 11577
rect 2617 11471 2651 11505
rect 2617 11399 2651 11433
rect 2617 11327 2651 11361
rect 2617 11255 2651 11289
rect 2617 11183 2651 11217
rect 2617 11111 2651 11145
rect 2617 11039 2651 11073
rect 2617 10967 2651 11001
rect 2617 10895 2651 10929
rect 2617 10823 2651 10857
rect 2617 10750 2651 10784
rect 2617 10677 2651 10711
rect 2617 10604 2651 10638
rect 2617 10531 2651 10565
rect 2617 10458 2651 10492
rect 2617 10385 2651 10419
rect 2617 10312 2651 10346
rect 2617 10239 2651 10273
rect 2617 10166 2651 10200
rect 2617 10093 2651 10127
rect 2617 10020 2651 10054
rect 2617 9947 2651 9981
rect 2617 9874 2651 9908
rect 2617 9801 2651 9835
rect 2617 9728 2651 9762
rect 2617 9655 2651 9689
rect 2617 9582 2651 9616
rect 2617 9509 2651 9543
rect 2617 9436 2651 9470
rect 2877 10817 3055 13371
rect 2877 10744 2911 10778
rect 2949 10744 2983 10778
rect 3021 10744 3055 10778
rect 2877 10671 2911 10705
rect 2949 10671 2983 10705
rect 3021 10671 3055 10705
rect 2877 10598 2911 10632
rect 2949 10598 2983 10632
rect 3021 10598 3055 10632
rect 2877 10525 2911 10559
rect 2949 10525 2983 10559
rect 3021 10525 3055 10559
rect 2877 10452 2911 10486
rect 2949 10452 2983 10486
rect 3021 10452 3055 10486
rect 2877 10379 2911 10413
rect 2949 10379 2983 10413
rect 3021 10379 3055 10413
rect 2877 10306 2911 10340
rect 2949 10306 2983 10340
rect 3021 10306 3055 10340
rect 2877 10233 2911 10267
rect 2949 10233 2983 10267
rect 3021 10233 3055 10267
rect 2877 10160 2911 10194
rect 2949 10160 2983 10194
rect 3021 10160 3055 10194
rect 2877 10087 2911 10121
rect 2949 10087 2983 10121
rect 3021 10087 3055 10121
rect 2877 10014 2911 10048
rect 2949 10014 2983 10048
rect 3021 10014 3055 10048
rect 2877 9941 2911 9975
rect 2949 9941 2983 9975
rect 3021 9941 3055 9975
rect 2877 9868 2911 9902
rect 2949 9868 2983 9902
rect 3021 9868 3055 9902
rect 2877 9795 2911 9829
rect 2949 9795 2983 9829
rect 3021 9795 3055 9829
rect 2877 9722 2911 9756
rect 2949 9722 2983 9756
rect 3021 9722 3055 9756
rect 2877 9649 2911 9683
rect 2949 9649 2983 9683
rect 3021 9649 3055 9683
rect 2877 9576 2911 9610
rect 2949 9576 2983 9610
rect 3021 9576 3055 9610
rect 2877 9503 2911 9537
rect 2949 9503 2983 9537
rect 3021 9503 3055 9537
rect 3797 10817 3975 13371
rect 3797 10744 3831 10778
rect 3869 10744 3903 10778
rect 3941 10744 3975 10778
rect 3797 10671 3831 10705
rect 3869 10671 3903 10705
rect 3941 10671 3975 10705
rect 3797 10598 3831 10632
rect 3869 10598 3903 10632
rect 3941 10598 3975 10632
rect 3797 10525 3831 10559
rect 3869 10525 3903 10559
rect 3941 10525 3975 10559
rect 3797 10452 3831 10486
rect 3869 10452 3903 10486
rect 3941 10452 3975 10486
rect 3797 10379 3831 10413
rect 3869 10379 3903 10413
rect 3941 10379 3975 10413
rect 3797 10306 3831 10340
rect 3869 10306 3903 10340
rect 3941 10306 3975 10340
rect 3797 10233 3831 10267
rect 3869 10233 3903 10267
rect 3941 10233 3975 10267
rect 3797 10160 3831 10194
rect 3869 10160 3903 10194
rect 3941 10160 3975 10194
rect 3797 10087 3831 10121
rect 3869 10087 3903 10121
rect 3941 10087 3975 10121
rect 3797 10014 3831 10048
rect 3869 10014 3903 10048
rect 3941 10014 3975 10048
rect 3797 9941 3831 9975
rect 3869 9941 3903 9975
rect 3941 9941 3975 9975
rect 3797 9868 3831 9902
rect 3869 9868 3903 9902
rect 3941 9868 3975 9902
rect 3797 9795 3831 9829
rect 3869 9795 3903 9829
rect 3941 9795 3975 9829
rect 3797 9722 3831 9756
rect 3869 9722 3903 9756
rect 3941 9722 3975 9756
rect 3797 9649 3831 9683
rect 3869 9649 3903 9683
rect 3941 9649 3975 9683
rect 3797 9576 3831 9610
rect 3869 9576 3903 9610
rect 3941 9576 3975 9610
rect 3797 9503 3831 9537
rect 3869 9503 3903 9537
rect 3941 9503 3975 9537
rect 4717 10160 4895 13362
rect 4717 10087 4751 10121
rect 4789 10087 4823 10121
rect 4861 10087 4895 10121
rect 4717 10014 4751 10048
rect 4789 10014 4823 10048
rect 4861 10014 4895 10048
rect 4717 9941 4751 9975
rect 4789 9941 4823 9975
rect 4861 9941 4895 9975
rect 4717 9868 4751 9902
rect 4789 9868 4823 9902
rect 4861 9868 4895 9902
rect 4717 9795 4751 9829
rect 4789 9795 4823 9829
rect 4861 9795 4895 9829
rect 4717 9722 4751 9756
rect 4789 9722 4823 9756
rect 4861 9722 4895 9756
rect 4717 9649 4751 9683
rect 4789 9649 4823 9683
rect 4861 9649 4895 9683
rect 4717 9576 4751 9610
rect 4789 9576 4823 9610
rect 4861 9576 4895 9610
rect 4717 9503 4751 9537
rect 4789 9503 4823 9537
rect 4861 9503 4895 9537
rect 5637 10160 5815 13362
rect 5637 10087 5671 10121
rect 5709 10087 5743 10121
rect 5781 10087 5815 10121
rect 5637 10014 5671 10048
rect 5709 10014 5743 10048
rect 5781 10014 5815 10048
rect 5637 9941 5671 9975
rect 5709 9941 5743 9975
rect 5781 9941 5815 9975
rect 5637 9868 5671 9902
rect 5709 9868 5743 9902
rect 5781 9868 5815 9902
rect 5637 9795 5671 9829
rect 5709 9795 5743 9829
rect 5781 9795 5815 9829
rect 5637 9722 5671 9756
rect 5709 9722 5743 9756
rect 5781 9722 5815 9756
rect 5637 9649 5671 9683
rect 5709 9649 5743 9683
rect 5781 9649 5815 9683
rect 5637 9576 5671 9610
rect 5709 9576 5743 9610
rect 5781 9576 5815 9610
rect 5637 9503 5671 9537
rect 5709 9503 5743 9537
rect 5781 9503 5815 9537
rect 6557 10160 6735 13362
rect 6557 10087 6591 10121
rect 6629 10087 6663 10121
rect 6701 10087 6735 10121
rect 6557 10014 6591 10048
rect 6629 10014 6663 10048
rect 6701 10014 6735 10048
rect 6557 9941 6591 9975
rect 6629 9941 6663 9975
rect 6701 9941 6735 9975
rect 6557 9868 6591 9902
rect 6629 9868 6663 9902
rect 6701 9868 6735 9902
rect 6557 9795 6591 9829
rect 6629 9795 6663 9829
rect 6701 9795 6735 9829
rect 6557 9722 6591 9756
rect 6629 9722 6663 9756
rect 6701 9722 6735 9756
rect 6557 9649 6591 9683
rect 6629 9649 6663 9683
rect 6701 9649 6735 9683
rect 6557 9576 6591 9610
rect 6629 9576 6663 9610
rect 6701 9576 6735 9610
rect 6557 9503 6591 9537
rect 6629 9503 6663 9537
rect 6701 9503 6735 9537
rect 7477 10160 7655 13362
rect 7477 10087 7511 10121
rect 7549 10087 7583 10121
rect 7621 10087 7655 10121
rect 7477 10014 7511 10048
rect 7549 10014 7583 10048
rect 7621 10014 7655 10048
rect 7477 9941 7511 9975
rect 7549 9941 7583 9975
rect 7621 9941 7655 9975
rect 7477 9868 7511 9902
rect 7549 9868 7583 9902
rect 7621 9868 7655 9902
rect 7477 9795 7511 9829
rect 7549 9795 7583 9829
rect 7621 9795 7655 9829
rect 7477 9722 7511 9756
rect 7549 9722 7583 9756
rect 7621 9722 7655 9756
rect 7477 9649 7511 9683
rect 7549 9649 7583 9683
rect 7621 9649 7655 9683
rect 7477 9576 7511 9610
rect 7549 9576 7583 9610
rect 7621 9576 7655 9610
rect 7477 9503 7511 9537
rect 7549 9503 7583 9537
rect 7621 9503 7655 9537
rect 8397 10160 8575 13362
rect 8397 10087 8431 10121
rect 8469 10087 8503 10121
rect 8541 10087 8575 10121
rect 8397 10014 8431 10048
rect 8469 10014 8503 10048
rect 8541 10014 8575 10048
rect 8397 9941 8431 9975
rect 8469 9941 8503 9975
rect 8541 9941 8575 9975
rect 8397 9868 8431 9902
rect 8469 9868 8503 9902
rect 8541 9868 8575 9902
rect 8397 9795 8431 9829
rect 8469 9795 8503 9829
rect 8541 9795 8575 9829
rect 8397 9722 8431 9756
rect 8469 9722 8503 9756
rect 8541 9722 8575 9756
rect 8397 9649 8431 9683
rect 8469 9649 8503 9683
rect 8541 9649 8575 9683
rect 8397 9576 8431 9610
rect 8469 9576 8503 9610
rect 8541 9576 8575 9610
rect 8397 9503 8431 9537
rect 8469 9503 8503 9537
rect 8541 9503 8575 9537
rect 9317 10160 9495 13362
rect 9317 10087 9351 10121
rect 9389 10087 9423 10121
rect 9461 10087 9495 10121
rect 9317 10014 9351 10048
rect 9389 10014 9423 10048
rect 9461 10014 9495 10048
rect 9317 9941 9351 9975
rect 9389 9941 9423 9975
rect 9461 9941 9495 9975
rect 9317 9868 9351 9902
rect 9389 9868 9423 9902
rect 9461 9868 9495 9902
rect 9317 9795 9351 9829
rect 9389 9795 9423 9829
rect 9461 9795 9495 9829
rect 9317 9722 9351 9756
rect 9389 9722 9423 9756
rect 9461 9722 9495 9756
rect 9317 9649 9351 9683
rect 9389 9649 9423 9683
rect 9461 9649 9495 9683
rect 9317 9576 9351 9610
rect 9389 9576 9423 9610
rect 9461 9576 9495 9610
rect 9317 9503 9351 9537
rect 9389 9503 9423 9537
rect 9461 9503 9495 9537
rect 10237 10160 10415 13362
rect 10237 10087 10271 10121
rect 10309 10087 10343 10121
rect 10381 10087 10415 10121
rect 10237 10014 10271 10048
rect 10309 10014 10343 10048
rect 10381 10014 10415 10048
rect 10237 9941 10271 9975
rect 10309 9941 10343 9975
rect 10381 9941 10415 9975
rect 10237 9868 10271 9902
rect 10309 9868 10343 9902
rect 10381 9868 10415 9902
rect 10237 9795 10271 9829
rect 10309 9795 10343 9829
rect 10381 9795 10415 9829
rect 10237 9722 10271 9756
rect 10309 9722 10343 9756
rect 10381 9722 10415 9756
rect 10237 9649 10271 9683
rect 10309 9649 10343 9683
rect 10381 9649 10415 9683
rect 10237 9576 10271 9610
rect 10309 9576 10343 9610
rect 10381 9576 10415 9610
rect 10237 9503 10271 9537
rect 10309 9503 10343 9537
rect 10381 9503 10415 9537
rect 11157 10160 11335 13362
rect 11157 10087 11191 10121
rect 11229 10087 11263 10121
rect 11301 10087 11335 10121
rect 11157 10014 11191 10048
rect 11229 10014 11263 10048
rect 11301 10014 11335 10048
rect 11157 9941 11191 9975
rect 11229 9941 11263 9975
rect 11301 9941 11335 9975
rect 11157 9868 11191 9902
rect 11229 9868 11263 9902
rect 11301 9868 11335 9902
rect 11157 9795 11191 9829
rect 11229 9795 11263 9829
rect 11301 9795 11335 9829
rect 11157 9722 11191 9756
rect 11229 9722 11263 9756
rect 11301 9722 11335 9756
rect 11157 9649 11191 9683
rect 11229 9649 11263 9683
rect 11301 9649 11335 9683
rect 11157 9576 11191 9610
rect 11229 9576 11263 9610
rect 11301 9576 11335 9610
rect 11157 9503 11191 9537
rect 11229 9503 11263 9537
rect 11301 9503 11335 9537
rect 12077 10160 12255 13362
rect 12077 10087 12111 10121
rect 12149 10087 12183 10121
rect 12221 10087 12255 10121
rect 12077 10014 12111 10048
rect 12149 10014 12183 10048
rect 12221 10014 12255 10048
rect 12077 9941 12111 9975
rect 12149 9941 12183 9975
rect 12221 9941 12255 9975
rect 12077 9868 12111 9902
rect 12149 9868 12183 9902
rect 12221 9868 12255 9902
rect 12077 9795 12111 9829
rect 12149 9795 12183 9829
rect 12221 9795 12255 9829
rect 12077 9722 12111 9756
rect 12149 9722 12183 9756
rect 12221 9722 12255 9756
rect 12077 9649 12111 9683
rect 12149 9649 12183 9683
rect 12221 9649 12255 9683
rect 12077 9576 12111 9610
rect 12149 9576 12183 9610
rect 12221 9576 12255 9610
rect 12077 9503 12111 9537
rect 12149 9503 12183 9537
rect 12221 9503 12255 9537
rect 12997 10160 13175 13362
rect 12997 10087 13031 10121
rect 13069 10087 13103 10121
rect 13141 10087 13175 10121
rect 12997 10014 13031 10048
rect 13069 10014 13103 10048
rect 13141 10014 13175 10048
rect 12997 9941 13031 9975
rect 13069 9941 13103 9975
rect 13141 9941 13175 9975
rect 12997 9868 13031 9902
rect 13069 9868 13103 9902
rect 13141 9868 13175 9902
rect 12997 9795 13031 9829
rect 13069 9795 13103 9829
rect 13141 9795 13175 9829
rect 12997 9722 13031 9756
rect 13069 9722 13103 9756
rect 13141 9722 13175 9756
rect 12997 9649 13031 9683
rect 13069 9649 13103 9683
rect 13141 9649 13175 9683
rect 12997 9576 13031 9610
rect 13069 9576 13103 9610
rect 13141 9576 13175 9610
rect 12997 9503 13031 9537
rect 13069 9503 13103 9537
rect 13141 9503 13175 9537
rect 2617 9363 2651 9397
rect 2697 9357 2731 9391
rect 2770 9357 2804 9391
rect 2843 9357 2877 9391
rect 2916 9357 2950 9391
rect 2989 9357 3023 9391
rect 3061 9357 3095 9391
rect 3133 9357 3167 9391
rect 3205 9364 3210 9391
rect 3210 9364 3239 9391
rect 3277 9364 3278 9391
rect 3278 9364 3311 9391
rect 3205 9357 3239 9364
rect 3277 9357 3311 9364
rect 3349 9357 3383 9391
rect 3421 9357 3455 9391
rect 3493 9357 3527 9391
rect 3565 9364 3578 9391
rect 3578 9364 3599 9391
rect 3637 9364 3646 9391
rect 3646 9364 3671 9391
rect 3565 9357 3599 9364
rect 3637 9357 3671 9364
rect 3709 9357 3743 9391
rect 3781 9357 3815 9391
rect 3853 9357 3887 9391
rect 3925 9357 3959 9391
rect 3997 9357 4031 9391
rect 4069 9364 4096 9391
rect 4096 9364 4103 9391
rect 4141 9364 4164 9391
rect 4164 9364 4175 9391
rect 4069 9357 4103 9364
rect 4141 9357 4175 9364
rect 4213 9357 4247 9391
rect 4285 9357 4319 9391
rect 4357 9357 4391 9391
rect 4429 9357 4463 9391
rect 4501 9364 4532 9391
rect 4532 9364 4535 9391
rect 4573 9364 4600 9391
rect 4600 9364 4607 9391
rect 4501 9357 4535 9364
rect 4573 9357 4607 9364
rect 4645 9357 4679 9391
rect 4717 9357 4751 9391
rect 4789 9357 4823 9391
rect 4861 9357 4895 9391
rect 4933 9357 4967 9391
rect 5005 9364 5016 9391
rect 5016 9364 5039 9391
rect 5077 9364 5084 9391
rect 5084 9364 5111 9391
rect 5005 9357 5039 9364
rect 5077 9357 5111 9364
rect 5149 9357 5183 9391
rect 5221 9357 5255 9391
rect 5293 9357 5327 9391
rect 5365 9357 5399 9391
rect 5437 9364 5452 9391
rect 5452 9364 5471 9391
rect 5509 9364 5520 9391
rect 5520 9364 5543 9391
rect 5437 9357 5471 9364
rect 5509 9357 5543 9364
rect 5581 9357 5615 9391
rect 5653 9357 5687 9391
rect 5725 9357 5759 9391
rect 5797 9357 5831 9391
rect 5869 9357 5903 9391
rect 5941 9364 5970 9391
rect 5970 9364 5975 9391
rect 6013 9364 6038 9391
rect 6038 9364 6047 9391
rect 5941 9357 5975 9364
rect 6013 9357 6047 9364
rect 6085 9357 6119 9391
rect 6157 9357 6191 9391
rect 6229 9357 6263 9391
rect 6301 9357 6335 9391
rect 6373 9364 6406 9391
rect 6406 9364 6407 9391
rect 6373 9357 6407 9364
rect 6445 9357 6479 9391
rect 6517 9357 6551 9391
rect 6589 9357 6623 9391
rect 6661 9357 6695 9391
rect 6733 9357 6767 9391
rect 6805 9357 6839 9391
rect 6877 9364 6890 9391
rect 6890 9364 6911 9391
rect 6949 9364 6958 9391
rect 6958 9364 6983 9391
rect 6877 9357 6911 9364
rect 6949 9357 6983 9364
rect 7021 9357 7055 9391
rect 7093 9357 7127 9391
rect 7165 9357 7199 9391
rect 7237 9364 7258 9391
rect 7258 9364 7271 9391
rect 7309 9364 7326 9391
rect 7326 9364 7343 9391
rect 7237 9357 7271 9364
rect 7309 9357 7343 9364
rect 7381 9357 7415 9391
rect 7453 9357 7487 9391
rect 7525 9357 7559 9391
rect 7597 9357 7631 9391
rect 7669 9357 7703 9391
rect 7741 9357 7775 9391
rect 7813 9364 7844 9391
rect 7844 9364 7847 9391
rect 7813 9357 7847 9364
rect 7885 9357 7919 9391
rect 7957 9357 7991 9391
rect 8029 9357 8063 9391
rect 8101 9357 8135 9391
rect 8173 9364 8178 9391
rect 8178 9364 8207 9391
rect 8245 9364 8246 9391
rect 8246 9364 8279 9391
rect 8173 9357 8207 9364
rect 8245 9357 8279 9364
rect 8317 9357 8351 9391
rect 8389 9357 8423 9391
rect 8461 9357 8495 9391
rect 8533 9357 8567 9391
rect 8605 9357 8639 9391
rect 8677 9364 8696 9391
rect 8696 9364 8711 9391
rect 8749 9364 8764 9391
rect 8764 9364 8783 9391
rect 8677 9357 8711 9364
rect 8749 9357 8783 9364
rect 8821 9357 8855 9391
rect 8893 9357 8927 9391
rect 8965 9357 8999 9391
rect 9037 9357 9071 9391
rect 9109 9364 9132 9391
rect 9132 9364 9143 9391
rect 9181 9364 9200 9391
rect 9200 9364 9215 9391
rect 9109 9357 9143 9364
rect 9181 9357 9215 9364
rect 9253 9357 9287 9391
rect 9325 9357 9359 9391
rect 9397 9357 9431 9391
rect 9469 9357 9503 9391
rect 9541 9357 9575 9391
rect 9613 9364 9616 9391
rect 9616 9364 9647 9391
rect 9685 9364 9718 9391
rect 9718 9364 9719 9391
rect 9613 9357 9647 9364
rect 9685 9357 9719 9364
rect 9757 9357 9791 9391
rect 9829 9357 9863 9391
rect 9901 9357 9935 9391
rect 9973 9357 10007 9391
rect 10045 9364 10052 9391
rect 10052 9364 10079 9391
rect 10117 9364 10120 9391
rect 10120 9364 10151 9391
rect 10045 9357 10079 9364
rect 10117 9357 10151 9364
rect 10189 9357 10223 9391
rect 10261 9357 10295 9391
rect 10333 9357 10367 9391
rect 10405 9357 10439 9391
rect 10477 9357 10511 9391
rect 10549 9364 10570 9391
rect 10570 9364 10583 9391
rect 10621 9364 10638 9391
rect 10638 9364 10655 9391
rect 10549 9357 10583 9364
rect 10621 9357 10655 9364
rect 10693 9357 10727 9391
rect 10765 9357 10799 9391
rect 10837 9357 10871 9391
rect 10909 9364 10938 9391
rect 10938 9364 10943 9391
rect 10981 9364 11006 9391
rect 11006 9364 11015 9391
rect 10909 9357 10943 9364
rect 10981 9357 11015 9364
rect 11053 9357 11087 9391
rect 11125 9357 11159 9391
rect 11197 9357 11231 9391
rect 11269 9357 11303 9391
rect 11341 9357 11375 9391
rect 11413 9357 11447 9391
rect 11485 9364 11490 9391
rect 11490 9364 11519 9391
rect 11557 9364 11558 9391
rect 11558 9364 11591 9391
rect 11485 9357 11519 9364
rect 11557 9357 11591 9364
rect 11629 9357 11663 9391
rect 11701 9357 11735 9391
rect 11773 9357 11807 9391
rect 11845 9364 11858 9391
rect 11858 9364 11879 9391
rect 11917 9364 11926 9391
rect 11926 9364 11951 9391
rect 11845 9357 11879 9364
rect 11917 9357 11951 9364
rect 11989 9357 12023 9391
rect 12061 9357 12095 9391
rect 12133 9357 12167 9391
rect 12205 9357 12239 9391
rect 12277 9357 12311 9391
rect 12349 9364 12376 9391
rect 12376 9364 12383 9391
rect 12421 9364 12444 9391
rect 12444 9364 12455 9391
rect 12349 9357 12383 9364
rect 12421 9357 12455 9364
rect 12493 9357 12527 9391
rect 12565 9357 12599 9391
rect 12637 9357 12671 9391
rect 12709 9357 12743 9391
rect 12781 9364 12812 9391
rect 12812 9364 12815 9391
rect 12853 9364 12880 9391
rect 12880 9364 12887 9391
rect 12781 9357 12815 9364
rect 12853 9357 12887 9364
rect 2365 9313 2395 9343
rect 2395 9313 2399 9343
rect 2365 9309 2399 9313
rect 2221 9245 2225 9271
rect 2225 9245 2255 9271
rect 2293 9245 2327 9271
rect 13453 9270 13458 16686
rect 2365 9266 13458 9270
rect 2221 9237 2255 9245
rect 2293 9237 2327 9245
rect 2365 9198 13411 9266
rect 13411 9232 13458 9266
rect 13458 9232 13628 16686
rect 13411 9198 13526 9232
rect 2221 9177 2225 9198
rect 2225 9177 2255 9198
rect 2221 9164 2255 9177
rect 2293 9096 13479 9198
rect 13479 9164 13526 9198
rect 13526 9164 13628 9232
rect 13628 9164 13631 16686
rect 13479 9130 13559 9164
rect 13479 9096 13513 9130
rect 13513 9096 13547 9130
rect 13547 9096 13559 9130
rect 2293 9092 13559 9096
rect 13775 9165 13781 28423
rect 13781 9165 14019 28423
rect 14019 9165 14025 28423
rect 1827 8992 1834 9026
rect 1834 8992 1861 9026
rect 1899 8992 1933 9026
rect 1971 9012 2005 9025
rect 2043 9012 2072 9024
rect 2072 9012 2077 9024
rect 1971 8991 2004 9012
rect 2004 8991 2005 9012
rect 2043 8990 2077 9012
rect 1827 8919 1834 8953
rect 1834 8919 1861 8953
rect 1899 8919 1933 8953
rect 1971 8944 2004 8952
rect 2004 8944 2005 8952
rect 13775 9082 13781 9116
rect 13781 9082 13809 9116
rect 13847 9085 13881 9119
rect 13919 9087 13953 9121
rect 13991 9087 14019 9121
rect 14019 9087 14025 9121
rect 13775 8999 13781 9033
rect 13781 8999 13809 9033
rect 13847 9005 13881 9039
rect 13919 9009 13953 9043
rect 13991 9009 14019 9043
rect 14019 9009 14025 9043
rect 1971 8918 2005 8944
rect 2043 8940 8845 8951
rect 8884 8940 8918 8951
rect 8957 8940 8991 8951
rect 9030 8940 9064 8951
rect 9103 8940 9137 8951
rect 9176 8940 9210 8951
rect 9249 8940 9283 8951
rect 9322 8940 9356 8951
rect 9395 8940 9429 8951
rect 9468 8940 9502 8951
rect 9541 8940 9575 8951
rect 9614 8940 9648 8951
rect 9687 8940 9721 8951
rect 9760 8940 9794 8951
rect 9833 8940 9867 8951
rect 9906 8940 9940 8951
rect 9979 8940 10013 8951
rect 10052 8940 10086 8951
rect 10125 8940 10159 8951
rect 10198 8940 10232 8951
rect 10271 8940 10305 8951
rect 10344 8940 10378 8951
rect 10417 8940 10451 8951
rect 10490 8940 10524 8951
rect 10563 8940 10597 8951
rect 10636 8940 10670 8951
rect 10709 8940 10743 8951
rect 10782 8940 10816 8951
rect 10855 8940 10889 8951
rect 10928 8940 10962 8951
rect 11001 8940 11035 8951
rect 11074 8940 11108 8951
rect 11147 8940 11181 8951
rect 11220 8940 11254 8951
rect 11293 8940 11327 8951
rect 11366 8940 11400 8951
rect 11439 8940 11473 8951
rect 11512 8940 11546 8951
rect 11585 8940 11619 8951
rect 11658 8940 11692 8951
rect 11731 8940 11765 8951
rect 11804 8940 11838 8951
rect 11877 8940 11911 8951
rect 11950 8940 11984 8951
rect 12023 8940 12057 8951
rect 12096 8940 12130 8951
rect 12169 8940 12203 8951
rect 12242 8940 12276 8951
rect 12315 8940 12349 8951
rect 12388 8940 12422 8951
rect 12461 8940 12495 8951
rect 12534 8940 12568 8951
rect 12607 8940 12641 8951
rect 12680 8940 12714 8951
rect 12753 8940 12787 8951
rect 12826 8940 12860 8951
rect 12899 8940 12933 8951
rect 12972 8940 13006 8951
rect 13045 8940 13079 8951
rect 13118 8940 13152 8951
rect 13191 8940 13225 8951
rect 13264 8940 13298 8951
rect 13337 8940 13371 8951
rect 13410 8940 13444 8951
rect 13483 8940 13517 8951
rect 13556 8940 13590 8951
rect 13629 8940 13663 8951
rect 1827 8876 1834 8880
rect 1834 8876 1861 8880
rect 1899 8876 1933 8880
rect 2043 8879 8845 8940
rect 8884 8917 8918 8940
rect 8957 8917 8991 8940
rect 9030 8917 9064 8940
rect 9103 8917 9137 8940
rect 9176 8917 9210 8940
rect 9249 8917 9283 8940
rect 9322 8917 9356 8940
rect 9395 8917 9429 8940
rect 9468 8917 9502 8940
rect 9541 8917 9575 8940
rect 9614 8917 9648 8940
rect 9687 8917 9721 8940
rect 9760 8917 9794 8940
rect 9833 8917 9867 8940
rect 9906 8917 9940 8940
rect 9979 8917 10013 8940
rect 10052 8917 10086 8940
rect 10125 8917 10159 8940
rect 10198 8917 10232 8940
rect 10271 8917 10305 8940
rect 10344 8917 10378 8940
rect 10417 8917 10451 8940
rect 10490 8917 10524 8940
rect 10563 8917 10597 8940
rect 10636 8917 10670 8940
rect 10709 8917 10743 8940
rect 10782 8917 10816 8940
rect 10855 8917 10889 8940
rect 10928 8917 10962 8940
rect 11001 8917 11035 8940
rect 11074 8917 11108 8940
rect 11147 8917 11181 8940
rect 11220 8917 11254 8940
rect 11293 8917 11327 8940
rect 11366 8917 11400 8940
rect 11439 8917 11473 8940
rect 11512 8917 11546 8940
rect 11585 8917 11619 8940
rect 11658 8917 11692 8940
rect 11731 8917 11765 8940
rect 11804 8917 11838 8940
rect 11877 8917 11911 8940
rect 11950 8917 11984 8940
rect 12023 8917 12057 8940
rect 12096 8917 12130 8940
rect 12169 8917 12203 8940
rect 12242 8917 12276 8940
rect 12315 8917 12349 8940
rect 12388 8917 12422 8940
rect 12461 8917 12495 8940
rect 12534 8917 12568 8940
rect 12607 8917 12641 8940
rect 12680 8917 12714 8940
rect 12753 8917 12787 8940
rect 12826 8917 12860 8940
rect 12899 8917 12933 8940
rect 12972 8917 13006 8940
rect 13045 8917 13079 8940
rect 13118 8917 13152 8940
rect 13191 8917 13225 8940
rect 13264 8917 13298 8940
rect 13337 8917 13371 8940
rect 13410 8917 13444 8940
rect 13483 8917 13517 8940
rect 13556 8917 13590 8940
rect 13629 8917 13663 8940
rect 13702 8917 13736 8951
rect 13775 8917 13781 8951
rect 13781 8917 13809 8951
rect 13847 8925 13881 8959
rect 13919 8932 13953 8966
rect 13991 8932 14019 8966
rect 14019 8932 14025 8966
rect 1827 8846 1861 8876
rect 1899 8846 1933 8876
rect 1971 8872 2038 8879
rect 2038 8872 8917 8879
rect 1971 8807 8917 8872
rect 8956 8845 8990 8879
rect 9029 8845 9063 8879
rect 9102 8845 9136 8879
rect 9175 8845 9209 8879
rect 9248 8845 9282 8879
rect 9321 8845 9355 8879
rect 9394 8845 9428 8879
rect 9467 8845 9501 8879
rect 9540 8845 9574 8879
rect 9613 8845 9647 8879
rect 9686 8845 9720 8879
rect 9759 8845 9793 8879
rect 9832 8845 9866 8879
rect 9905 8845 9939 8879
rect 9978 8845 10012 8879
rect 10051 8845 10085 8879
rect 10124 8845 10158 8879
rect 10197 8845 10231 8879
rect 10270 8845 10304 8879
rect 10343 8845 10377 8879
rect 10416 8845 10450 8879
rect 10489 8845 10523 8879
rect 10562 8845 10596 8879
rect 10635 8845 10669 8879
rect 10708 8845 10742 8879
rect 10781 8845 10815 8879
rect 10854 8845 10888 8879
rect 10927 8845 10961 8879
rect 11000 8845 11034 8879
rect 11073 8845 11107 8879
rect 11146 8845 11180 8879
rect 11219 8845 11253 8879
rect 11292 8845 11326 8879
rect 11365 8845 11399 8879
rect 11438 8845 11472 8879
rect 11511 8845 11545 8879
rect 11584 8845 11618 8879
rect 11657 8845 11691 8879
rect 11730 8845 11764 8879
rect 11803 8845 11837 8879
rect 11876 8845 11910 8879
rect 11949 8845 11983 8879
rect 12022 8845 12056 8879
rect 12095 8845 12129 8879
rect 12168 8845 12202 8879
rect 12241 8845 12275 8879
rect 12314 8845 12348 8879
rect 12387 8845 12421 8879
rect 12460 8845 12494 8879
rect 12533 8845 12567 8879
rect 12606 8845 12640 8879
rect 12679 8845 12713 8879
rect 12752 8845 12786 8879
rect 12825 8845 12859 8879
rect 12898 8845 12932 8879
rect 12971 8845 13005 8879
rect 13044 8845 13078 8879
rect 13117 8845 13151 8879
rect 13190 8845 13224 8879
rect 13263 8845 13297 8879
rect 13336 8845 13370 8879
rect 13409 8845 13443 8879
rect 13482 8845 13516 8879
rect 13555 8845 13589 8879
rect 13628 8845 13662 8879
rect 13701 8872 13735 8879
rect 13701 8845 13735 8872
rect 13774 8845 13808 8879
rect 13847 8845 13849 8879
rect 13849 8845 13881 8879
rect 13919 8855 13953 8889
rect 13991 8855 14019 8889
rect 14019 8855 14025 8889
rect 1827 8773 1861 8807
rect 1899 8804 1970 8807
rect 1970 8804 8989 8807
rect 229 8728 263 8762
rect 1899 8702 1902 8804
rect 1902 8702 8989 8804
rect 9028 8773 9062 8807
rect 9101 8773 9135 8807
rect 9174 8773 9208 8807
rect 9247 8773 9281 8807
rect 9320 8773 9354 8807
rect 9393 8773 9427 8807
rect 9466 8773 9500 8807
rect 9539 8773 9573 8807
rect 9612 8773 9646 8807
rect 9685 8773 9719 8807
rect 9758 8773 9792 8807
rect 9831 8773 9865 8807
rect 9904 8773 9938 8807
rect 9977 8773 10011 8807
rect 10050 8773 10084 8807
rect 10123 8773 10157 8807
rect 10196 8773 10230 8807
rect 10269 8773 10303 8807
rect 10342 8773 10376 8807
rect 10415 8773 10449 8807
rect 10488 8773 10522 8807
rect 10561 8773 10595 8807
rect 10634 8773 10668 8807
rect 10707 8773 10741 8807
rect 10780 8773 10814 8807
rect 10853 8773 10887 8807
rect 10926 8773 10960 8807
rect 10999 8773 11033 8807
rect 11072 8773 11106 8807
rect 11145 8773 11179 8807
rect 11218 8773 11252 8807
rect 11291 8773 11325 8807
rect 11364 8773 11398 8807
rect 11437 8773 11471 8807
rect 11510 8773 11544 8807
rect 11583 8773 11617 8807
rect 11656 8773 11690 8807
rect 11729 8773 11763 8807
rect 11802 8773 11836 8807
rect 11875 8773 11909 8807
rect 11948 8773 11982 8807
rect 12021 8773 12055 8807
rect 12094 8773 12128 8807
rect 12167 8773 12201 8807
rect 12240 8773 12274 8807
rect 12313 8773 12347 8807
rect 12386 8773 12420 8807
rect 12459 8773 12493 8807
rect 12532 8773 12566 8807
rect 12605 8773 12639 8807
rect 12678 8773 12712 8807
rect 12751 8773 12785 8807
rect 12824 8773 12858 8807
rect 12897 8773 12931 8807
rect 12970 8773 13004 8807
rect 13043 8773 13077 8807
rect 13116 8773 13150 8807
rect 13189 8773 13223 8807
rect 13262 8773 13296 8807
rect 13335 8773 13369 8807
rect 13408 8773 13442 8807
rect 13481 8773 13515 8807
rect 13554 8773 13588 8807
rect 13627 8773 13661 8807
rect 13700 8773 13734 8807
rect 13773 8804 13807 8807
rect 13773 8773 13807 8804
rect 13846 8773 13880 8807
rect 13919 8773 13953 8807
rect 13991 8778 14019 8812
rect 14019 8778 14025 8812
rect 9028 8702 9062 8735
rect 9101 8702 9135 8735
rect 9174 8702 9208 8735
rect 9247 8702 9281 8735
rect 9320 8702 9354 8735
rect 9393 8702 9427 8735
rect 9466 8702 9500 8735
rect 9539 8702 9573 8735
rect 9612 8702 9646 8735
rect 9685 8702 9719 8735
rect 9758 8702 9792 8735
rect 9831 8702 9865 8735
rect 9904 8702 9938 8735
rect 9977 8702 10011 8735
rect 10050 8702 10084 8735
rect 10123 8702 10157 8735
rect 10196 8702 10230 8735
rect 10269 8702 10303 8735
rect 10342 8702 10376 8735
rect 10415 8702 10449 8735
rect 10488 8702 10522 8735
rect 10561 8702 10595 8735
rect 10634 8702 10668 8735
rect 10707 8702 10741 8735
rect 10780 8702 10814 8735
rect 10853 8702 10887 8735
rect 10926 8702 10960 8735
rect 10999 8702 11033 8735
rect 11072 8702 11106 8735
rect 11145 8702 11179 8735
rect 11218 8702 11252 8735
rect 11291 8702 11325 8735
rect 11364 8702 11398 8735
rect 11437 8702 11471 8735
rect 11510 8702 11544 8735
rect 11583 8702 11617 8735
rect 11656 8702 11690 8735
rect 11729 8702 11763 8735
rect 11802 8702 11836 8735
rect 11875 8702 11909 8735
rect 11948 8702 11982 8735
rect 12021 8702 12055 8735
rect 12094 8702 12128 8735
rect 12167 8702 12201 8735
rect 12240 8702 12274 8735
rect 12313 8702 12347 8735
rect 12386 8702 12420 8735
rect 12459 8702 12493 8735
rect 12532 8702 12566 8735
rect 12605 8702 12639 8735
rect 12678 8702 12712 8735
rect 12751 8702 12785 8735
rect 12824 8702 12858 8735
rect 12897 8702 12931 8735
rect 12970 8702 13004 8735
rect 13043 8702 13077 8735
rect 13116 8702 13150 8735
rect 13189 8702 13223 8735
rect 13262 8702 13296 8735
rect 13335 8702 13369 8735
rect 13408 8702 13442 8735
rect 13481 8702 13515 8735
rect 13554 8702 13588 8735
rect 13627 8702 13661 8735
rect 13700 8702 13734 8735
rect 13773 8702 13807 8735
rect 13846 8702 13870 8735
rect 13870 8702 13880 8735
rect 1899 8701 8989 8702
rect 9028 8701 9062 8702
rect 9101 8701 9135 8702
rect 9174 8701 9208 8702
rect 9247 8701 9281 8702
rect 9320 8701 9354 8702
rect 9393 8701 9427 8702
rect 9466 8701 9500 8702
rect 9539 8701 9573 8702
rect 9612 8701 9646 8702
rect 9685 8701 9719 8702
rect 9758 8701 9792 8702
rect 9831 8701 9865 8702
rect 9904 8701 9938 8702
rect 9977 8701 10011 8702
rect 10050 8701 10084 8702
rect 10123 8701 10157 8702
rect 10196 8701 10230 8702
rect 10269 8701 10303 8702
rect 10342 8701 10376 8702
rect 10415 8701 10449 8702
rect 10488 8701 10522 8702
rect 10561 8701 10595 8702
rect 10634 8701 10668 8702
rect 10707 8701 10741 8702
rect 10780 8701 10814 8702
rect 10853 8701 10887 8702
rect 10926 8701 10960 8702
rect 10999 8701 11033 8702
rect 11072 8701 11106 8702
rect 11145 8701 11179 8702
rect 11218 8701 11252 8702
rect 11291 8701 11325 8702
rect 11364 8701 11398 8702
rect 11437 8701 11471 8702
rect 11510 8701 11544 8702
rect 11583 8701 11617 8702
rect 11656 8701 11690 8702
rect 11729 8701 11763 8702
rect 11802 8701 11836 8702
rect 11875 8701 11909 8702
rect 11948 8701 11982 8702
rect 12021 8701 12055 8702
rect 12094 8701 12128 8702
rect 12167 8701 12201 8702
rect 12240 8701 12274 8702
rect 12313 8701 12347 8702
rect 12386 8701 12420 8702
rect 12459 8701 12493 8702
rect 12532 8701 12566 8702
rect 12605 8701 12639 8702
rect 12678 8701 12712 8702
rect 12751 8701 12785 8702
rect 12824 8701 12858 8702
rect 12897 8701 12931 8702
rect 12970 8701 13004 8702
rect 13043 8701 13077 8702
rect 13116 8701 13150 8702
rect 13189 8701 13223 8702
rect 13262 8701 13296 8702
rect 13335 8701 13369 8702
rect 13408 8701 13442 8702
rect 13481 8701 13515 8702
rect 13554 8701 13588 8702
rect 13627 8701 13661 8702
rect 13700 8701 13734 8702
rect 13773 8701 13807 8702
rect 13846 8701 13880 8702
rect 13919 8701 13953 8735
rect 229 8656 263 8690
rect 1610 8654 1644 8688
rect 1682 8654 1716 8688
rect 14094 8564 14128 8598
rect 14166 8564 14200 8598
rect 10536 8465 10570 8499
rect 10609 8465 10643 8499
rect 10682 8465 10716 8499
rect 10755 8465 10789 8499
rect 10828 8465 10862 8499
rect 10901 8465 10935 8499
rect 10974 8465 11008 8499
rect 11047 8465 11081 8499
rect 11120 8465 11154 8499
rect 11193 8465 11227 8499
rect 11266 8465 11300 8499
rect 11339 8465 11373 8499
rect 11412 8465 11446 8499
rect 11485 8465 11519 8499
rect 11558 8465 11592 8499
rect 11631 8465 11665 8499
rect 11704 8465 11738 8499
rect 11777 8465 11811 8499
rect 11850 8465 11884 8499
rect 11923 8465 11957 8499
rect 11996 8465 12030 8499
rect 12069 8465 12103 8499
rect 12142 8465 12176 8499
rect 12215 8465 12249 8499
rect 12288 8465 12322 8499
rect 12361 8465 12395 8499
rect 12434 8465 12468 8499
rect 12507 8465 12541 8499
rect 12580 8465 12614 8499
rect 12653 8465 12687 8499
rect 12726 8465 12760 8499
rect 12799 8465 12833 8499
rect 12872 8465 12906 8499
rect 12945 8465 12979 8499
rect 13018 8465 13052 8499
rect 13091 8457 13701 8499
rect 10464 8392 10498 8426
rect 10536 8393 10570 8427
rect 10609 8423 10638 8427
rect 10638 8423 10643 8427
rect 10682 8423 10706 8427
rect 10706 8423 10716 8427
rect 10755 8423 10774 8427
rect 10774 8423 10789 8427
rect 10828 8423 10842 8427
rect 10842 8423 10862 8427
rect 10901 8423 10910 8427
rect 10910 8423 10935 8427
rect 10974 8423 10978 8427
rect 10978 8423 11008 8427
rect 11047 8423 11080 8427
rect 11080 8423 11081 8427
rect 11120 8423 11148 8427
rect 11148 8423 11154 8427
rect 11193 8423 11216 8427
rect 11216 8423 11227 8427
rect 11266 8423 11284 8427
rect 11284 8423 11300 8427
rect 11339 8423 11352 8427
rect 11352 8423 11373 8427
rect 11412 8423 11420 8427
rect 11420 8423 11446 8427
rect 11485 8423 11488 8427
rect 11488 8423 11519 8427
rect 11558 8423 11590 8427
rect 11590 8423 11592 8427
rect 11631 8423 11658 8427
rect 11658 8423 11665 8427
rect 11704 8423 11726 8427
rect 11726 8423 11738 8427
rect 11777 8423 11794 8427
rect 11794 8423 11811 8427
rect 11850 8423 11862 8427
rect 11862 8423 11884 8427
rect 11923 8423 11930 8427
rect 11930 8423 11957 8427
rect 11996 8423 11998 8427
rect 11998 8423 12030 8427
rect 12069 8423 12100 8427
rect 12100 8423 12103 8427
rect 12142 8423 12168 8427
rect 12168 8423 12176 8427
rect 12215 8423 12236 8427
rect 12236 8423 12249 8427
rect 12288 8423 12304 8427
rect 12304 8423 12322 8427
rect 12361 8423 12372 8427
rect 12372 8423 12395 8427
rect 12434 8423 12440 8427
rect 12440 8423 12468 8427
rect 12507 8423 12508 8427
rect 12508 8423 12541 8427
rect 12580 8423 12610 8427
rect 12610 8423 12614 8427
rect 12653 8423 12678 8427
rect 12678 8423 12687 8427
rect 12726 8423 12746 8427
rect 12746 8423 12760 8427
rect 12799 8423 12814 8427
rect 12814 8423 12833 8427
rect 12872 8423 12882 8427
rect 12882 8423 12906 8427
rect 12945 8423 12950 8427
rect 12950 8423 12979 8427
rect 10609 8393 10643 8423
rect 10682 8393 10716 8423
rect 10755 8393 10789 8423
rect 10828 8393 10862 8423
rect 10901 8393 10935 8423
rect 10974 8393 11008 8423
rect 11047 8393 11081 8423
rect 11120 8393 11154 8423
rect 11193 8393 11227 8423
rect 11266 8393 11300 8423
rect 11339 8393 11373 8423
rect 11412 8393 11446 8423
rect 11485 8393 11519 8423
rect 11558 8393 11592 8423
rect 11631 8393 11665 8423
rect 11704 8393 11738 8423
rect 11777 8393 11811 8423
rect 11850 8393 11884 8423
rect 11923 8393 11957 8423
rect 11996 8393 12030 8423
rect 12069 8393 12103 8423
rect 12142 8393 12176 8423
rect 12215 8393 12249 8423
rect 12288 8393 12322 8423
rect 12361 8393 12395 8423
rect 12434 8393 12468 8423
rect 12507 8393 12541 8423
rect 12580 8393 12614 8423
rect 12653 8393 12687 8423
rect 12726 8393 12760 8423
rect 12799 8393 12833 8423
rect 12872 8393 12906 8423
rect 12945 8393 12979 8423
rect 13018 8393 13052 8427
rect 13091 8423 13120 8457
rect 13120 8423 13154 8457
rect 13154 8423 13188 8457
rect 13188 8423 13222 8457
rect 13222 8423 13256 8457
rect 13256 8423 13290 8457
rect 13290 8423 13324 8457
rect 13324 8423 13358 8457
rect 13358 8423 13392 8457
rect 13392 8423 13426 8457
rect 13426 8423 13460 8457
rect 13460 8423 13494 8457
rect 13494 8423 13528 8457
rect 13528 8423 13562 8457
rect 13562 8423 13596 8457
rect 13596 8423 13630 8457
rect 13630 8423 13664 8457
rect 13664 8423 13698 8457
rect 13698 8423 13701 8457
rect 13091 8393 13701 8423
rect 13739 8393 13773 8427
rect 10464 8321 10498 8353
rect 10464 8319 10473 8321
rect 10473 8319 10498 8321
rect 10536 8319 10570 8353
rect 10608 8325 10642 8355
rect 10681 8325 10715 8355
rect 10754 8325 10788 8355
rect 10827 8325 10861 8355
rect 10900 8325 10934 8355
rect 10973 8325 11007 8355
rect 11046 8325 11080 8355
rect 11119 8325 11153 8355
rect 11192 8325 11226 8355
rect 11265 8325 11299 8355
rect 11338 8325 11372 8355
rect 11411 8325 11445 8355
rect 11484 8325 11518 8355
rect 11557 8325 11591 8355
rect 11630 8325 11664 8355
rect 11703 8325 11737 8355
rect 11776 8325 11810 8355
rect 11849 8325 11883 8355
rect 11922 8325 11956 8355
rect 11995 8325 12029 8355
rect 12068 8325 12102 8355
rect 12141 8325 12175 8355
rect 12214 8325 12248 8355
rect 12287 8325 12321 8355
rect 12360 8325 12394 8355
rect 12433 8325 12467 8355
rect 12506 8325 12540 8355
rect 12579 8325 12613 8355
rect 12652 8325 12686 8355
rect 12725 8325 12759 8355
rect 12798 8325 12832 8355
rect 12871 8325 12905 8355
rect 12944 8325 12978 8355
rect 13017 8325 13051 8355
rect 10608 8321 10639 8325
rect 10639 8321 10642 8325
rect 10681 8321 10710 8325
rect 10710 8321 10715 8325
rect 10754 8321 10778 8325
rect 10778 8321 10788 8325
rect 10827 8321 10846 8325
rect 10846 8321 10861 8325
rect 10900 8321 10914 8325
rect 10914 8321 10934 8325
rect 10973 8321 10982 8325
rect 10982 8321 11007 8325
rect 11046 8321 11050 8325
rect 11050 8321 11080 8325
rect 11119 8321 11152 8325
rect 11152 8321 11153 8325
rect 11192 8321 11220 8325
rect 11220 8321 11226 8325
rect 11265 8321 11288 8325
rect 11288 8321 11299 8325
rect 11338 8321 11356 8325
rect 11356 8321 11372 8325
rect 11411 8321 11424 8325
rect 11424 8321 11445 8325
rect 11484 8321 11492 8325
rect 11492 8321 11518 8325
rect 11557 8321 11560 8325
rect 11560 8321 11591 8325
rect 11630 8321 11662 8325
rect 11662 8321 11664 8325
rect 11703 8321 11730 8325
rect 11730 8321 11737 8325
rect 11776 8321 11798 8325
rect 11798 8321 11810 8325
rect 11849 8321 11866 8325
rect 11866 8321 11883 8325
rect 11922 8321 11934 8325
rect 11934 8321 11956 8325
rect 11995 8321 12002 8325
rect 12002 8321 12029 8325
rect 12068 8321 12070 8325
rect 12070 8321 12102 8325
rect 12141 8321 12172 8325
rect 12172 8321 12175 8325
rect 12214 8321 12240 8325
rect 12240 8321 12248 8325
rect 12287 8321 12308 8325
rect 12308 8321 12321 8325
rect 12360 8321 12376 8325
rect 12376 8321 12394 8325
rect 12433 8321 12444 8325
rect 12444 8321 12467 8325
rect 12506 8321 12512 8325
rect 12512 8321 12540 8325
rect 12579 8321 12580 8325
rect 12580 8321 12613 8325
rect 12652 8321 12682 8325
rect 12682 8321 12686 8325
rect 12725 8321 12750 8325
rect 12750 8321 12759 8325
rect 12798 8321 12818 8325
rect 12818 8321 12832 8325
rect 12871 8321 12886 8325
rect 12886 8321 12905 8325
rect 12944 8321 12954 8325
rect 12954 8321 12978 8325
rect 13017 8321 13022 8325
rect 13022 8321 13051 8325
rect 13090 8321 13124 8355
rect 13163 8325 13557 8393
rect 13595 8325 13629 8326
rect 13163 8321 13192 8325
rect 13192 8321 13226 8325
rect 13226 8321 13260 8325
rect 13260 8321 13294 8325
rect 13294 8321 13328 8325
rect 13328 8321 13362 8325
rect 13362 8321 13396 8325
rect 13396 8321 13430 8325
rect 13430 8321 13464 8325
rect 13464 8321 13498 8325
rect 13498 8321 13532 8325
rect 13532 8321 13557 8325
rect 13595 8292 13600 8325
rect 13600 8292 13629 8325
rect 10464 8253 10498 8280
rect 10464 8246 10473 8253
rect 10473 8246 10498 8253
rect 10536 8246 10570 8280
rect 10608 8257 10642 8282
rect 13667 8263 13701 8297
rect 13739 8290 13766 8297
rect 13766 8290 13773 8297
rect 13739 8263 13773 8290
rect 10608 8248 10639 8257
rect 10639 8248 10642 8257
rect 10464 8185 10498 8207
rect 10464 8173 10473 8185
rect 10473 8173 10498 8185
rect 10536 8173 10570 8207
rect 10608 8189 10642 8209
rect 10608 8175 10639 8189
rect 10639 8175 10642 8189
rect 10464 8117 10498 8134
rect 10464 8100 10473 8117
rect 10473 8100 10498 8117
rect 10536 8100 10570 8134
rect 10608 8121 10642 8136
rect 10608 8102 10639 8121
rect 10639 8102 10642 8121
rect 10464 8049 10498 8061
rect 10464 8027 10473 8049
rect 10473 8027 10498 8049
rect 10536 8027 10570 8061
rect 10608 8053 10642 8063
rect 10608 8029 10639 8053
rect 10639 8029 10642 8053
rect 10464 7981 10498 7988
rect 10464 7954 10473 7981
rect 10473 7954 10498 7981
rect 10536 7954 10570 7988
rect 10608 7985 10642 7990
rect 10608 7956 10639 7985
rect 10639 7956 10642 7985
rect 698 7913 732 7917
rect 771 7913 805 7917
rect 844 7913 878 7917
rect 917 7913 951 7917
rect 990 7913 1024 7917
rect 1063 7913 1097 7917
rect 1136 7913 1170 7917
rect 1209 7913 1243 7917
rect 1282 7913 1316 7917
rect 1355 7913 1389 7917
rect 1428 7913 1462 7917
rect 1501 7913 1535 7917
rect 1574 7913 1608 7917
rect 1647 7913 1681 7917
rect 1720 7913 1754 7917
rect 1793 7913 1827 7917
rect 1866 7913 1900 7917
rect 1939 7913 1973 7917
rect 2012 7913 2046 7917
rect 2085 7913 2119 7917
rect 2158 7913 2192 7917
rect 2231 7913 2265 7917
rect 2304 7913 2338 7917
rect 2377 7913 2411 7917
rect 2450 7913 2484 7917
rect 2523 7913 2557 7917
rect 2596 7913 2630 7917
rect 2669 7913 2703 7917
rect 2742 7913 2776 7917
rect 2815 7913 2849 7917
rect 2888 7913 2922 7917
rect 2961 7913 2995 7917
rect 3034 7913 3068 7917
rect 3107 7913 3141 7917
rect 3180 7913 3214 7917
rect 3253 7913 3287 7917
rect 3326 7913 3360 7917
rect 3399 7913 3433 7917
rect 3472 7913 3506 7917
rect 3545 7913 3579 7917
rect 3618 7913 3652 7917
rect 3691 7913 3725 7917
rect 3764 7913 3798 7917
rect 3837 7913 3871 7917
rect 3910 7913 3944 7917
rect 3983 7913 4017 7917
rect 4056 7913 4090 7917
rect 4129 7913 4163 7917
rect 4202 7913 4236 7917
rect 4275 7913 4309 7917
rect 4348 7913 4382 7917
rect 4421 7913 4455 7917
rect 4494 7913 9568 7917
rect 698 7883 728 7913
rect 728 7883 732 7913
rect 771 7883 805 7913
rect 844 7883 878 7913
rect 917 7883 951 7913
rect 990 7883 1024 7913
rect 1063 7883 1097 7913
rect 1136 7883 1170 7913
rect 1209 7883 1243 7913
rect 1282 7883 1316 7913
rect 1355 7883 1389 7913
rect 1428 7883 1462 7913
rect 1501 7883 1535 7913
rect 1574 7883 1608 7913
rect 1647 7883 1681 7913
rect 1720 7883 1754 7913
rect 1793 7883 1827 7913
rect 1866 7883 1900 7913
rect 1939 7883 1973 7913
rect 2012 7883 2046 7913
rect 2085 7883 2119 7913
rect 2158 7883 2192 7913
rect 2231 7883 2265 7913
rect 2304 7883 2338 7913
rect 2377 7883 2411 7913
rect 2450 7883 2484 7913
rect 2523 7883 2557 7913
rect 2596 7883 2630 7913
rect 2669 7883 2703 7913
rect 2742 7883 2776 7913
rect 2815 7883 2849 7913
rect 2888 7883 2922 7913
rect 2961 7883 2995 7913
rect 3034 7883 3068 7913
rect 3107 7883 3141 7913
rect 3180 7883 3214 7913
rect 3253 7883 3287 7913
rect 3326 7883 3360 7913
rect 3399 7883 3433 7913
rect 3472 7883 3506 7913
rect 3545 7883 3579 7913
rect 3618 7883 3652 7913
rect 3691 7883 3725 7913
rect 3764 7883 3798 7913
rect 3837 7883 3871 7913
rect 3910 7883 3944 7913
rect 3983 7883 4017 7913
rect 4056 7883 4090 7913
rect 4129 7883 4163 7913
rect 4202 7883 4236 7913
rect 4275 7883 4309 7913
rect 4348 7883 4382 7913
rect 4421 7883 4455 7913
rect 626 7777 722 7845
rect 722 7777 732 7845
rect 771 7811 805 7845
rect 844 7811 878 7845
rect 917 7811 951 7845
rect 990 7811 1024 7845
rect 1063 7811 1097 7845
rect 1136 7811 1170 7845
rect 1209 7811 1243 7845
rect 1282 7811 1316 7845
rect 1355 7811 1389 7845
rect 1428 7811 1462 7845
rect 1501 7811 1535 7845
rect 1574 7811 1608 7845
rect 1647 7811 1681 7845
rect 1720 7811 1754 7845
rect 1793 7811 1827 7845
rect 1866 7811 1900 7845
rect 1939 7811 1973 7845
rect 2012 7811 2046 7845
rect 2085 7811 2119 7845
rect 2158 7811 2192 7845
rect 2231 7811 2265 7845
rect 2304 7811 2338 7845
rect 2377 7811 2411 7845
rect 2450 7811 2484 7845
rect 2523 7811 2557 7845
rect 2596 7811 2630 7845
rect 2669 7811 2703 7845
rect 2742 7811 2776 7845
rect 2815 7811 2849 7845
rect 2888 7811 2922 7845
rect 2961 7811 2995 7845
rect 3034 7811 3068 7845
rect 3107 7811 3141 7845
rect 3180 7811 3214 7845
rect 3253 7811 3287 7845
rect 3326 7811 3360 7845
rect 3399 7811 3433 7845
rect 3472 7811 3506 7845
rect 3545 7811 3579 7845
rect 3618 7811 3652 7845
rect 3691 7811 3725 7845
rect 3764 7811 3798 7845
rect 3837 7811 3871 7845
rect 3910 7811 3944 7845
rect 3983 7811 4017 7845
rect 4056 7811 4090 7845
rect 4129 7811 4163 7845
rect 4202 7811 4236 7845
rect 4275 7811 4309 7845
rect 4348 7811 4382 7845
rect 4421 7811 4455 7845
rect 4494 7811 9568 7913
rect 9606 7811 9640 7845
rect 626 7773 732 7777
rect 626 6083 790 7773
rect 790 6083 804 7773
rect 843 7743 877 7773
rect 916 7743 950 7773
rect 989 7743 1023 7773
rect 1062 7743 1096 7773
rect 1135 7743 1169 7773
rect 1208 7743 1242 7773
rect 1281 7743 1315 7773
rect 1354 7743 1388 7773
rect 1427 7743 1461 7773
rect 1500 7743 1534 7773
rect 1573 7743 1607 7773
rect 1646 7743 1680 7773
rect 1719 7743 1753 7773
rect 1792 7743 1826 7773
rect 1865 7743 1899 7773
rect 1938 7743 1972 7773
rect 2011 7743 2045 7773
rect 2084 7743 2118 7773
rect 2157 7743 2191 7773
rect 2230 7743 2264 7773
rect 2303 7743 2337 7773
rect 2376 7743 2410 7773
rect 2449 7743 2483 7773
rect 2522 7743 2556 7773
rect 2595 7743 2629 7773
rect 2668 7743 2702 7773
rect 2741 7743 2775 7773
rect 2814 7743 2848 7773
rect 2887 7743 2921 7773
rect 2960 7743 2994 7773
rect 3033 7743 3067 7773
rect 3106 7743 3140 7773
rect 3179 7743 3213 7773
rect 3252 7743 3286 7773
rect 3325 7743 3359 7773
rect 3398 7743 3432 7773
rect 3471 7743 3505 7773
rect 3544 7743 3578 7773
rect 3617 7743 3651 7773
rect 3690 7743 3724 7773
rect 3763 7743 3797 7773
rect 3836 7743 3870 7773
rect 3909 7743 3943 7773
rect 3982 7743 4016 7773
rect 4055 7743 4089 7773
rect 4128 7743 4162 7773
rect 4201 7743 4235 7773
rect 4274 7743 4308 7773
rect 4347 7743 4381 7773
rect 4420 7743 4454 7773
rect 4493 7743 4527 7773
rect 4566 7743 9496 7811
rect 843 7739 877 7743
rect 916 7739 950 7743
rect 989 7739 1023 7743
rect 1062 7739 1096 7743
rect 1135 7739 1169 7743
rect 1208 7739 1242 7743
rect 1281 7739 1315 7743
rect 1354 7739 1388 7743
rect 1427 7739 1461 7743
rect 1500 7739 1534 7743
rect 1573 7739 1607 7743
rect 1646 7739 1680 7743
rect 1719 7739 1753 7743
rect 1792 7739 1826 7743
rect 1865 7739 1899 7743
rect 1938 7739 1972 7743
rect 2011 7739 2045 7743
rect 2084 7739 2118 7743
rect 2157 7739 2191 7743
rect 2230 7739 2264 7743
rect 2303 7739 2337 7743
rect 2376 7739 2410 7743
rect 2449 7739 2483 7743
rect 2522 7739 2556 7743
rect 2595 7739 2629 7743
rect 2668 7739 2702 7743
rect 2741 7739 2775 7743
rect 2814 7739 2848 7743
rect 2887 7739 2921 7743
rect 2960 7739 2994 7743
rect 3033 7739 3067 7743
rect 3106 7739 3140 7743
rect 3179 7739 3213 7743
rect 3252 7739 3286 7743
rect 3325 7739 3359 7743
rect 3398 7739 3432 7743
rect 3471 7739 3505 7743
rect 3544 7739 3578 7743
rect 3617 7739 3651 7743
rect 3690 7739 3724 7743
rect 3763 7739 3797 7743
rect 3836 7739 3870 7743
rect 3909 7739 3943 7743
rect 3982 7739 4016 7743
rect 4055 7739 4089 7743
rect 4128 7739 4162 7743
rect 4201 7739 4235 7743
rect 4274 7739 4308 7743
rect 4347 7739 4381 7743
rect 4420 7739 4454 7743
rect 4493 7739 4527 7743
rect 4566 7739 9496 7743
rect 9534 7737 9568 7771
rect 9606 7744 9636 7771
rect 9636 7744 9640 7771
rect 9606 7737 9640 7744
rect 9462 7665 9496 7699
rect 9534 7663 9568 7697
rect 9606 7663 9636 7697
rect 9636 7663 9640 7697
rect 9462 7591 9466 7625
rect 9466 7591 9496 7625
rect 9534 7589 9568 7623
rect 9606 7589 9636 7623
rect 9636 7589 9640 7623
rect 626 6011 732 6083
rect 770 6010 790 6044
rect 790 6010 804 6044
rect 626 5938 660 5972
rect 698 5938 732 5972
rect 770 5937 790 5971
rect 790 5937 804 5971
rect 626 5865 660 5899
rect 698 5865 732 5899
rect 770 5864 790 5898
rect 790 5864 804 5898
rect 626 5792 660 5826
rect 698 5792 732 5826
rect 1019 7485 1053 7519
rect 1091 7485 1093 7519
rect 1093 7485 1125 7519
rect 1163 7485 1195 7519
rect 1195 7485 1197 7519
rect 1235 7485 1263 7519
rect 1263 7485 1269 7519
rect 1307 7485 1331 7519
rect 1331 7485 1341 7519
rect 1379 7485 1399 7519
rect 1399 7485 1413 7519
rect 1451 7485 1467 7519
rect 1467 7485 1485 7519
rect 1523 7485 1535 7519
rect 1535 7485 1557 7519
rect 1595 7485 1603 7519
rect 1603 7485 1629 7519
rect 1667 7485 1671 7519
rect 1671 7485 1701 7519
rect 1739 7485 1773 7519
rect 1811 7485 1841 7519
rect 1841 7485 1845 7519
rect 1883 7485 1909 7519
rect 1909 7485 1917 7519
rect 1955 7485 1977 7519
rect 1977 7485 1989 7519
rect 2027 7485 2045 7519
rect 2045 7485 2061 7519
rect 2099 7485 2113 7519
rect 2113 7485 2133 7519
rect 2171 7485 2181 7519
rect 2181 7485 2205 7519
rect 2243 7485 2249 7519
rect 2249 7485 2277 7519
rect 2315 7485 2317 7519
rect 2317 7485 2349 7519
rect 2387 7485 2419 7519
rect 2419 7485 2421 7519
rect 2459 7485 2487 7519
rect 2487 7485 2493 7519
rect 2531 7485 2555 7519
rect 2555 7485 2565 7519
rect 2603 7485 2623 7519
rect 2623 7485 2637 7519
rect 2675 7485 2691 7519
rect 2691 7485 2709 7519
rect 2747 7485 2759 7519
rect 2759 7485 2781 7519
rect 2819 7485 2827 7519
rect 2827 7485 2853 7519
rect 2891 7485 2895 7519
rect 2895 7485 2925 7519
rect 2963 7485 2997 7519
rect 3035 7485 3065 7519
rect 3065 7485 3069 7519
rect 3107 7485 3133 7519
rect 3133 7485 3141 7519
rect 3179 7485 3201 7519
rect 3201 7485 3213 7519
rect 3251 7485 3269 7519
rect 3269 7485 3285 7519
rect 3323 7485 3337 7519
rect 3337 7485 3357 7519
rect 3395 7485 3405 7519
rect 3405 7485 3429 7519
rect 3467 7485 3473 7519
rect 3473 7485 3501 7519
rect 3539 7485 3541 7519
rect 3541 7485 3573 7519
rect 3611 7485 3643 7519
rect 3643 7485 3645 7519
rect 3683 7485 3711 7519
rect 3711 7485 3717 7519
rect 3755 7485 3779 7519
rect 3779 7485 3789 7519
rect 3827 7485 3847 7519
rect 3847 7485 3861 7519
rect 3899 7485 3915 7519
rect 3915 7485 3933 7519
rect 3971 7485 3983 7519
rect 3983 7485 4005 7519
rect 4043 7485 4051 7519
rect 4051 7485 4077 7519
rect 4115 7485 4119 7519
rect 4119 7485 4149 7519
rect 4187 7485 4221 7519
rect 4259 7485 4289 7519
rect 4289 7485 4293 7519
rect 4331 7485 4357 7519
rect 4357 7485 4365 7519
rect 4403 7485 4425 7519
rect 4425 7485 4437 7519
rect 4475 7485 4493 7519
rect 4493 7485 4509 7519
rect 4547 7485 4561 7519
rect 4561 7485 4581 7519
rect 4619 7485 4629 7519
rect 4629 7485 4653 7519
rect 4691 7485 4697 7519
rect 4697 7485 4725 7519
rect 4763 7485 4765 7519
rect 4765 7485 4797 7519
rect 4835 7485 4867 7519
rect 4867 7485 4869 7519
rect 4907 7485 4935 7519
rect 4935 7485 4941 7519
rect 4979 7485 5003 7519
rect 5003 7485 5013 7519
rect 5051 7485 5071 7519
rect 5071 7485 5085 7519
rect 5123 7485 5139 7519
rect 5139 7485 5157 7519
rect 5195 7485 5207 7519
rect 5207 7485 5229 7519
rect 5267 7485 5275 7519
rect 5275 7485 5301 7519
rect 5339 7485 5343 7519
rect 5343 7485 5373 7519
rect 5411 7485 5445 7519
rect 5483 7485 5513 7519
rect 5513 7485 5517 7519
rect 5555 7485 5581 7519
rect 5581 7485 5589 7519
rect 5627 7485 5649 7519
rect 5649 7485 5661 7519
rect 5699 7485 5717 7519
rect 5717 7485 5733 7519
rect 5771 7485 5785 7519
rect 5785 7485 5805 7519
rect 5843 7485 5853 7519
rect 5853 7485 5877 7519
rect 5915 7485 5921 7519
rect 5921 7485 5949 7519
rect 5987 7485 5989 7519
rect 5989 7485 6021 7519
rect 6059 7485 6091 7519
rect 6091 7485 6093 7519
rect 6131 7485 6159 7519
rect 6159 7485 6165 7519
rect 6203 7485 6227 7519
rect 6227 7485 6237 7519
rect 6275 7485 6295 7519
rect 6295 7485 6309 7519
rect 6347 7485 6363 7519
rect 6363 7485 6381 7519
rect 6419 7485 6431 7519
rect 6431 7485 6453 7519
rect 6491 7485 6499 7519
rect 6499 7485 6525 7519
rect 6563 7485 6567 7519
rect 6567 7485 6597 7519
rect 6635 7485 6669 7519
rect 6707 7485 6737 7519
rect 6737 7485 6741 7519
rect 6779 7485 6805 7519
rect 6805 7485 6813 7519
rect 6851 7485 6873 7519
rect 6873 7485 6885 7519
rect 6923 7485 6941 7519
rect 6941 7485 6957 7519
rect 6995 7485 7009 7519
rect 7009 7485 7029 7519
rect 7067 7485 7077 7519
rect 7077 7485 7101 7519
rect 7139 7485 7145 7519
rect 7145 7485 7173 7519
rect 7211 7485 7213 7519
rect 7213 7485 7245 7519
rect 7283 7485 7315 7519
rect 7315 7485 7317 7519
rect 7355 7485 7383 7519
rect 7383 7485 7389 7519
rect 7427 7485 7451 7519
rect 7451 7485 7461 7519
rect 7499 7485 7519 7519
rect 7519 7485 7533 7519
rect 7571 7485 7587 7519
rect 7587 7485 7605 7519
rect 7643 7485 7655 7519
rect 7655 7485 7677 7519
rect 7715 7485 7723 7519
rect 7723 7485 7749 7519
rect 7787 7485 7791 7519
rect 7791 7485 7821 7519
rect 7859 7485 7893 7519
rect 7931 7485 7961 7519
rect 7961 7485 7965 7519
rect 8003 7485 8029 7519
rect 8029 7485 8037 7519
rect 8075 7485 8097 7519
rect 8097 7485 8109 7519
rect 8147 7485 8165 7519
rect 8165 7485 8181 7519
rect 8219 7485 8233 7519
rect 8233 7485 8253 7519
rect 8291 7485 8301 7519
rect 8301 7485 8325 7519
rect 8363 7485 8369 7519
rect 8369 7485 8397 7519
rect 8435 7485 8437 7519
rect 8437 7485 8469 7519
rect 8507 7485 8539 7519
rect 8539 7485 8541 7519
rect 8579 7485 8607 7519
rect 8607 7485 8613 7519
rect 8651 7485 8675 7519
rect 8675 7485 8685 7519
rect 8723 7485 8743 7519
rect 8743 7485 8757 7519
rect 8795 7485 8811 7519
rect 8811 7485 8829 7519
rect 8867 7485 8879 7519
rect 8879 7485 8901 7519
rect 8939 7485 8947 7519
rect 8947 7485 8973 7519
rect 9012 7485 9015 7519
rect 9015 7485 9046 7519
rect 9085 7485 9117 7519
rect 9117 7485 9119 7519
rect 947 7417 981 7447
rect 947 7413 981 7417
rect 1269 7412 1284 7428
rect 1284 7412 1303 7428
rect 1342 7412 1353 7428
rect 1353 7412 1376 7428
rect 1415 7412 1422 7428
rect 1422 7412 1449 7428
rect 1488 7412 1491 7428
rect 1491 7412 1522 7428
rect 1561 7412 1594 7428
rect 1594 7412 1595 7428
rect 1634 7412 1663 7428
rect 1663 7412 1668 7428
rect 1707 7412 1732 7428
rect 1732 7412 1741 7428
rect 1780 7412 1801 7428
rect 1801 7412 1814 7428
rect 1853 7412 1870 7428
rect 1870 7412 1887 7428
rect 1926 7412 1939 7428
rect 1939 7412 1960 7428
rect 1999 7412 2008 7428
rect 2008 7412 2033 7428
rect 2072 7412 2077 7428
rect 2077 7412 2106 7428
rect 2145 7412 2146 7428
rect 2146 7412 2179 7428
rect 2218 7412 2250 7428
rect 2250 7412 2252 7428
rect 2291 7412 2319 7428
rect 2319 7412 2325 7428
rect 2364 7412 2388 7428
rect 2388 7412 2398 7428
rect 2437 7412 2457 7428
rect 2457 7412 2471 7428
rect 2510 7412 2526 7428
rect 2526 7412 2544 7428
rect 2583 7412 2595 7428
rect 2595 7412 2617 7428
rect 2656 7412 2664 7428
rect 2664 7412 2690 7428
rect 2729 7412 2733 7428
rect 2733 7412 2763 7428
rect 2802 7412 2836 7428
rect 2875 7412 2905 7428
rect 2905 7412 2909 7428
rect 2948 7412 2974 7428
rect 2974 7412 2982 7428
rect 3021 7412 3043 7428
rect 3043 7412 3055 7428
rect 3094 7412 3112 7428
rect 3112 7412 3128 7428
rect 3167 7412 3181 7428
rect 3181 7412 3201 7428
rect 3240 7412 3250 7428
rect 3250 7412 3274 7428
rect 3313 7412 3319 7428
rect 3319 7412 3347 7428
rect 3386 7412 3388 7428
rect 3388 7412 3420 7428
rect 3459 7412 3492 7428
rect 3492 7412 3493 7428
rect 3532 7412 3561 7428
rect 3561 7412 3566 7428
rect 3605 7412 3630 7428
rect 3630 7412 3639 7428
rect 3678 7412 3699 7428
rect 3699 7412 3712 7428
rect 3751 7412 3768 7428
rect 3768 7412 3785 7428
rect 3824 7412 3837 7428
rect 3837 7412 3858 7428
rect 3897 7412 3906 7428
rect 3906 7412 3931 7428
rect 3970 7412 3975 7428
rect 3975 7412 4004 7428
rect 4043 7412 4044 7428
rect 4044 7412 4077 7428
rect 4116 7412 4147 7428
rect 4147 7412 4150 7428
rect 4189 7412 4216 7428
rect 4216 7412 4223 7428
rect 4262 7412 4285 7428
rect 4285 7412 4296 7428
rect 4335 7412 4354 7428
rect 4354 7412 4369 7428
rect 4408 7412 4423 7428
rect 4423 7412 4442 7428
rect 4481 7412 4492 7428
rect 4492 7412 4515 7428
rect 4554 7412 4561 7428
rect 4561 7412 4588 7428
rect 4627 7412 4630 7428
rect 4630 7412 4661 7428
rect 1269 7394 1303 7412
rect 1342 7394 1376 7412
rect 1415 7394 1449 7412
rect 1488 7394 1522 7412
rect 1561 7394 1595 7412
rect 1634 7394 1668 7412
rect 1707 7394 1741 7412
rect 1780 7394 1814 7412
rect 1853 7394 1887 7412
rect 1926 7394 1960 7412
rect 1999 7394 2033 7412
rect 2072 7394 2106 7412
rect 2145 7394 2179 7412
rect 2218 7394 2252 7412
rect 2291 7394 2325 7412
rect 2364 7394 2398 7412
rect 2437 7394 2471 7412
rect 2510 7394 2544 7412
rect 2583 7394 2617 7412
rect 2656 7394 2690 7412
rect 2729 7394 2763 7412
rect 2802 7394 2836 7412
rect 2875 7394 2909 7412
rect 2948 7394 2982 7412
rect 3021 7394 3055 7412
rect 3094 7394 3128 7412
rect 3167 7394 3201 7412
rect 3240 7394 3274 7412
rect 3313 7394 3347 7412
rect 3386 7394 3420 7412
rect 3459 7394 3493 7412
rect 3532 7394 3566 7412
rect 3605 7394 3639 7412
rect 3678 7394 3712 7412
rect 3751 7394 3785 7412
rect 3824 7394 3858 7412
rect 3897 7394 3931 7412
rect 3970 7394 4004 7412
rect 4043 7394 4077 7412
rect 4116 7394 4150 7412
rect 4189 7394 4223 7412
rect 4262 7394 4296 7412
rect 4335 7394 4369 7412
rect 4408 7394 4442 7412
rect 4481 7394 4515 7412
rect 4554 7394 4588 7412
rect 4627 7394 4661 7412
rect 4700 7394 4734 7428
rect 4773 7412 4803 7428
rect 4803 7412 4807 7428
rect 4846 7412 4872 7428
rect 4872 7412 4880 7428
rect 4919 7412 4941 7428
rect 4941 7412 4953 7428
rect 4992 7412 5010 7428
rect 5010 7412 5026 7428
rect 5065 7412 5079 7428
rect 5079 7412 5099 7428
rect 5138 7412 5148 7428
rect 5148 7412 5172 7428
rect 5211 7412 5217 7428
rect 5217 7412 5245 7428
rect 5284 7412 5286 7428
rect 5286 7412 5318 7428
rect 5357 7412 5389 7428
rect 5389 7412 5391 7428
rect 5430 7412 5458 7428
rect 5458 7412 5464 7428
rect 5503 7412 5527 7428
rect 5527 7412 5537 7428
rect 5576 7412 5596 7428
rect 5596 7412 5610 7428
rect 5649 7412 5664 7428
rect 5664 7412 5683 7428
rect 5722 7412 5732 7428
rect 5732 7412 5756 7428
rect 5795 7412 5800 7428
rect 5800 7412 5829 7428
rect 4773 7394 4807 7412
rect 4846 7394 4880 7412
rect 4919 7394 4953 7412
rect 4992 7394 5026 7412
rect 5065 7394 5099 7412
rect 5138 7394 5172 7412
rect 5211 7394 5245 7412
rect 5284 7394 5318 7412
rect 5357 7394 5391 7412
rect 5430 7394 5464 7412
rect 5503 7394 5537 7412
rect 5576 7394 5610 7412
rect 5649 7394 5683 7412
rect 5722 7394 5756 7412
rect 5795 7394 5829 7412
rect 5868 7394 5902 7428
rect 5941 7412 5970 7428
rect 5970 7412 5975 7428
rect 6014 7412 6038 7428
rect 6038 7412 6048 7428
rect 6087 7412 6106 7428
rect 6106 7412 6121 7428
rect 6160 7412 6174 7428
rect 6174 7412 6194 7428
rect 6233 7412 6242 7428
rect 6242 7412 6267 7428
rect 6306 7412 6310 7428
rect 6310 7412 6340 7428
rect 6379 7412 6412 7428
rect 6412 7412 6413 7428
rect 6451 7412 6480 7428
rect 6480 7412 6485 7428
rect 6523 7412 6548 7428
rect 6548 7412 6557 7428
rect 6595 7412 6616 7428
rect 6616 7412 6629 7428
rect 6667 7412 6684 7428
rect 6684 7412 6701 7428
rect 6739 7412 6752 7428
rect 6752 7412 6773 7428
rect 6811 7412 6820 7428
rect 6820 7412 6845 7428
rect 6883 7412 6888 7428
rect 6888 7412 6917 7428
rect 6955 7412 6956 7428
rect 6956 7412 6989 7428
rect 7027 7412 7058 7428
rect 7058 7412 7061 7428
rect 7099 7412 7126 7428
rect 7126 7412 7133 7428
rect 7171 7412 7194 7428
rect 7194 7412 7205 7428
rect 7243 7412 7262 7428
rect 7262 7412 7277 7428
rect 7315 7412 7330 7428
rect 7330 7412 7349 7428
rect 7387 7412 7398 7428
rect 7398 7412 7421 7428
rect 7459 7412 7466 7428
rect 7466 7412 7493 7428
rect 7531 7412 7534 7428
rect 7534 7412 7565 7428
rect 7603 7412 7636 7428
rect 7636 7412 7637 7428
rect 7675 7412 7704 7428
rect 7704 7412 7709 7428
rect 7747 7412 7772 7428
rect 7772 7412 7781 7428
rect 7819 7412 7840 7428
rect 7840 7412 7853 7428
rect 7891 7412 7908 7428
rect 7908 7412 7925 7428
rect 7963 7412 7976 7428
rect 7976 7412 7997 7428
rect 8035 7412 8044 7428
rect 8044 7412 8069 7428
rect 8107 7412 8112 7428
rect 8112 7412 8141 7428
rect 8179 7412 8180 7428
rect 8180 7412 8213 7428
rect 8251 7412 8282 7428
rect 8282 7412 8285 7428
rect 8323 7412 8350 7428
rect 8350 7412 8357 7428
rect 8395 7412 8418 7428
rect 8418 7412 8429 7428
rect 8467 7412 8486 7428
rect 8486 7412 8501 7428
rect 8539 7412 8554 7428
rect 8554 7412 8573 7428
rect 8611 7412 8622 7428
rect 8622 7412 8645 7428
rect 8683 7412 8690 7428
rect 8690 7412 8717 7428
rect 8755 7412 8758 7428
rect 8758 7412 8789 7428
rect 8827 7412 8860 7428
rect 8860 7412 8861 7428
rect 8899 7412 8928 7428
rect 8928 7412 8933 7428
rect 8971 7412 8996 7428
rect 8996 7412 9005 7428
rect 5941 7394 5975 7412
rect 6014 7394 6048 7412
rect 6087 7394 6121 7412
rect 6160 7394 6194 7412
rect 6233 7394 6267 7412
rect 6306 7394 6340 7412
rect 6379 7394 6413 7412
rect 6451 7394 6485 7412
rect 6523 7394 6557 7412
rect 6595 7394 6629 7412
rect 6667 7394 6701 7412
rect 6739 7394 6773 7412
rect 6811 7394 6845 7412
rect 6883 7394 6917 7412
rect 6955 7394 6989 7412
rect 7027 7394 7061 7412
rect 7099 7394 7133 7412
rect 7171 7394 7205 7412
rect 7243 7394 7277 7412
rect 7315 7394 7349 7412
rect 7387 7394 7421 7412
rect 7459 7394 7493 7412
rect 7531 7394 7565 7412
rect 7603 7394 7637 7412
rect 7675 7394 7709 7412
rect 7747 7394 7781 7412
rect 7819 7394 7853 7412
rect 7891 7394 7925 7412
rect 7963 7394 7997 7412
rect 8035 7394 8069 7412
rect 8107 7394 8141 7412
rect 8179 7394 8213 7412
rect 8251 7394 8285 7412
rect 8323 7394 8357 7412
rect 8395 7394 8429 7412
rect 8467 7394 8501 7412
rect 8539 7394 8573 7412
rect 8611 7394 8645 7412
rect 8683 7394 8717 7412
rect 8755 7394 8789 7412
rect 8827 7394 8861 7412
rect 8899 7394 8933 7412
rect 8971 7394 9005 7412
rect 9157 7416 9185 7445
rect 9185 7416 9191 7445
rect 9157 7411 9191 7416
rect 947 7349 981 7372
rect 947 7338 981 7349
rect 9157 7348 9185 7371
rect 9185 7348 9191 7371
rect 9157 7337 9191 7348
rect 947 7281 981 7297
rect 947 7263 981 7281
rect 947 7213 981 7222
rect 947 7188 981 7213
rect 947 7145 981 7147
rect 947 7113 981 7145
rect 947 7043 981 7072
rect 947 7038 981 7043
rect 947 6975 981 6997
rect 947 6963 981 6975
rect 947 6907 981 6922
rect 947 6888 981 6907
rect 947 6839 981 6847
rect 947 6813 981 6839
rect 947 6771 981 6772
rect 947 6738 981 6771
rect 947 6669 981 6697
rect 947 6663 981 6669
rect 1223 7264 1257 7298
rect 1223 7190 1257 7224
rect 1223 7116 1257 7150
rect 1223 7042 1257 7076
rect 1223 6968 1257 7002
rect 1223 6893 1257 6927
rect 1223 6818 1257 6852
rect 1223 6743 1257 6777
rect 1223 6668 1257 6702
rect 1535 7264 1569 7298
rect 1535 7190 1569 7224
rect 1535 7116 1569 7150
rect 1535 7042 1569 7076
rect 1535 6967 1569 7001
rect 1535 6892 1569 6926
rect 1535 6817 1569 6851
rect 1535 6742 1569 6776
rect 1535 6667 1569 6701
rect 1847 7264 1881 7298
rect 1847 7190 1881 7224
rect 1847 7116 1881 7150
rect 1847 7042 1881 7076
rect 1847 6968 1881 7002
rect 1847 6893 1881 6927
rect 1847 6818 1881 6852
rect 1847 6743 1881 6777
rect 1847 6668 1881 6702
rect 2159 7264 2193 7298
rect 2159 7190 2193 7224
rect 2159 7116 2193 7150
rect 2159 7042 2193 7076
rect 2159 6967 2193 7001
rect 2159 6892 2193 6926
rect 2159 6817 2193 6851
rect 2159 6742 2193 6776
rect 2159 6667 2193 6701
rect 2471 7264 2505 7298
rect 2471 7190 2505 7224
rect 2471 7116 2505 7150
rect 2471 7042 2505 7076
rect 2471 6968 2505 7002
rect 2471 6893 2505 6927
rect 2471 6818 2505 6852
rect 2471 6743 2505 6777
rect 2471 6668 2505 6702
rect 2783 7264 2817 7298
rect 2783 7190 2817 7224
rect 2783 7116 2817 7150
rect 2783 7042 2817 7076
rect 2783 6967 2817 7001
rect 2783 6892 2817 6926
rect 2783 6817 2817 6851
rect 2783 6742 2817 6776
rect 2783 6667 2817 6701
rect 3095 7264 3129 7298
rect 3095 7190 3129 7224
rect 3095 7116 3129 7150
rect 3095 7042 3129 7076
rect 3095 6968 3129 7002
rect 3095 6893 3129 6927
rect 3095 6818 3129 6852
rect 3095 6743 3129 6777
rect 3095 6668 3129 6702
rect 3407 7264 3441 7298
rect 3407 7190 3441 7224
rect 3407 7116 3441 7150
rect 3407 7042 3441 7076
rect 3407 6967 3441 7001
rect 3407 6892 3441 6926
rect 3407 6817 3441 6851
rect 3407 6742 3441 6776
rect 3407 6667 3441 6701
rect 3719 7264 3753 7298
rect 3719 7190 3753 7224
rect 3719 7116 3753 7150
rect 3719 7042 3753 7076
rect 3719 6968 3753 7002
rect 3719 6893 3753 6927
rect 3719 6818 3753 6852
rect 3719 6743 3753 6777
rect 3719 6668 3753 6702
rect 4031 7264 4065 7298
rect 4031 7190 4065 7224
rect 4031 7116 4065 7150
rect 4031 7042 4065 7076
rect 4031 6967 4065 7001
rect 4031 6892 4065 6926
rect 4031 6817 4065 6851
rect 4031 6742 4065 6776
rect 4031 6667 4065 6701
rect 4343 7264 4377 7298
rect 4343 7190 4377 7224
rect 4343 7116 4377 7150
rect 4343 7042 4377 7076
rect 4343 6968 4377 7002
rect 4343 6893 4377 6927
rect 4343 6818 4377 6852
rect 4343 6743 4377 6777
rect 4343 6668 4377 6702
rect 4655 7264 4689 7298
rect 4655 7190 4689 7224
rect 4655 7116 4689 7150
rect 4655 7042 4689 7076
rect 4655 6967 4689 7001
rect 4655 6892 4689 6926
rect 4655 6817 4689 6851
rect 4655 6742 4689 6776
rect 4655 6667 4689 6701
rect 4967 7264 5001 7298
rect 4967 7190 5001 7224
rect 4967 7116 5001 7150
rect 4967 7042 5001 7076
rect 4967 6968 5001 7002
rect 4967 6893 5001 6927
rect 4967 6818 5001 6852
rect 4967 6743 5001 6777
rect 4967 6668 5001 6702
rect 5279 7264 5313 7298
rect 5279 7190 5313 7224
rect 5279 7116 5313 7150
rect 5279 7042 5313 7076
rect 5279 6967 5313 7001
rect 5279 6892 5313 6926
rect 5279 6817 5313 6851
rect 5279 6742 5313 6776
rect 5279 6667 5313 6701
rect 5591 7264 5625 7298
rect 5591 7190 5625 7224
rect 5591 7116 5625 7150
rect 5591 7042 5625 7076
rect 5591 6968 5625 7002
rect 5591 6893 5625 6927
rect 5591 6818 5625 6852
rect 5591 6743 5625 6777
rect 5591 6668 5625 6702
rect 5903 7264 5937 7298
rect 5903 7190 5937 7224
rect 5903 7116 5937 7150
rect 5903 7042 5937 7076
rect 5903 6967 5937 7001
rect 5903 6892 5937 6926
rect 5903 6817 5937 6851
rect 5903 6742 5937 6776
rect 5903 6667 5937 6701
rect 6215 7264 6249 7298
rect 6215 7190 6249 7224
rect 6215 7116 6249 7150
rect 6215 7042 6249 7076
rect 6215 6968 6249 7002
rect 6215 6893 6249 6927
rect 6215 6818 6249 6852
rect 6215 6743 6249 6777
rect 6215 6668 6249 6702
rect 6527 7264 6561 7298
rect 6527 7190 6561 7224
rect 6527 7116 6561 7150
rect 6527 7042 6561 7076
rect 6527 6967 6561 7001
rect 6527 6892 6561 6926
rect 6527 6817 6561 6851
rect 6527 6742 6561 6776
rect 6527 6667 6561 6701
rect 6839 7264 6873 7298
rect 6839 7190 6873 7224
rect 6839 7116 6873 7150
rect 6839 7042 6873 7076
rect 6839 6968 6873 7002
rect 6839 6893 6873 6927
rect 6839 6818 6873 6852
rect 6839 6743 6873 6777
rect 6839 6668 6873 6702
rect 7151 7264 7185 7298
rect 7151 7190 7185 7224
rect 7151 7116 7185 7150
rect 7151 7042 7185 7076
rect 7151 6967 7185 7001
rect 7151 6892 7185 6926
rect 7151 6817 7185 6851
rect 7151 6742 7185 6776
rect 7151 6667 7185 6701
rect 7463 7264 7497 7298
rect 7463 7190 7497 7224
rect 7463 7116 7497 7150
rect 7463 7042 7497 7076
rect 7463 6968 7497 7002
rect 7463 6893 7497 6927
rect 7463 6818 7497 6852
rect 7463 6743 7497 6777
rect 7463 6668 7497 6702
rect 7775 7264 7809 7298
rect 7775 7190 7809 7224
rect 7775 7116 7809 7150
rect 7775 7042 7809 7076
rect 7775 6967 7809 7001
rect 7775 6892 7809 6926
rect 7775 6817 7809 6851
rect 7775 6742 7809 6776
rect 7775 6667 7809 6701
rect 8087 7264 8121 7298
rect 8087 7190 8121 7224
rect 8087 7116 8121 7150
rect 8087 7042 8121 7076
rect 8087 6967 8121 7001
rect 8087 6892 8121 6926
rect 8087 6817 8121 6851
rect 8087 6742 8121 6776
rect 8087 6667 8121 6701
rect 8399 7264 8433 7298
rect 8399 7190 8433 7224
rect 8399 7116 8433 7150
rect 8399 7042 8433 7076
rect 8399 6968 8433 7002
rect 8399 6893 8433 6927
rect 8399 6818 8433 6852
rect 8399 6743 8433 6777
rect 8399 6668 8433 6702
rect 8711 7264 8745 7298
rect 8711 7190 8745 7224
rect 8711 7116 8745 7150
rect 8711 7042 8745 7076
rect 8711 6967 8745 7001
rect 8711 6892 8745 6926
rect 8711 6817 8745 6851
rect 8711 6742 8745 6776
rect 8711 6667 8745 6701
rect 9023 7264 9057 7298
rect 9023 7190 9057 7224
rect 9023 7116 9057 7150
rect 9023 7042 9057 7076
rect 9023 6968 9057 7002
rect 9023 6893 9057 6927
rect 9023 6818 9057 6852
rect 9023 6743 9057 6777
rect 9023 6668 9057 6702
rect 9157 7280 9185 7297
rect 9185 7280 9191 7297
rect 9157 7263 9191 7280
rect 9157 7212 9185 7223
rect 9185 7212 9191 7223
rect 9157 7189 9191 7212
rect 9157 7144 9185 7149
rect 9185 7144 9191 7149
rect 9157 7115 9191 7144
rect 9157 7042 9191 7075
rect 9157 7041 9185 7042
rect 9185 7041 9191 7042
rect 9157 6974 9191 7001
rect 9157 6967 9185 6974
rect 9185 6967 9191 6974
rect 9157 6906 9191 6926
rect 9157 6892 9185 6906
rect 9185 6892 9191 6906
rect 9157 6838 9191 6851
rect 9157 6817 9185 6838
rect 9185 6817 9191 6838
rect 9157 6770 9191 6776
rect 9157 6742 9185 6770
rect 9185 6742 9191 6770
rect 9157 6668 9185 6701
rect 9185 6668 9191 6701
rect 9157 6667 9191 6668
rect 947 6601 981 6622
rect 947 6588 981 6601
rect 9157 6600 9185 6626
rect 9185 6600 9191 6626
rect 9157 6592 9191 6600
rect 947 6533 981 6547
rect 947 6513 981 6533
rect 947 6465 981 6472
rect 947 6438 981 6465
rect 947 6397 981 6398
rect 947 6364 981 6397
rect 947 6295 981 6324
rect 947 6290 981 6295
rect 947 6227 981 6250
rect 947 6216 981 6227
rect 947 6159 981 6176
rect 947 6142 981 6159
rect 947 6091 981 6102
rect 947 6068 981 6091
rect 947 6023 981 6028
rect 947 5994 981 6023
rect 1379 6538 1413 6572
rect 1379 6466 1413 6500
rect 1379 6393 1413 6427
rect 1379 6320 1413 6354
rect 1379 6247 1413 6281
rect 1379 6174 1413 6208
rect 1379 6101 1413 6135
rect 1379 6028 1413 6062
rect 1379 5955 1413 5989
rect 1691 6538 1725 6572
rect 1691 6465 1725 6499
rect 1691 6392 1725 6426
rect 1691 6319 1725 6353
rect 1691 6246 1725 6280
rect 1691 6173 1725 6207
rect 1691 6100 1725 6134
rect 1691 6027 1725 6061
rect 1691 5954 1725 5988
rect 2003 6538 2037 6572
rect 2003 6466 2037 6500
rect 2003 6393 2037 6427
rect 2003 6320 2037 6354
rect 2003 6247 2037 6281
rect 2003 6174 2037 6208
rect 2003 6101 2037 6135
rect 2003 6028 2037 6062
rect 2003 5955 2037 5989
rect 2315 6538 2349 6572
rect 2315 6465 2349 6499
rect 2315 6392 2349 6426
rect 2315 6319 2349 6353
rect 2315 6246 2349 6280
rect 2315 6173 2349 6207
rect 2315 6100 2349 6134
rect 2315 6027 2349 6061
rect 2315 5954 2349 5988
rect 2627 6538 2661 6572
rect 2627 6466 2661 6500
rect 2627 6393 2661 6427
rect 2627 6320 2661 6354
rect 2627 6247 2661 6281
rect 2627 6174 2661 6208
rect 2627 6101 2661 6135
rect 2627 6028 2661 6062
rect 2627 5955 2661 5989
rect 2939 6538 2973 6572
rect 2939 6465 2973 6499
rect 2939 6392 2973 6426
rect 2939 6319 2973 6353
rect 2939 6246 2973 6280
rect 2939 6173 2973 6207
rect 2939 6100 2973 6134
rect 2939 6027 2973 6061
rect 2939 5954 2973 5988
rect 3251 6538 3285 6572
rect 3251 6465 3285 6499
rect 3251 6392 3285 6426
rect 3251 6319 3285 6353
rect 3251 6246 3285 6280
rect 3251 6173 3285 6207
rect 3251 6100 3285 6134
rect 3251 6027 3285 6061
rect 3251 5954 3285 5988
rect 3563 6538 3597 6572
rect 3563 6465 3597 6499
rect 3563 6392 3597 6426
rect 3563 6319 3597 6353
rect 3563 6246 3597 6280
rect 3563 6173 3597 6207
rect 3563 6100 3597 6134
rect 3563 6027 3597 6061
rect 3563 5954 3597 5988
rect 3875 6538 3909 6572
rect 3875 6466 3909 6500
rect 3875 6393 3909 6427
rect 3875 6320 3909 6354
rect 3875 6247 3909 6281
rect 3875 6174 3909 6208
rect 3875 6101 3909 6135
rect 3875 6028 3909 6062
rect 3875 5955 3909 5989
rect 4187 6538 4221 6572
rect 4187 6465 4221 6499
rect 4187 6392 4221 6426
rect 4187 6319 4221 6353
rect 4187 6246 4221 6280
rect 4187 6173 4221 6207
rect 4187 6100 4221 6134
rect 4187 6027 4221 6061
rect 4187 5954 4221 5988
rect 4499 6538 4533 6572
rect 4499 6466 4533 6500
rect 4499 6393 4533 6427
rect 4499 6320 4533 6354
rect 4499 6247 4533 6281
rect 4499 6174 4533 6208
rect 4499 6101 4533 6135
rect 4499 6028 4533 6062
rect 4499 5955 4533 5989
rect 4811 6538 4845 6572
rect 4811 6465 4845 6499
rect 4811 6392 4845 6426
rect 4811 6319 4845 6353
rect 4811 6246 4845 6280
rect 4811 6173 4845 6207
rect 4811 6100 4845 6134
rect 4811 6027 4845 6061
rect 4811 5954 4845 5988
rect 5123 6538 5157 6572
rect 5123 6466 5157 6500
rect 5123 6393 5157 6427
rect 5123 6320 5157 6354
rect 5123 6247 5157 6281
rect 5123 6174 5157 6208
rect 5123 6101 5157 6135
rect 5123 6028 5157 6062
rect 5123 5955 5157 5989
rect 5435 6538 5469 6572
rect 5435 6465 5469 6499
rect 5435 6392 5469 6426
rect 5435 6319 5469 6353
rect 5435 6246 5469 6280
rect 5435 6173 5469 6207
rect 5435 6100 5469 6134
rect 5435 6027 5469 6061
rect 5435 5954 5469 5988
rect 5747 6538 5781 6572
rect 5747 6466 5781 6500
rect 5747 6393 5781 6427
rect 5747 6320 5781 6354
rect 5747 6247 5781 6281
rect 5747 6174 5781 6208
rect 5747 6101 5781 6135
rect 5747 6028 5781 6062
rect 5747 5955 5781 5989
rect 6059 6538 6093 6572
rect 6059 6465 6093 6499
rect 6059 6392 6093 6426
rect 6059 6319 6093 6353
rect 6059 6246 6093 6280
rect 6059 6173 6093 6207
rect 6059 6100 6093 6134
rect 6059 6027 6093 6061
rect 6059 5954 6093 5988
rect 6371 6538 6405 6572
rect 6371 6466 6405 6500
rect 6371 6393 6405 6427
rect 6371 6320 6405 6354
rect 6371 6247 6405 6281
rect 6371 6174 6405 6208
rect 6371 6101 6405 6135
rect 6371 6028 6405 6062
rect 6371 5955 6405 5989
rect 6683 6538 6717 6572
rect 6683 6465 6717 6499
rect 6683 6392 6717 6426
rect 6683 6319 6717 6353
rect 6683 6246 6717 6280
rect 6683 6173 6717 6207
rect 6683 6100 6717 6134
rect 6683 6027 6717 6061
rect 6683 5954 6717 5988
rect 6995 6538 7029 6572
rect 6995 6466 7029 6500
rect 6995 6393 7029 6427
rect 6995 6320 7029 6354
rect 6995 6247 7029 6281
rect 6995 6174 7029 6208
rect 6995 6101 7029 6135
rect 6995 6028 7029 6062
rect 6995 5955 7029 5989
rect 7307 6538 7341 6572
rect 7307 6465 7341 6499
rect 7307 6392 7341 6426
rect 7307 6319 7341 6353
rect 7307 6246 7341 6280
rect 7307 6173 7341 6207
rect 7307 6100 7341 6134
rect 7307 6027 7341 6061
rect 7307 5954 7341 5988
rect 7619 6538 7653 6572
rect 7619 6466 7653 6500
rect 7619 6393 7653 6427
rect 7619 6320 7653 6354
rect 7619 6247 7653 6281
rect 7619 6174 7653 6208
rect 7619 6101 7653 6135
rect 7619 6028 7653 6062
rect 7619 5955 7653 5989
rect 7931 6538 7965 6572
rect 7931 6465 7965 6499
rect 7931 6392 7965 6426
rect 7931 6319 7965 6353
rect 7931 6246 7965 6280
rect 7931 6173 7965 6207
rect 7931 6100 7965 6134
rect 7931 6027 7965 6061
rect 7931 5954 7965 5988
rect 8243 6538 8277 6572
rect 8243 6465 8277 6499
rect 8243 6392 8277 6426
rect 8243 6319 8277 6353
rect 8243 6246 8277 6280
rect 8243 6173 8277 6207
rect 8243 6100 8277 6134
rect 8243 6027 8277 6061
rect 8243 5954 8277 5988
rect 8555 6538 8589 6572
rect 8555 6466 8589 6500
rect 8555 6393 8589 6427
rect 8555 6320 8589 6354
rect 8555 6247 8589 6281
rect 8555 6174 8589 6208
rect 8555 6101 8589 6135
rect 8555 6028 8589 6062
rect 8555 5955 8589 5989
rect 8867 6538 8901 6572
rect 8867 6465 8901 6499
rect 8867 6392 8901 6426
rect 8867 6319 8901 6353
rect 8867 6246 8901 6280
rect 8867 6173 8901 6207
rect 8867 6100 8901 6134
rect 8867 6027 8901 6061
rect 8867 5954 8901 5988
rect 9157 6532 9185 6551
rect 9185 6532 9191 6551
rect 9157 6517 9191 6532
rect 9157 6464 9185 6476
rect 9185 6464 9191 6476
rect 9157 6442 9191 6464
rect 9157 6396 9185 6401
rect 9185 6396 9191 6401
rect 9157 6367 9191 6396
rect 9157 6294 9191 6326
rect 9157 6292 9185 6294
rect 9185 6292 9191 6294
rect 9157 6226 9191 6251
rect 9157 6217 9185 6226
rect 9185 6217 9191 6226
rect 9157 6158 9191 6176
rect 9157 6142 9185 6158
rect 9185 6142 9191 6158
rect 9157 6090 9191 6101
rect 9157 6067 9185 6090
rect 9185 6067 9191 6090
rect 9157 6022 9191 6026
rect 9157 5992 9185 6022
rect 9185 5992 9191 6022
rect 947 5920 981 5954
rect 9157 5920 9185 5951
rect 9185 5920 9191 5951
rect 9157 5917 9191 5920
rect 9462 7517 9466 7551
rect 9466 7517 9496 7551
rect 9534 7515 9568 7549
rect 9606 7515 9636 7549
rect 9636 7515 9640 7549
rect 9462 7443 9466 7477
rect 9466 7443 9496 7477
rect 9534 7441 9568 7475
rect 9606 7441 9636 7475
rect 9636 7441 9640 7475
rect 9462 7369 9466 7403
rect 9466 7369 9496 7403
rect 9534 7367 9568 7401
rect 9606 7367 9636 7401
rect 9636 7367 9640 7401
rect 9462 7295 9466 7329
rect 9466 7295 9496 7329
rect 9534 7293 9568 7327
rect 9606 7293 9636 7327
rect 9636 7293 9640 7327
rect 9462 7221 9466 7255
rect 9466 7221 9496 7255
rect 9534 7219 9568 7253
rect 9606 7219 9636 7253
rect 9636 7219 9640 7253
rect 9462 7147 9466 7181
rect 9466 7147 9496 7181
rect 9534 7146 9568 7180
rect 9606 7146 9636 7180
rect 9636 7146 9640 7180
rect 9462 7073 9466 7107
rect 9466 7073 9496 7107
rect 9534 7073 9568 7107
rect 9606 7073 9636 7107
rect 9636 7073 9640 7107
rect 9462 7000 9466 7034
rect 9466 7000 9496 7034
rect 9534 7000 9568 7034
rect 9606 7000 9636 7034
rect 9636 7000 9640 7034
rect 9462 6927 9466 6961
rect 9466 6927 9496 6961
rect 9534 6927 9568 6961
rect 9606 6927 9636 6961
rect 9636 6927 9640 6961
rect 9462 6854 9466 6888
rect 9466 6854 9496 6888
rect 9534 6854 9568 6888
rect 9606 6854 9636 6888
rect 9636 6854 9640 6888
rect 9462 6781 9466 6815
rect 9466 6781 9496 6815
rect 9534 6781 9568 6815
rect 9606 6781 9636 6815
rect 9636 6781 9640 6815
rect 9462 6708 9466 6742
rect 9466 6708 9496 6742
rect 9534 6708 9568 6742
rect 9606 6708 9636 6742
rect 9636 6708 9640 6742
rect 9462 6635 9466 6669
rect 9466 6635 9496 6669
rect 9534 6635 9568 6669
rect 9606 6635 9636 6669
rect 9636 6635 9640 6669
rect 9462 6562 9466 6596
rect 9466 6562 9496 6596
rect 9534 6562 9568 6596
rect 9606 6562 9636 6596
rect 9636 6562 9640 6596
rect 9462 6489 9466 6523
rect 9466 6489 9496 6523
rect 9534 6489 9568 6523
rect 9606 6489 9636 6523
rect 9636 6489 9640 6523
rect 9462 6416 9466 6450
rect 9466 6416 9496 6450
rect 9534 6416 9568 6450
rect 9606 6416 9636 6450
rect 9636 6416 9640 6450
rect 9462 6343 9466 6377
rect 9466 6343 9496 6377
rect 9534 6343 9568 6377
rect 9606 6343 9636 6377
rect 9636 6343 9640 6377
rect 9462 6270 9466 6304
rect 9466 6270 9496 6304
rect 9534 6270 9568 6304
rect 9606 6270 9636 6304
rect 9636 6270 9640 6304
rect 9462 6197 9466 6231
rect 9466 6197 9496 6231
rect 9534 6197 9568 6231
rect 9606 6197 9636 6231
rect 9636 6197 9640 6231
rect 9462 6124 9466 6158
rect 9466 6124 9496 6158
rect 9534 6124 9568 6158
rect 9606 6124 9636 6158
rect 9636 6124 9640 6158
rect 9462 6051 9466 6085
rect 9466 6051 9496 6085
rect 9534 6051 9568 6085
rect 9606 6051 9636 6085
rect 9636 6051 9640 6085
rect 9462 5978 9466 6012
rect 9466 5978 9496 6012
rect 9534 5978 9568 6012
rect 9606 5978 9636 6012
rect 9636 5978 9640 6012
rect 9462 5905 9466 5939
rect 9466 5905 9496 5939
rect 9534 5905 9568 5939
rect 9606 5905 9636 5939
rect 9636 5905 9640 5939
rect 10464 7913 10498 7915
rect 10464 7881 10473 7913
rect 10473 7881 10498 7913
rect 10536 7881 10570 7915
rect 10608 7883 10639 7917
rect 10639 7883 10642 7917
rect 10464 7811 10473 7842
rect 10473 7811 10498 7842
rect 10464 7808 10498 7811
rect 10536 7808 10570 7842
rect 10608 7815 10639 7844
rect 10639 7815 10642 7844
rect 10608 7810 10642 7815
rect 10464 7743 10473 7769
rect 10473 7743 10498 7769
rect 10464 7735 10498 7743
rect 10536 7735 10570 7769
rect 10608 7747 10639 7771
rect 10639 7747 10642 7771
rect 10608 7737 10642 7747
rect 10464 7675 10473 7696
rect 10473 7675 10498 7696
rect 10464 7662 10498 7675
rect 10536 7662 10570 7696
rect 10608 7679 10639 7698
rect 10639 7679 10642 7698
rect 10608 7664 10642 7679
rect 10464 7607 10473 7623
rect 10473 7607 10498 7623
rect 10464 7589 10498 7607
rect 10536 7589 10570 7623
rect 10608 7611 10639 7625
rect 10639 7611 10642 7625
rect 10608 7591 10642 7611
rect 10464 7539 10473 7550
rect 10473 7539 10498 7550
rect 10464 7516 10498 7539
rect 10536 7516 10570 7550
rect 10608 7543 10639 7552
rect 10639 7543 10642 7552
rect 10608 7518 10642 7543
rect 10464 7471 10473 7477
rect 10473 7471 10498 7477
rect 10464 7443 10498 7471
rect 10536 7443 10570 7477
rect 10608 7475 10639 7479
rect 10639 7475 10642 7479
rect 10608 7445 10642 7475
rect 10464 7403 10473 7404
rect 10473 7403 10498 7404
rect 10464 7370 10498 7403
rect 10536 7370 10570 7404
rect 10608 7373 10642 7406
rect 10608 7372 10639 7373
rect 10639 7372 10642 7373
rect 10464 7301 10498 7331
rect 10464 7297 10473 7301
rect 10473 7297 10498 7301
rect 10536 7297 10570 7331
rect 10608 7305 10642 7333
rect 10608 7299 10639 7305
rect 10639 7299 10642 7305
rect 10464 7233 10498 7258
rect 10464 7224 10473 7233
rect 10473 7224 10498 7233
rect 10536 7224 10570 7258
rect 10608 7237 10642 7260
rect 10608 7226 10639 7237
rect 10639 7226 10642 7237
rect 10464 7165 10498 7185
rect 10464 7151 10473 7165
rect 10473 7151 10498 7165
rect 10536 7151 10570 7185
rect 10608 7169 10642 7187
rect 10608 7153 10639 7169
rect 10639 7153 10642 7169
rect 10464 7097 10498 7112
rect 10464 7078 10473 7097
rect 10473 7078 10498 7097
rect 10536 7078 10570 7112
rect 10608 7101 10642 7113
rect 10608 7079 10639 7101
rect 10639 7079 10642 7101
rect 10464 7029 10498 7039
rect 10464 7005 10473 7029
rect 10473 7005 10498 7029
rect 10536 7005 10570 7039
rect 10608 7033 10642 7039
rect 10608 7005 10639 7033
rect 10639 7005 10642 7033
rect 10464 6961 10498 6965
rect 10464 6931 10473 6961
rect 10473 6931 10498 6961
rect 10536 6931 10570 6965
rect 10608 6931 10639 6965
rect 10639 6931 10642 6965
rect 10464 6859 10473 6891
rect 10473 6859 10498 6891
rect 10464 6857 10498 6859
rect 10536 6857 10570 6891
rect 10608 6863 10639 6891
rect 10639 6863 10642 6891
rect 10608 6857 10642 6863
rect 10464 6791 10473 6817
rect 10473 6791 10498 6817
rect 10464 6783 10498 6791
rect 10536 6783 10570 6817
rect 10608 6795 10639 6817
rect 10639 6795 10642 6817
rect 10608 6783 10642 6795
rect 10464 6723 10473 6743
rect 10473 6723 10498 6743
rect 10464 6709 10498 6723
rect 10536 6709 10570 6743
rect 10608 6727 10639 6743
rect 10639 6727 10642 6743
rect 10608 6709 10642 6727
rect 10464 6655 10473 6669
rect 10473 6655 10498 6669
rect 10464 6635 10498 6655
rect 10536 6635 10570 6669
rect 10608 6659 10639 6669
rect 10639 6659 10642 6669
rect 10608 6635 10642 6659
rect 10464 6587 10473 6595
rect 10473 6587 10498 6595
rect 10464 6561 10498 6587
rect 10536 6561 10570 6595
rect 10608 6591 10639 6595
rect 10639 6591 10642 6595
rect 10608 6561 10642 6591
rect 10464 6519 10473 6521
rect 10473 6519 10498 6521
rect 10464 6487 10498 6519
rect 10536 6487 10570 6521
rect 10608 6489 10642 6521
rect 10608 6487 10639 6489
rect 10639 6487 10642 6489
rect 10464 6394 10498 6428
rect 10536 6394 10570 6428
rect 10608 6394 10642 6428
rect 10864 8082 10878 8116
rect 10878 8082 10898 8116
rect 10936 8082 10946 8116
rect 10946 8082 10970 8116
rect 11008 8082 11014 8116
rect 11014 8082 11042 8116
rect 11080 8082 11082 8116
rect 11082 8082 11114 8116
rect 11152 8082 11184 8116
rect 11184 8082 11186 8116
rect 11224 8082 11252 8116
rect 11252 8082 11258 8116
rect 11296 8082 11320 8116
rect 11320 8082 11330 8116
rect 11368 8082 11388 8116
rect 11388 8082 11402 8116
rect 11440 8082 11456 8116
rect 11456 8082 11474 8116
rect 11512 8082 11524 8116
rect 11524 8082 11546 8116
rect 11584 8082 11592 8116
rect 11592 8082 11618 8116
rect 11656 8082 11660 8116
rect 11660 8082 11690 8116
rect 11728 8082 11762 8116
rect 11800 8082 11830 8116
rect 11830 8082 11834 8116
rect 11872 8082 11898 8116
rect 11898 8082 11906 8116
rect 11944 8082 11966 8116
rect 11966 8082 11978 8116
rect 12016 8082 12034 8116
rect 12034 8082 12050 8116
rect 12088 8082 12102 8116
rect 12102 8082 12122 8116
rect 12160 8082 12170 8116
rect 12170 8082 12194 8116
rect 12232 8082 12238 8116
rect 12238 8082 12266 8116
rect 12304 8082 12306 8116
rect 12306 8082 12338 8116
rect 12376 8082 12408 8116
rect 12408 8082 12410 8116
rect 12448 8082 12476 8116
rect 12476 8082 12482 8116
rect 12520 8082 12544 8116
rect 12544 8082 12554 8116
rect 12592 8082 12612 8116
rect 12612 8082 12626 8116
rect 12664 8082 12680 8116
rect 12680 8082 12698 8116
rect 12736 8082 12748 8116
rect 12748 8082 12770 8116
rect 12808 8082 12816 8116
rect 12816 8082 12842 8116
rect 12880 8082 12884 8116
rect 12884 8082 12914 8116
rect 12952 8082 12986 8116
rect 13024 8082 13054 8116
rect 13054 8082 13058 8116
rect 13096 8082 13122 8116
rect 13122 8082 13130 8116
rect 13169 8082 13190 8116
rect 13190 8082 13203 8116
rect 13242 8082 13258 8116
rect 13258 8082 13276 8116
rect 13315 8082 13326 8116
rect 13326 8082 13349 8116
rect 13387 8033 13421 8041
rect 13387 8007 13394 8033
rect 13394 8007 13421 8033
rect 10995 7954 11004 7988
rect 11004 7954 11029 7988
rect 11070 7954 11074 7988
rect 11074 7954 11104 7988
rect 11145 7954 11178 7988
rect 11178 7954 11179 7988
rect 11220 7954 11248 7988
rect 11248 7954 11254 7988
rect 11295 7954 11318 7988
rect 11318 7954 11329 7988
rect 11370 7954 11388 7988
rect 11388 7954 11404 7988
rect 11445 7954 11457 7988
rect 11457 7954 11479 7988
rect 11519 7954 11526 7988
rect 11526 7954 11553 7988
rect 11593 7954 11595 7988
rect 11595 7954 11627 7988
rect 11667 7954 11699 7988
rect 11699 7954 11701 7988
rect 11741 7954 11768 7988
rect 11768 7954 11775 7988
rect 11815 7954 11837 7988
rect 11837 7954 11849 7988
rect 11889 7954 11906 7988
rect 11906 7954 11923 7988
rect 11963 7954 11975 7988
rect 11975 7954 11997 7988
rect 12037 7954 12044 7988
rect 12044 7954 12071 7988
rect 12111 7954 12113 7988
rect 12113 7954 12145 7988
rect 12185 7954 12216 7988
rect 12216 7954 12219 7988
rect 12259 7954 12285 7988
rect 12285 7954 12293 7988
rect 12333 7954 12354 7988
rect 12354 7954 12367 7988
rect 12407 7954 12423 7988
rect 12423 7954 12441 7988
rect 12481 7954 12492 7988
rect 12492 7954 12515 7988
rect 12555 7954 12561 7988
rect 12561 7954 12589 7988
rect 12629 7954 12630 7988
rect 12630 7954 12663 7988
rect 12703 7954 12734 7988
rect 12734 7954 12737 7988
rect 12777 7954 12803 7988
rect 12803 7954 12811 7988
rect 12851 7954 12872 7988
rect 12872 7954 12885 7988
rect 12925 7954 12941 7988
rect 12941 7954 12959 7988
rect 12999 7954 13010 7988
rect 13010 7954 13033 7988
rect 13073 7954 13079 7988
rect 13079 7954 13107 7988
rect 13147 7954 13148 7988
rect 13148 7954 13181 7988
rect 13221 7954 13251 7988
rect 13251 7954 13255 7988
rect 13387 7965 13421 7966
rect 13387 7932 13394 7965
rect 13394 7932 13421 7965
rect 13387 7863 13394 7891
rect 13394 7863 13421 7891
rect 10792 7844 10826 7858
rect 10792 7824 10826 7844
rect 10792 7776 10826 7784
rect 10792 7750 10826 7776
rect 10792 7708 10826 7710
rect 10792 7676 10826 7708
rect 10792 7606 10826 7636
rect 10792 7602 10826 7606
rect 10792 7538 10826 7563
rect 10792 7529 10826 7538
rect 10792 7470 10826 7490
rect 10792 7456 10826 7470
rect 10792 7402 10826 7417
rect 10792 7383 10826 7402
rect 10792 7334 10826 7344
rect 10792 7310 10826 7334
rect 10792 7266 10826 7271
rect 10792 7237 10826 7266
rect 10939 7824 10973 7858
rect 10939 7751 10973 7785
rect 10939 7678 10973 7712
rect 10939 7605 10973 7639
rect 10939 7532 10973 7566
rect 10939 7459 10973 7493
rect 10939 7386 10973 7420
rect 10939 7312 10973 7346
rect 10939 7238 10973 7272
rect 11251 7824 11285 7858
rect 11251 7751 11285 7785
rect 11251 7678 11285 7712
rect 11251 7605 11285 7639
rect 11251 7532 11285 7566
rect 11251 7459 11285 7493
rect 11251 7386 11285 7420
rect 11251 7312 11285 7346
rect 11251 7238 11285 7272
rect 11563 7824 11597 7858
rect 11563 7751 11597 7785
rect 11563 7678 11597 7712
rect 11563 7605 11597 7639
rect 11563 7532 11597 7566
rect 11563 7459 11597 7493
rect 11563 7386 11597 7420
rect 11563 7312 11597 7346
rect 11563 7238 11597 7272
rect 11875 7824 11909 7858
rect 11875 7751 11909 7785
rect 11875 7678 11909 7712
rect 11875 7605 11909 7639
rect 11875 7532 11909 7566
rect 11875 7459 11909 7493
rect 11875 7386 11909 7420
rect 11875 7312 11909 7346
rect 11875 7238 11909 7272
rect 12187 7824 12221 7858
rect 12187 7751 12221 7785
rect 12187 7678 12221 7712
rect 12187 7605 12221 7639
rect 12187 7532 12221 7566
rect 12187 7459 12221 7493
rect 12187 7386 12221 7420
rect 12187 7312 12221 7346
rect 12187 7238 12221 7272
rect 12499 7824 12533 7858
rect 12499 7751 12533 7785
rect 12499 7678 12533 7712
rect 12499 7605 12533 7639
rect 12499 7532 12533 7566
rect 12499 7459 12533 7493
rect 12499 7386 12533 7420
rect 12499 7312 12533 7346
rect 12499 7238 12533 7272
rect 12811 7824 12845 7858
rect 12811 7751 12845 7785
rect 12811 7678 12845 7712
rect 12811 7605 12845 7639
rect 12811 7532 12845 7566
rect 12811 7459 12845 7493
rect 12811 7386 12845 7420
rect 12811 7312 12845 7346
rect 12811 7238 12845 7272
rect 13123 7824 13157 7858
rect 13123 7751 13157 7785
rect 13123 7678 13157 7712
rect 13123 7605 13157 7639
rect 13123 7532 13157 7566
rect 13123 7459 13157 7493
rect 13123 7386 13157 7420
rect 13123 7312 13157 7346
rect 13123 7238 13157 7272
rect 13387 7857 13421 7863
rect 13387 7795 13394 7816
rect 13394 7795 13421 7816
rect 13387 7782 13421 7795
rect 13387 7727 13394 7741
rect 13394 7727 13421 7741
rect 13387 7707 13421 7727
rect 13387 7659 13394 7666
rect 13394 7659 13421 7666
rect 13387 7632 13421 7659
rect 13387 7557 13421 7591
rect 13387 7489 13421 7516
rect 13387 7482 13394 7489
rect 13394 7482 13421 7489
rect 13387 7421 13421 7441
rect 13387 7407 13394 7421
rect 13394 7407 13421 7421
rect 13387 7353 13421 7365
rect 13387 7331 13394 7353
rect 13394 7331 13421 7353
rect 13387 7285 13421 7289
rect 13387 7255 13394 7285
rect 13394 7255 13421 7285
rect 13387 7183 13394 7213
rect 13394 7183 13421 7213
rect 13387 7179 13421 7183
rect 11093 7120 11127 7154
rect 11093 7046 11127 7080
rect 11093 6972 11127 7006
rect 11093 6898 11127 6932
rect 11093 6824 11127 6858
rect 11093 6749 11127 6783
rect 11093 6674 11127 6708
rect 11093 6599 11127 6633
rect 11093 6524 11127 6558
rect 11405 7120 11439 7154
rect 11405 7046 11439 7080
rect 11405 6972 11439 7006
rect 11405 6898 11439 6932
rect 11405 6824 11439 6858
rect 11405 6749 11439 6783
rect 11405 6674 11439 6708
rect 11405 6599 11439 6633
rect 11405 6524 11439 6558
rect 11717 7120 11751 7154
rect 11717 7046 11751 7080
rect 11717 6972 11751 7006
rect 11717 6898 11751 6932
rect 11717 6824 11751 6858
rect 11717 6749 11751 6783
rect 11717 6674 11751 6708
rect 11717 6599 11751 6633
rect 11717 6524 11751 6558
rect 12029 7120 12063 7154
rect 12029 7046 12063 7080
rect 12029 6972 12063 7006
rect 12029 6898 12063 6932
rect 12029 6824 12063 6858
rect 12029 6749 12063 6783
rect 12029 6674 12063 6708
rect 12029 6599 12063 6633
rect 12029 6524 12063 6558
rect 12341 7120 12375 7154
rect 12341 7046 12375 7080
rect 12341 6972 12375 7006
rect 12341 6898 12375 6932
rect 12341 6824 12375 6858
rect 12341 6749 12375 6783
rect 12341 6674 12375 6708
rect 12341 6599 12375 6633
rect 12341 6524 12375 6558
rect 12653 7120 12687 7154
rect 12653 7046 12687 7080
rect 12653 6972 12687 7006
rect 12653 6898 12687 6932
rect 12653 6824 12687 6858
rect 12653 6749 12687 6783
rect 12653 6674 12687 6708
rect 12653 6599 12687 6633
rect 12653 6524 12687 6558
rect 12965 7120 12999 7154
rect 12965 7046 12999 7080
rect 12965 6972 12999 7006
rect 12965 6898 12999 6932
rect 12965 6824 12999 6858
rect 12965 6749 12999 6783
rect 12965 6674 12999 6708
rect 12965 6599 12999 6633
rect 12965 6524 12999 6558
rect 13277 7120 13311 7154
rect 13277 7046 13311 7080
rect 13277 6972 13311 7006
rect 13277 6898 13311 6932
rect 13277 6824 13311 6858
rect 13277 6749 13311 6783
rect 13277 6674 13311 6708
rect 13277 6599 13311 6633
rect 13277 6524 13311 6558
rect 13387 7115 13394 7139
rect 13394 7115 13421 7139
rect 13387 7105 13421 7115
rect 13387 7047 13394 7065
rect 13394 7047 13421 7065
rect 13387 7031 13421 7047
rect 13387 6979 13394 6991
rect 13394 6979 13421 6991
rect 13387 6957 13421 6979
rect 13387 6911 13394 6917
rect 13394 6911 13421 6917
rect 13387 6883 13421 6911
rect 13387 6809 13421 6843
rect 13387 6741 13421 6769
rect 13387 6735 13394 6741
rect 13394 6735 13421 6741
rect 13387 6673 13421 6695
rect 13387 6661 13394 6673
rect 13394 6661 13421 6673
rect 13387 6605 13421 6621
rect 13387 6587 13394 6605
rect 13394 6587 13421 6605
rect 13387 6537 13421 6547
rect 13387 6513 13394 6537
rect 13394 6513 13421 6537
rect 13387 6469 13421 6473
rect 13387 6439 13394 6469
rect 13394 6439 13421 6469
rect 10864 6367 10894 6401
rect 10894 6367 10898 6401
rect 10937 6367 10962 6401
rect 10962 6367 10971 6401
rect 11010 6367 11030 6401
rect 11030 6367 11044 6401
rect 11083 6367 11098 6401
rect 11098 6367 11117 6401
rect 11155 6367 11166 6401
rect 11166 6367 11189 6401
rect 11227 6367 11234 6401
rect 11234 6367 11261 6401
rect 11299 6367 11302 6401
rect 11302 6367 11333 6401
rect 11371 6367 11404 6401
rect 11404 6367 11405 6401
rect 11443 6367 11472 6401
rect 11472 6367 11477 6401
rect 11515 6367 11540 6401
rect 11540 6367 11549 6401
rect 11587 6367 11608 6401
rect 11608 6367 11621 6401
rect 11659 6367 11676 6401
rect 11676 6367 11693 6401
rect 11731 6367 11744 6401
rect 11744 6367 11765 6401
rect 11803 6367 11812 6401
rect 11812 6367 11837 6401
rect 11875 6367 11880 6401
rect 11880 6367 11909 6401
rect 11947 6367 11948 6401
rect 11948 6367 11981 6401
rect 12019 6367 12050 6401
rect 12050 6367 12053 6401
rect 12091 6367 12118 6401
rect 12118 6367 12125 6401
rect 12163 6367 12186 6401
rect 12186 6367 12197 6401
rect 12235 6367 12254 6401
rect 12254 6367 12269 6401
rect 12307 6367 12322 6401
rect 12322 6367 12341 6401
rect 12379 6367 12390 6401
rect 12390 6367 12413 6401
rect 12451 6367 12458 6401
rect 12458 6367 12485 6401
rect 12523 6367 12526 6401
rect 12526 6367 12557 6401
rect 12595 6367 12628 6401
rect 12628 6367 12629 6401
rect 12667 6367 12696 6401
rect 12696 6367 12701 6401
rect 12739 6367 12764 6401
rect 12764 6367 12773 6401
rect 12811 6367 12832 6401
rect 12832 6367 12845 6401
rect 12883 6367 12900 6401
rect 12900 6367 12917 6401
rect 12955 6367 12968 6401
rect 12968 6367 12989 6401
rect 13027 6367 13036 6401
rect 13036 6367 13061 6401
rect 13099 6367 13104 6401
rect 13104 6367 13133 6401
rect 13171 6367 13172 6401
rect 13172 6367 13205 6401
rect 13243 6367 13274 6401
rect 13274 6367 13277 6401
rect 13315 6367 13342 6401
rect 13342 6367 13349 6401
rect 13595 8082 13600 8096
rect 13600 8082 13629 8096
rect 13595 8062 13629 8082
rect 13667 8062 13701 8096
rect 13739 8086 13766 8096
rect 13766 8086 13773 8096
rect 13739 8062 13773 8086
rect 13595 8014 13600 8022
rect 13600 8014 13629 8022
rect 13595 7988 13629 8014
rect 13667 7988 13701 8022
rect 13739 8018 13766 8022
rect 13766 8018 13773 8022
rect 13739 7988 13773 8018
rect 13595 7946 13600 7948
rect 13600 7946 13629 7948
rect 13595 7914 13629 7946
rect 13667 7914 13701 7948
rect 13739 7916 13773 7948
rect 13739 7914 13766 7916
rect 13766 7914 13773 7916
rect 13595 7844 13629 7874
rect 13595 7840 13600 7844
rect 13600 7840 13629 7844
rect 13667 7840 13701 7874
rect 13739 7848 13773 7874
rect 13739 7840 13766 7848
rect 13766 7840 13773 7848
rect 13595 7776 13629 7800
rect 13595 7766 13600 7776
rect 13600 7766 13629 7776
rect 13667 7766 13701 7800
rect 13739 7780 13773 7800
rect 13739 7766 13766 7780
rect 13766 7766 13773 7780
rect 13595 7708 13629 7726
rect 13595 7692 13600 7708
rect 13600 7692 13629 7708
rect 13667 7692 13701 7726
rect 13739 7712 13773 7726
rect 13739 7692 13766 7712
rect 13766 7692 13773 7712
rect 13595 7640 13629 7652
rect 13595 7618 13600 7640
rect 13600 7618 13629 7640
rect 13667 7618 13701 7652
rect 13739 7644 13773 7652
rect 13739 7618 13766 7644
rect 13766 7618 13773 7644
rect 13595 7572 13629 7578
rect 13595 7544 13600 7572
rect 13600 7544 13629 7572
rect 13667 7544 13701 7578
rect 13739 7576 13773 7578
rect 13739 7544 13766 7576
rect 13766 7544 13773 7576
rect 13595 7470 13600 7504
rect 13600 7470 13629 7504
rect 13667 7470 13701 7504
rect 13739 7474 13766 7504
rect 13766 7474 13773 7504
rect 13739 7470 13773 7474
rect 13595 7402 13600 7430
rect 13600 7402 13629 7430
rect 13595 7396 13629 7402
rect 13667 7397 13701 7431
rect 13739 7406 13766 7431
rect 13766 7406 13773 7431
rect 13739 7397 13773 7406
rect 13595 7334 13600 7356
rect 13600 7334 13629 7356
rect 13595 7322 13629 7334
rect 13667 7324 13701 7358
rect 13739 7338 13766 7358
rect 13766 7338 13773 7358
rect 13739 7324 13773 7338
rect 13595 7266 13600 7283
rect 13600 7266 13629 7283
rect 13595 7249 13629 7266
rect 13667 7251 13701 7285
rect 13739 7270 13766 7285
rect 13766 7270 13773 7285
rect 13739 7251 13773 7270
rect 13595 7198 13600 7210
rect 13600 7198 13629 7210
rect 13595 7176 13629 7198
rect 13667 7178 13701 7212
rect 13739 7202 13766 7212
rect 13766 7202 13773 7212
rect 13739 7178 13773 7202
rect 13595 7130 13600 7137
rect 13600 7130 13629 7137
rect 13595 7103 13629 7130
rect 13667 7105 13701 7139
rect 13739 7134 13766 7139
rect 13766 7134 13773 7139
rect 13739 7105 13773 7134
rect 13595 7062 13600 7064
rect 13600 7062 13629 7064
rect 13595 7030 13629 7062
rect 13667 7032 13701 7066
rect 13739 7032 13773 7066
rect 13595 6960 13629 6991
rect 13595 6957 13600 6960
rect 13600 6957 13629 6960
rect 13667 6959 13701 6993
rect 13739 6964 13773 6993
rect 13739 6959 13766 6964
rect 13766 6959 13773 6964
rect 13595 6892 13629 6918
rect 13595 6884 13600 6892
rect 13600 6884 13629 6892
rect 13667 6886 13701 6920
rect 13739 6896 13773 6920
rect 13739 6886 13766 6896
rect 13766 6886 13773 6896
rect 13595 6824 13629 6845
rect 13595 6811 13600 6824
rect 13600 6811 13629 6824
rect 13667 6813 13701 6847
rect 13739 6828 13773 6847
rect 13739 6813 13766 6828
rect 13766 6813 13773 6828
rect 13595 6756 13629 6772
rect 13595 6738 13600 6756
rect 13600 6738 13629 6756
rect 13667 6740 13701 6774
rect 13739 6760 13773 6774
rect 13739 6740 13766 6760
rect 13766 6740 13773 6760
rect 13595 6688 13629 6699
rect 13595 6665 13600 6688
rect 13600 6665 13629 6688
rect 13667 6667 13701 6701
rect 13739 6692 13773 6701
rect 13739 6667 13766 6692
rect 13766 6667 13773 6692
rect 13595 6620 13629 6626
rect 13595 6592 13600 6620
rect 13600 6592 13629 6620
rect 13667 6594 13701 6628
rect 13739 6624 13773 6628
rect 13739 6594 13766 6624
rect 13766 6594 13773 6624
rect 13595 6552 13629 6553
rect 13595 6519 13600 6552
rect 13600 6519 13629 6552
rect 13667 6521 13701 6555
rect 13739 6522 13766 6555
rect 13766 6522 13773 6555
rect 13739 6521 13773 6522
rect 13595 6450 13600 6480
rect 13600 6450 13629 6480
rect 13595 6446 13629 6450
rect 13667 6448 13701 6482
rect 13739 6454 13766 6482
rect 13766 6454 13773 6482
rect 13739 6448 13773 6454
rect 13595 6382 13600 6407
rect 13600 6382 13629 6407
rect 13595 6373 13629 6382
rect 13667 6375 13701 6409
rect 13739 6386 13766 6409
rect 13766 6386 13773 6409
rect 13739 6375 13773 6386
rect 10464 6329 10498 6350
rect 10464 6316 10473 6329
rect 10473 6316 10498 6329
rect 10536 6316 10570 6350
rect 10608 6329 10642 6348
rect 10608 6314 10639 6329
rect 10639 6314 10642 6329
rect 10464 6261 10498 6272
rect 10464 6238 10473 6261
rect 10473 6238 10498 6261
rect 10536 6238 10570 6272
rect 10608 6234 10642 6268
rect 13595 6314 13600 6334
rect 13600 6314 13629 6334
rect 13595 6300 13629 6314
rect 13667 6302 13701 6336
rect 13739 6318 13766 6336
rect 13766 6318 13773 6336
rect 13739 6302 13773 6318
rect 13595 6246 13600 6261
rect 13600 6246 13629 6261
rect 13595 6227 13629 6246
rect 13667 6229 13701 6263
rect 13739 6250 13766 6263
rect 13766 6250 13773 6263
rect 13739 6229 13773 6250
rect 10464 6193 10498 6194
rect 10464 6160 10473 6193
rect 10473 6160 10498 6193
rect 10536 6160 10570 6194
rect 10608 6178 10639 6188
rect 10639 6178 10673 6188
rect 10673 6178 10707 6188
rect 10707 6178 10741 6188
rect 10741 6178 10775 6188
rect 10775 6178 10809 6188
rect 10809 6178 10843 6188
rect 10843 6178 10877 6188
rect 10877 6178 10911 6188
rect 10911 6178 10945 6188
rect 10945 6178 10979 6188
rect 10979 6178 11013 6188
rect 11013 6178 11047 6188
rect 11047 6178 11074 6188
rect 11113 6178 11115 6188
rect 11115 6178 11147 6188
rect 11186 6178 11217 6188
rect 11217 6178 11220 6188
rect 11259 6178 11285 6188
rect 11285 6178 11293 6188
rect 11332 6178 11353 6188
rect 11353 6178 11366 6188
rect 11405 6178 11421 6188
rect 11421 6178 11439 6188
rect 11478 6178 11489 6188
rect 11489 6178 11512 6188
rect 11551 6178 11557 6188
rect 11557 6178 11585 6188
rect 11624 6178 11625 6188
rect 11625 6178 11658 6188
rect 11697 6178 11727 6188
rect 11727 6178 11731 6188
rect 11770 6178 11795 6188
rect 11795 6178 11804 6188
rect 11843 6178 11863 6188
rect 11863 6178 11877 6188
rect 11916 6178 11931 6188
rect 11931 6178 11950 6188
rect 11989 6178 11999 6188
rect 11999 6178 12023 6188
rect 12062 6178 12067 6188
rect 12067 6178 12096 6188
rect 10608 6116 11074 6178
rect 11113 6154 11147 6178
rect 11186 6154 11220 6178
rect 11259 6154 11293 6178
rect 11332 6154 11366 6178
rect 11405 6154 11439 6178
rect 11478 6154 11512 6178
rect 11551 6154 11585 6178
rect 11624 6154 11658 6178
rect 11697 6154 11731 6178
rect 11770 6154 11804 6178
rect 11843 6154 11877 6178
rect 11916 6154 11950 6178
rect 11989 6154 12023 6178
rect 12062 6154 12096 6178
rect 12135 6154 12169 6188
rect 12208 6178 12237 6188
rect 12237 6178 12242 6188
rect 12281 6178 12305 6188
rect 12305 6178 12315 6188
rect 12354 6178 12373 6188
rect 12373 6178 12388 6188
rect 12427 6178 12441 6188
rect 12441 6178 12461 6188
rect 12500 6178 12509 6188
rect 12509 6178 12534 6188
rect 12573 6178 12577 6188
rect 12577 6178 12607 6188
rect 12646 6178 12679 6188
rect 12679 6178 12680 6188
rect 12719 6178 12747 6188
rect 12747 6178 12753 6188
rect 12792 6178 12815 6188
rect 12815 6178 12826 6188
rect 12865 6178 12883 6188
rect 12883 6178 12899 6188
rect 12938 6178 12951 6188
rect 12951 6178 12972 6188
rect 13011 6178 13019 6188
rect 13019 6178 13045 6188
rect 13084 6178 13087 6188
rect 13087 6178 13118 6188
rect 13157 6178 13189 6188
rect 13189 6178 13191 6188
rect 13230 6178 13257 6188
rect 13257 6178 13264 6188
rect 13303 6178 13325 6188
rect 13325 6178 13337 6188
rect 13376 6178 13393 6188
rect 13393 6178 13410 6188
rect 13449 6178 13461 6188
rect 13461 6178 13483 6188
rect 13522 6178 13529 6188
rect 13529 6178 13556 6188
rect 13595 6178 13600 6188
rect 13600 6178 13629 6188
rect 12208 6154 12242 6178
rect 12281 6154 12315 6178
rect 12354 6154 12388 6178
rect 12427 6154 12461 6178
rect 12500 6154 12534 6178
rect 12573 6154 12607 6178
rect 12646 6154 12680 6178
rect 12719 6154 12753 6178
rect 12792 6154 12826 6178
rect 12865 6154 12899 6178
rect 12938 6154 12972 6178
rect 13011 6154 13045 6178
rect 13084 6154 13118 6178
rect 13157 6154 13191 6178
rect 13230 6154 13264 6178
rect 13303 6154 13337 6178
rect 13376 6154 13410 6178
rect 13449 6154 13483 6178
rect 13522 6154 13556 6178
rect 13595 6154 13629 6178
rect 13667 6156 13701 6190
rect 13739 6182 13766 6190
rect 13766 6182 13773 6190
rect 13739 6156 13773 6182
rect 10464 6082 10498 6116
rect 10536 6080 11146 6116
rect 11185 6082 11219 6116
rect 11258 6082 11292 6116
rect 11331 6082 11365 6116
rect 11404 6082 11438 6116
rect 11477 6082 11511 6116
rect 11550 6082 11584 6116
rect 11623 6082 11657 6116
rect 11696 6082 11730 6116
rect 11769 6082 11803 6116
rect 11842 6082 11876 6116
rect 11915 6082 11949 6116
rect 11988 6082 12022 6116
rect 12061 6082 12095 6116
rect 12134 6082 12168 6116
rect 12207 6082 12241 6116
rect 12280 6082 12314 6116
rect 12353 6082 12387 6116
rect 12426 6082 12460 6116
rect 12499 6082 12533 6116
rect 12572 6082 12606 6116
rect 12645 6082 12679 6116
rect 12718 6082 12752 6116
rect 12791 6082 12825 6116
rect 12864 6082 12898 6116
rect 12937 6082 12971 6116
rect 13010 6082 13044 6116
rect 13083 6082 13117 6116
rect 13156 6082 13190 6116
rect 13229 6082 13263 6116
rect 13302 6082 13336 6116
rect 13375 6082 13409 6116
rect 13448 6082 13482 6116
rect 13521 6082 13555 6116
rect 13594 6082 13628 6116
rect 13667 6082 13701 6116
rect 13739 6114 13766 6117
rect 13766 6114 13773 6117
rect 13739 6083 13773 6114
rect 10536 6046 10541 6080
rect 10541 6046 10575 6080
rect 10575 6046 10609 6080
rect 10609 6046 10643 6080
rect 10643 6046 10677 6080
rect 10677 6046 10711 6080
rect 10711 6046 10745 6080
rect 10745 6046 10779 6080
rect 10779 6046 10813 6080
rect 10813 6046 10847 6080
rect 10847 6046 10881 6080
rect 10881 6046 10915 6080
rect 10915 6046 10949 6080
rect 10949 6046 10983 6080
rect 10983 6046 11017 6080
rect 11017 6046 11051 6080
rect 11051 6046 11085 6080
rect 11085 6046 11119 6080
rect 11119 6046 11146 6080
rect 10536 6010 11146 6046
rect 11185 6010 11219 6044
rect 11258 6010 11292 6044
rect 11331 6010 11365 6044
rect 11404 6010 11438 6044
rect 11477 6010 11511 6044
rect 11550 6010 11584 6044
rect 11623 6010 11657 6044
rect 11696 6010 11730 6044
rect 11769 6010 11803 6044
rect 11842 6010 11876 6044
rect 11915 6010 11949 6044
rect 11988 6010 12022 6044
rect 12061 6010 12095 6044
rect 12134 6010 12168 6044
rect 12207 6010 12241 6044
rect 12280 6010 12314 6044
rect 12353 6010 12387 6044
rect 12426 6010 12460 6044
rect 12499 6010 12533 6044
rect 12572 6010 12606 6044
rect 12645 6010 12679 6044
rect 12718 6010 12752 6044
rect 12791 6010 12825 6044
rect 12864 6010 12898 6044
rect 12937 6010 12971 6044
rect 13010 6010 13044 6044
rect 13083 6010 13117 6044
rect 13156 6010 13190 6044
rect 13229 6010 13263 6044
rect 13302 6010 13336 6044
rect 13375 6010 13409 6044
rect 13448 6010 13482 6044
rect 13521 6010 13555 6044
rect 13594 6010 13628 6044
rect 13667 6010 13701 6044
rect 10473 5916 10507 5950
rect 10546 5916 10580 5950
rect 10619 5916 10653 5950
rect 10692 5916 10726 5950
rect 10765 5916 10799 5950
rect 10838 5916 10872 5950
rect 10911 5916 10945 5950
rect 10984 5916 11018 5950
rect 11057 5916 11091 5950
rect 11130 5916 11164 5950
rect 11203 5916 11237 5950
rect 11276 5916 11310 5950
rect 11349 5916 11383 5950
rect 11422 5916 11456 5950
rect 11495 5916 11529 5950
rect 11568 5916 11602 5950
rect 11641 5916 11675 5950
rect 11714 5916 11748 5950
rect 11787 5916 11821 5950
rect 11860 5916 11894 5950
rect 11933 5916 11967 5950
rect 12005 5916 12039 5950
rect 12077 5916 12111 5950
rect 12149 5916 12183 5950
rect 12221 5916 12255 5950
rect 12293 5916 12327 5950
rect 12365 5916 12399 5950
rect 12437 5916 12471 5950
rect 12509 5916 12543 5950
rect 12581 5916 12615 5950
rect 12653 5916 12687 5950
rect 12725 5916 12759 5950
rect 12797 5916 12831 5950
rect 12869 5916 12903 5950
rect 12941 5916 12975 5950
rect 13013 5916 13047 5950
rect 13085 5916 13119 5950
rect 13157 5916 13191 5950
rect 13229 5916 13263 5950
rect 13301 5916 13335 5950
rect 13373 5916 13407 5950
rect 13445 5916 13479 5950
rect 13517 5916 13551 5950
rect 13589 5916 13623 5950
rect 13661 5916 13695 5950
rect 13733 5916 13767 5950
rect 1019 5852 1049 5880
rect 1049 5852 1053 5880
rect 1092 5852 1117 5880
rect 1117 5852 1126 5880
rect 1165 5852 1185 5880
rect 1185 5852 1199 5880
rect 1237 5852 1253 5880
rect 1253 5852 1271 5880
rect 1309 5852 1321 5880
rect 1321 5852 1343 5880
rect 1381 5852 1389 5880
rect 1389 5852 1415 5880
rect 1453 5852 1457 5880
rect 1457 5852 1487 5880
rect 1019 5846 1053 5852
rect 1092 5846 1126 5852
rect 1165 5846 1199 5852
rect 1237 5846 1271 5852
rect 1309 5846 1343 5852
rect 1381 5846 1415 5852
rect 1453 5846 1487 5852
rect 1525 5846 1559 5880
rect 1597 5852 1627 5880
rect 1627 5852 1631 5880
rect 1669 5852 1695 5880
rect 1695 5852 1703 5880
rect 1741 5852 1763 5880
rect 1763 5852 1775 5880
rect 1813 5852 1831 5880
rect 1831 5852 1847 5880
rect 1885 5852 1899 5880
rect 1899 5852 1919 5880
rect 1957 5852 1967 5880
rect 1967 5852 1991 5880
rect 2029 5852 2035 5880
rect 2035 5852 2063 5880
rect 2101 5852 2103 5880
rect 2103 5852 2135 5880
rect 2173 5852 2205 5880
rect 2205 5852 2207 5880
rect 2245 5852 2273 5880
rect 2273 5852 2279 5880
rect 2317 5852 2341 5880
rect 2341 5852 2351 5880
rect 2389 5852 2409 5880
rect 2409 5852 2423 5880
rect 2461 5852 2477 5880
rect 2477 5852 2495 5880
rect 2533 5852 2545 5880
rect 2545 5852 2567 5880
rect 2605 5852 2613 5880
rect 2613 5852 2639 5880
rect 2677 5852 2681 5880
rect 2681 5852 2711 5880
rect 1597 5846 1631 5852
rect 1669 5846 1703 5852
rect 1741 5846 1775 5852
rect 1813 5846 1847 5852
rect 1885 5846 1919 5852
rect 1957 5846 1991 5852
rect 2029 5846 2063 5852
rect 2101 5846 2135 5852
rect 2173 5846 2207 5852
rect 2245 5846 2279 5852
rect 2317 5846 2351 5852
rect 2389 5846 2423 5852
rect 2461 5846 2495 5852
rect 2533 5846 2567 5852
rect 2605 5846 2639 5852
rect 2677 5846 2711 5852
rect 2749 5846 2783 5880
rect 2821 5852 2851 5880
rect 2851 5852 2855 5880
rect 2893 5852 2919 5880
rect 2919 5852 2927 5880
rect 2965 5852 2987 5880
rect 2987 5852 2999 5880
rect 3037 5852 3055 5880
rect 3055 5852 3071 5880
rect 3109 5852 3123 5880
rect 3123 5852 3143 5880
rect 3181 5852 3191 5880
rect 3191 5852 3215 5880
rect 3253 5852 3259 5880
rect 3259 5852 3287 5880
rect 3325 5852 3327 5880
rect 3327 5852 3359 5880
rect 3397 5852 3429 5880
rect 3429 5852 3431 5880
rect 3469 5852 3497 5880
rect 3497 5852 3503 5880
rect 3541 5852 3565 5880
rect 3565 5852 3575 5880
rect 3613 5852 3633 5880
rect 3633 5852 3647 5880
rect 3685 5852 3701 5880
rect 3701 5852 3719 5880
rect 3757 5852 3769 5880
rect 3769 5852 3791 5880
rect 3829 5852 3837 5880
rect 3837 5852 3863 5880
rect 3901 5852 3905 5880
rect 3905 5852 3935 5880
rect 2821 5846 2855 5852
rect 2893 5846 2927 5852
rect 2965 5846 2999 5852
rect 3037 5846 3071 5852
rect 3109 5846 3143 5852
rect 3181 5846 3215 5852
rect 3253 5846 3287 5852
rect 3325 5846 3359 5852
rect 3397 5846 3431 5852
rect 3469 5846 3503 5852
rect 3541 5846 3575 5852
rect 3613 5846 3647 5852
rect 3685 5846 3719 5852
rect 3757 5846 3791 5852
rect 3829 5846 3863 5852
rect 3901 5846 3935 5852
rect 3973 5846 4007 5880
rect 4045 5852 4075 5880
rect 4075 5852 4079 5880
rect 4117 5852 4143 5880
rect 4143 5852 4151 5880
rect 4189 5852 4211 5880
rect 4211 5852 4223 5880
rect 4261 5852 4279 5880
rect 4279 5852 4295 5880
rect 4333 5852 4347 5880
rect 4347 5852 4367 5880
rect 4405 5852 4415 5880
rect 4415 5852 4439 5880
rect 4477 5852 4483 5880
rect 4483 5852 4511 5880
rect 4549 5852 4551 5880
rect 4551 5852 4583 5880
rect 4621 5852 4653 5880
rect 4653 5852 4655 5880
rect 4693 5852 4721 5880
rect 4721 5852 4727 5880
rect 4765 5852 4789 5880
rect 4789 5852 4799 5880
rect 4837 5852 4857 5880
rect 4857 5852 4871 5880
rect 4909 5852 4925 5880
rect 4925 5852 4943 5880
rect 4981 5852 4993 5880
rect 4993 5852 5015 5880
rect 5053 5852 5061 5880
rect 5061 5852 5087 5880
rect 5125 5852 5129 5880
rect 5129 5852 5159 5880
rect 4045 5846 4079 5852
rect 4117 5846 4151 5852
rect 4189 5846 4223 5852
rect 4261 5846 4295 5852
rect 4333 5846 4367 5852
rect 4405 5846 4439 5852
rect 4477 5846 4511 5852
rect 4549 5846 4583 5852
rect 4621 5846 4655 5852
rect 4693 5846 4727 5852
rect 4765 5846 4799 5852
rect 4837 5846 4871 5852
rect 4909 5846 4943 5852
rect 4981 5846 5015 5852
rect 5053 5846 5087 5852
rect 5125 5846 5159 5852
rect 5197 5846 5231 5880
rect 5269 5852 5299 5880
rect 5299 5852 5303 5880
rect 5341 5852 5367 5880
rect 5367 5852 5375 5880
rect 5413 5852 5435 5880
rect 5435 5852 5447 5880
rect 5485 5852 5503 5880
rect 5503 5852 5519 5880
rect 5557 5852 5571 5880
rect 5571 5852 5591 5880
rect 5629 5852 5639 5880
rect 5639 5852 5663 5880
rect 5701 5852 5707 5880
rect 5707 5852 5735 5880
rect 5773 5852 5775 5880
rect 5775 5852 5807 5880
rect 5845 5852 5877 5880
rect 5877 5852 5879 5880
rect 5917 5852 5945 5880
rect 5945 5852 5951 5880
rect 5989 5852 6013 5880
rect 6013 5852 6023 5880
rect 6061 5852 6081 5880
rect 6081 5852 6095 5880
rect 6133 5852 6149 5880
rect 6149 5852 6167 5880
rect 6205 5852 6217 5880
rect 6217 5852 6239 5880
rect 6277 5852 6285 5880
rect 6285 5852 6311 5880
rect 6349 5852 6353 5880
rect 6353 5852 6383 5880
rect 5269 5846 5303 5852
rect 5341 5846 5375 5852
rect 5413 5846 5447 5852
rect 5485 5846 5519 5852
rect 5557 5846 5591 5852
rect 5629 5846 5663 5852
rect 5701 5846 5735 5852
rect 5773 5846 5807 5852
rect 5845 5846 5879 5852
rect 5917 5846 5951 5852
rect 5989 5846 6023 5852
rect 6061 5846 6095 5852
rect 6133 5846 6167 5852
rect 6205 5846 6239 5852
rect 6277 5846 6311 5852
rect 6349 5846 6383 5852
rect 6421 5846 6455 5880
rect 6493 5852 6523 5880
rect 6523 5852 6527 5880
rect 6565 5852 6591 5880
rect 6591 5852 6599 5880
rect 6637 5852 6659 5880
rect 6659 5852 6671 5880
rect 6709 5852 6727 5880
rect 6727 5852 6743 5880
rect 6781 5852 6795 5880
rect 6795 5852 6815 5880
rect 6853 5852 6863 5880
rect 6863 5852 6887 5880
rect 6925 5852 6931 5880
rect 6931 5852 6959 5880
rect 6997 5852 6999 5880
rect 6999 5852 7031 5880
rect 7069 5852 7101 5880
rect 7101 5852 7103 5880
rect 7141 5852 7169 5880
rect 7169 5852 7175 5880
rect 7213 5852 7237 5880
rect 7237 5852 7247 5880
rect 7285 5852 7305 5880
rect 7305 5852 7319 5880
rect 7357 5852 7373 5880
rect 7373 5852 7391 5880
rect 7429 5852 7441 5880
rect 7441 5852 7463 5880
rect 7501 5852 7509 5880
rect 7509 5852 7535 5880
rect 7573 5852 7577 5880
rect 7577 5852 7607 5880
rect 6493 5846 6527 5852
rect 6565 5846 6599 5852
rect 6637 5846 6671 5852
rect 6709 5846 6743 5852
rect 6781 5846 6815 5852
rect 6853 5846 6887 5852
rect 6925 5846 6959 5852
rect 6997 5846 7031 5852
rect 7069 5846 7103 5852
rect 7141 5846 7175 5852
rect 7213 5846 7247 5852
rect 7285 5846 7319 5852
rect 7357 5846 7391 5852
rect 7429 5846 7463 5852
rect 7501 5846 7535 5852
rect 7573 5846 7607 5852
rect 7645 5846 7679 5880
rect 7717 5852 7747 5880
rect 7747 5852 7751 5880
rect 7789 5852 7815 5880
rect 7815 5852 7823 5880
rect 7861 5852 7883 5880
rect 7883 5852 7895 5880
rect 7933 5852 7951 5880
rect 7951 5852 7967 5880
rect 8005 5852 8019 5880
rect 8019 5852 8039 5880
rect 8077 5852 8087 5880
rect 8087 5852 8111 5880
rect 8149 5852 8155 5880
rect 8155 5852 8183 5880
rect 8221 5852 8223 5880
rect 8223 5852 8255 5880
rect 8293 5852 8325 5880
rect 8325 5852 8327 5880
rect 8365 5852 8393 5880
rect 8393 5852 8399 5880
rect 8437 5852 8461 5880
rect 8461 5852 8471 5880
rect 8509 5852 8529 5880
rect 8529 5852 8543 5880
rect 8581 5852 8597 5880
rect 8597 5852 8615 5880
rect 8653 5852 8665 5880
rect 8665 5852 8687 5880
rect 8725 5852 8733 5880
rect 8733 5852 8759 5880
rect 8797 5852 8801 5880
rect 8801 5852 8831 5880
rect 7717 5846 7751 5852
rect 7789 5846 7823 5852
rect 7861 5846 7895 5852
rect 7933 5846 7967 5852
rect 8005 5846 8039 5852
rect 8077 5846 8111 5852
rect 8149 5846 8183 5852
rect 8221 5846 8255 5852
rect 8293 5846 8327 5852
rect 8365 5846 8399 5852
rect 8437 5846 8471 5852
rect 8509 5846 8543 5852
rect 8581 5846 8615 5852
rect 8653 5846 8687 5852
rect 8725 5846 8759 5852
rect 8797 5846 8831 5852
rect 8869 5846 8903 5880
rect 8941 5852 8971 5880
rect 8971 5852 8975 5880
rect 9013 5852 9039 5880
rect 9039 5852 9047 5880
rect 8941 5846 8975 5852
rect 9013 5846 9047 5852
rect 9085 5846 9119 5880
rect 770 5791 790 5825
rect 790 5791 804 5825
rect 626 5719 660 5753
rect 698 5719 732 5753
rect 770 5718 790 5752
rect 790 5718 804 5752
rect 626 5646 660 5680
rect 698 5646 732 5680
rect 770 5645 804 5679
rect 626 5597 654 5607
rect 654 5597 660 5607
rect 698 5597 722 5607
rect 722 5597 732 5607
rect 9462 5809 9466 5843
rect 9466 5809 9496 5843
rect 9534 5809 9568 5843
rect 9606 5809 9636 5843
rect 9636 5809 9640 5843
rect 9462 5730 9466 5764
rect 9466 5730 9496 5764
rect 9534 5732 9568 5766
rect 9606 5732 9636 5766
rect 9636 5732 9640 5766
rect 9462 5651 9466 5685
rect 9466 5651 9496 5685
rect 9534 5656 9568 5690
rect 9606 5656 9636 5690
rect 9636 5656 9640 5690
rect 770 5602 5700 5606
rect 5739 5602 5773 5606
rect 5812 5602 5846 5606
rect 5885 5602 5919 5606
rect 5958 5602 5992 5606
rect 6031 5602 6065 5606
rect 6104 5602 6138 5606
rect 6177 5602 6211 5606
rect 6250 5602 6284 5606
rect 6323 5602 6357 5606
rect 6396 5602 6430 5606
rect 6469 5602 6503 5606
rect 6542 5602 6576 5606
rect 6615 5602 6649 5606
rect 6688 5602 6722 5606
rect 6761 5602 6795 5606
rect 6834 5602 6868 5606
rect 6907 5602 6941 5606
rect 6980 5602 7014 5606
rect 7053 5602 7087 5606
rect 7126 5602 7160 5606
rect 7199 5602 7233 5606
rect 7272 5602 7306 5606
rect 7345 5602 7379 5606
rect 7418 5602 7452 5606
rect 7491 5602 7525 5606
rect 7564 5602 7598 5606
rect 7637 5602 7671 5606
rect 7710 5602 7744 5606
rect 7783 5602 7817 5606
rect 7856 5602 7890 5606
rect 7929 5602 7963 5606
rect 8002 5602 8036 5606
rect 8075 5602 8109 5606
rect 8148 5602 8182 5606
rect 8221 5602 8255 5606
rect 8294 5602 8328 5606
rect 8367 5602 8401 5606
rect 8440 5602 8474 5606
rect 8513 5602 8547 5606
rect 8586 5602 8620 5606
rect 8659 5602 8693 5606
rect 8732 5602 8766 5606
rect 8805 5602 8839 5606
rect 8878 5602 8912 5606
rect 8951 5602 8985 5606
rect 9024 5602 9058 5606
rect 9097 5602 9131 5606
rect 9170 5602 9204 5606
rect 9243 5602 9277 5606
rect 9316 5602 9350 5606
rect 9389 5602 9423 5606
rect 626 5573 660 5597
rect 698 5573 732 5597
rect 770 5534 5700 5602
rect 5739 5572 5773 5602
rect 5812 5572 5846 5602
rect 5885 5572 5919 5602
rect 5958 5572 5992 5602
rect 6031 5572 6065 5602
rect 6104 5572 6138 5602
rect 6177 5572 6211 5602
rect 6250 5572 6284 5602
rect 6323 5572 6357 5602
rect 6396 5572 6430 5602
rect 6469 5572 6503 5602
rect 6542 5572 6576 5602
rect 6615 5572 6649 5602
rect 6688 5572 6722 5602
rect 6761 5572 6795 5602
rect 6834 5572 6868 5602
rect 6907 5572 6941 5602
rect 6980 5572 7014 5602
rect 7053 5572 7087 5602
rect 7126 5572 7160 5602
rect 7199 5572 7233 5602
rect 7272 5572 7306 5602
rect 7345 5572 7379 5602
rect 7418 5572 7452 5602
rect 7491 5572 7525 5602
rect 7564 5572 7598 5602
rect 7637 5572 7671 5602
rect 7710 5572 7744 5602
rect 7783 5572 7817 5602
rect 7856 5572 7890 5602
rect 7929 5572 7963 5602
rect 8002 5572 8036 5602
rect 8075 5572 8109 5602
rect 8148 5572 8182 5602
rect 8221 5572 8255 5602
rect 8294 5572 8328 5602
rect 8367 5572 8401 5602
rect 8440 5572 8474 5602
rect 8513 5572 8547 5602
rect 8586 5572 8620 5602
rect 8659 5572 8693 5602
rect 8732 5572 8766 5602
rect 8805 5572 8839 5602
rect 8878 5572 8912 5602
rect 8951 5572 8985 5602
rect 9024 5572 9058 5602
rect 9097 5572 9131 5602
rect 9170 5572 9204 5602
rect 9243 5572 9277 5602
rect 9316 5572 9350 5602
rect 9389 5572 9423 5602
rect 9462 5572 9466 5606
rect 9466 5572 9496 5606
rect 9534 5580 9568 5614
rect 9606 5580 9636 5614
rect 9636 5580 9640 5614
rect 626 5529 654 5534
rect 654 5529 660 5534
rect 626 5500 660 5529
rect 698 5432 5772 5534
rect 5811 5500 5845 5534
rect 5884 5500 5918 5534
rect 5957 5500 5991 5534
rect 6030 5500 6064 5534
rect 6103 5500 6137 5534
rect 6176 5500 6210 5534
rect 6249 5500 6283 5534
rect 6322 5500 6356 5534
rect 6395 5500 6429 5534
rect 6468 5500 6502 5534
rect 6541 5500 6575 5534
rect 6614 5500 6648 5534
rect 6687 5500 6721 5534
rect 6760 5500 6794 5534
rect 6833 5500 6867 5534
rect 6906 5500 6940 5534
rect 6979 5500 7013 5534
rect 7052 5500 7086 5534
rect 7125 5500 7159 5534
rect 7198 5500 7232 5534
rect 7271 5500 7305 5534
rect 7344 5500 7378 5534
rect 7417 5500 7451 5534
rect 7490 5500 7524 5534
rect 7563 5500 7597 5534
rect 7636 5500 7670 5534
rect 7709 5500 7743 5534
rect 7782 5500 7816 5534
rect 7855 5500 7889 5534
rect 7928 5500 7962 5534
rect 8001 5500 8035 5534
rect 8074 5500 8108 5534
rect 8147 5500 8181 5534
rect 8220 5500 8254 5534
rect 8293 5500 8327 5534
rect 8366 5500 8400 5534
rect 8439 5500 8473 5534
rect 8512 5500 8546 5534
rect 8585 5500 8619 5534
rect 8658 5500 8692 5534
rect 8731 5500 8765 5534
rect 8804 5500 8838 5534
rect 8877 5500 8911 5534
rect 8950 5500 8984 5534
rect 9023 5500 9057 5534
rect 9096 5500 9130 5534
rect 9169 5500 9203 5534
rect 9242 5500 9276 5534
rect 9315 5500 9349 5534
rect 9388 5500 9422 5534
rect 9461 5500 9494 5534
rect 9494 5500 9495 5534
rect 9534 5500 9568 5534
rect 9606 5504 9636 5538
rect 9636 5504 9640 5538
rect 5811 5432 5845 5462
rect 5884 5432 5918 5462
rect 5957 5432 5991 5462
rect 6030 5432 6064 5462
rect 6103 5432 6137 5462
rect 6176 5432 6210 5462
rect 6249 5432 6283 5462
rect 6322 5432 6356 5462
rect 6395 5432 6429 5462
rect 6468 5432 6502 5462
rect 6541 5432 6575 5462
rect 6614 5432 6648 5462
rect 6687 5432 6721 5462
rect 6760 5432 6794 5462
rect 6833 5432 6867 5462
rect 6906 5432 6940 5462
rect 6979 5432 7013 5462
rect 7052 5432 7086 5462
rect 7125 5432 7159 5462
rect 7198 5432 7232 5462
rect 7271 5432 7305 5462
rect 7344 5432 7378 5462
rect 7417 5432 7451 5462
rect 7490 5432 7524 5462
rect 7563 5432 7597 5462
rect 7636 5432 7670 5462
rect 7709 5432 7743 5462
rect 7782 5432 7816 5462
rect 7855 5432 7889 5462
rect 7928 5432 7962 5462
rect 8001 5432 8035 5462
rect 8074 5432 8108 5462
rect 8147 5432 8181 5462
rect 8220 5432 8254 5462
rect 8293 5432 8327 5462
rect 8366 5432 8400 5462
rect 8439 5432 8473 5462
rect 8512 5432 8546 5462
rect 8585 5432 8619 5462
rect 8658 5432 8692 5462
rect 8731 5432 8765 5462
rect 8804 5432 8838 5462
rect 8877 5432 8911 5462
rect 8950 5432 8984 5462
rect 9023 5432 9057 5462
rect 9096 5432 9130 5462
rect 9169 5432 9203 5462
rect 9242 5432 9276 5462
rect 9315 5432 9349 5462
rect 9388 5432 9422 5462
rect 9461 5432 9494 5462
rect 9494 5432 9495 5462
rect 9534 5432 9562 5462
rect 9562 5432 9568 5462
rect 698 5428 5772 5432
rect 5811 5428 5845 5432
rect 5884 5428 5918 5432
rect 5957 5428 5991 5432
rect 6030 5428 6064 5432
rect 6103 5428 6137 5432
rect 6176 5428 6210 5432
rect 6249 5428 6283 5432
rect 6322 5428 6356 5432
rect 6395 5428 6429 5432
rect 6468 5428 6502 5432
rect 6541 5428 6575 5432
rect 6614 5428 6648 5432
rect 6687 5428 6721 5432
rect 6760 5428 6794 5432
rect 6833 5428 6867 5432
rect 6906 5428 6940 5432
rect 6979 5428 7013 5432
rect 7052 5428 7086 5432
rect 7125 5428 7159 5432
rect 7198 5428 7232 5432
rect 7271 5428 7305 5432
rect 7344 5428 7378 5432
rect 7417 5428 7451 5432
rect 7490 5428 7524 5432
rect 7563 5428 7597 5432
rect 7636 5428 7670 5432
rect 7709 5428 7743 5432
rect 7782 5428 7816 5432
rect 7855 5428 7889 5432
rect 7928 5428 7962 5432
rect 8001 5428 8035 5432
rect 8074 5428 8108 5432
rect 8147 5428 8181 5432
rect 8220 5428 8254 5432
rect 8293 5428 8327 5432
rect 8366 5428 8400 5432
rect 8439 5428 8473 5432
rect 8512 5428 8546 5432
rect 8585 5428 8619 5432
rect 8658 5428 8692 5432
rect 8731 5428 8765 5432
rect 8804 5428 8838 5432
rect 8877 5428 8911 5432
rect 8950 5428 8984 5432
rect 9023 5428 9057 5432
rect 9096 5428 9130 5432
rect 9169 5428 9203 5432
rect 9242 5428 9276 5432
rect 9315 5428 9349 5432
rect 9388 5428 9422 5432
rect 9461 5428 9495 5432
rect 9534 5428 9568 5432
rect 10904 5826 10964 5847
rect 10964 5826 10998 5847
rect 10998 5826 11032 5847
rect 10904 5792 11032 5826
rect 10832 5741 10836 5775
rect 10836 5741 10866 5775
rect 10904 5741 10938 5792
rect 10938 5758 11032 5792
rect 11032 5758 12594 5847
rect 12633 5813 12667 5847
rect 12706 5813 12740 5847
rect 12779 5813 12813 5847
rect 12852 5813 12886 5847
rect 12925 5813 12959 5847
rect 12998 5813 13032 5847
rect 13071 5813 13105 5847
rect 13144 5813 13178 5847
rect 13217 5813 13251 5847
rect 13290 5813 13324 5847
rect 13363 5813 13397 5847
rect 13436 5813 13470 5847
rect 13509 5813 13543 5847
rect 13582 5813 13616 5847
rect 13655 5813 13689 5847
rect 13728 5813 13762 5847
rect 13801 5813 13835 5847
rect 13874 5813 13908 5847
rect 13947 5813 13981 5847
rect 14020 5813 14054 5847
rect 10938 5741 11100 5758
rect 11100 5741 12594 5758
rect 12633 5741 12667 5775
rect 12706 5741 12740 5775
rect 12779 5741 12813 5775
rect 12852 5741 12886 5775
rect 12925 5741 12959 5775
rect 12998 5741 13032 5775
rect 13071 5741 13105 5775
rect 13144 5741 13178 5775
rect 13217 5741 13251 5775
rect 13290 5741 13324 5775
rect 13363 5741 13397 5775
rect 13436 5741 13470 5775
rect 13509 5741 13543 5775
rect 13582 5741 13616 5775
rect 13655 5741 13689 5775
rect 13728 5741 13762 5775
rect 13801 5741 13835 5775
rect 13874 5741 13908 5775
rect 13947 5741 13981 5775
rect 14020 5758 14058 5775
rect 14058 5758 14126 5775
rect 10976 5724 11100 5741
rect 10832 5665 10836 5699
rect 10836 5665 10866 5699
rect 10904 5666 10938 5700
rect 10976 5669 11006 5724
rect 11006 5690 11100 5724
rect 11100 5690 12522 5741
rect 14020 5746 14126 5758
rect 14020 5712 14092 5746
rect 14092 5712 14126 5746
rect 14020 5703 14126 5712
rect 12561 5690 12595 5703
rect 12634 5690 12668 5703
rect 12707 5690 12741 5703
rect 12780 5690 12814 5703
rect 12853 5690 12887 5703
rect 12926 5690 12960 5703
rect 12999 5690 13033 5703
rect 13072 5690 13106 5703
rect 13145 5690 13179 5703
rect 13218 5690 13252 5703
rect 13291 5690 13325 5703
rect 13364 5690 13398 5703
rect 13437 5690 13471 5703
rect 13510 5690 13544 5703
rect 13583 5690 13617 5703
rect 13656 5690 13690 5703
rect 13729 5690 13763 5703
rect 13802 5690 13836 5703
rect 13875 5690 13909 5703
rect 13948 5690 13990 5703
rect 13990 5690 14126 5703
rect 11006 5669 12522 5690
rect 12561 5669 12595 5690
rect 12634 5669 12668 5690
rect 12707 5669 12741 5690
rect 12780 5669 12814 5690
rect 12853 5669 12887 5690
rect 12926 5669 12960 5690
rect 12999 5669 13033 5690
rect 13072 5669 13106 5690
rect 13145 5669 13179 5690
rect 13218 5669 13252 5690
rect 13291 5669 13325 5690
rect 13364 5669 13398 5690
rect 13437 5669 13471 5690
rect 13510 5669 13544 5690
rect 13583 5669 13617 5690
rect 13656 5669 13690 5690
rect 13729 5669 13763 5690
rect 13802 5669 13836 5690
rect 13875 5669 13909 5690
rect 13948 5678 14126 5690
rect 10832 5589 10836 5623
rect 10836 5589 10866 5623
rect 10904 5591 10938 5625
rect 10976 5594 11006 5628
rect 11006 5594 11010 5628
rect 10832 5514 10836 5548
rect 10836 5514 10866 5548
rect 10904 5516 10938 5550
rect 10976 5519 11006 5553
rect 11006 5519 11010 5553
rect 13948 5610 14024 5678
rect 14024 5610 14126 5678
rect 10832 5439 10836 5473
rect 10836 5439 10866 5473
rect 10904 5441 10938 5475
rect 10976 5444 11006 5478
rect 11006 5444 11010 5478
rect 10832 5364 10836 5398
rect 10836 5364 10866 5398
rect 10904 5366 10938 5400
rect 10976 5369 11006 5403
rect 11006 5369 11010 5403
rect 10832 5289 10836 5323
rect 10836 5289 10866 5323
rect 10904 5291 10938 5325
rect 10976 5294 11006 5328
rect 11006 5294 11010 5328
rect 10832 5214 10836 5248
rect 10836 5214 10866 5248
rect 10904 5216 10938 5250
rect 10976 5219 11006 5253
rect 11006 5219 11010 5253
rect 10832 5139 10836 5173
rect 10836 5139 10866 5173
rect 10904 5141 10938 5175
rect 10976 5144 11006 5178
rect 11006 5144 11010 5178
rect 10832 5064 10836 5098
rect 10836 5064 10866 5098
rect 10904 5066 10938 5100
rect 10976 5069 11006 5103
rect 11006 5069 11010 5103
rect 10832 4989 10836 5023
rect 10836 4989 10866 5023
rect 10904 4991 10938 5025
rect 10976 4994 11006 5028
rect 11006 4994 11010 5028
rect 10832 4914 10836 4948
rect 10836 4914 10866 4948
rect 10904 4916 10938 4950
rect 10976 4919 11006 4953
rect 11006 4919 11010 4953
rect 10832 4839 10836 4873
rect 10836 4839 10866 4873
rect 10904 4841 10938 4875
rect 10976 4844 11006 4878
rect 11006 4844 11010 4878
rect 10832 4764 10836 4798
rect 10836 4764 10866 4798
rect 10904 4766 10938 4800
rect 10976 4769 11006 4803
rect 11006 4769 11010 4803
rect 10832 4689 10836 4723
rect 10836 4689 10866 4723
rect 10904 4692 10938 4726
rect 10976 4694 11006 4728
rect 11006 4694 11010 4728
rect 11468 5503 11502 5537
rect 11540 5503 11570 5537
rect 11570 5503 11574 5537
rect 11612 5503 11638 5537
rect 11638 5503 11646 5537
rect 11684 5503 11706 5537
rect 11706 5503 11718 5537
rect 11756 5503 11774 5537
rect 11774 5503 11790 5537
rect 11828 5503 11842 5537
rect 11842 5503 11862 5537
rect 11900 5503 11910 5537
rect 11910 5503 11934 5537
rect 11972 5503 11978 5537
rect 11978 5503 12006 5537
rect 12044 5503 12046 5537
rect 12046 5503 12078 5537
rect 12116 5503 12148 5537
rect 12148 5503 12150 5537
rect 12188 5503 12216 5537
rect 12216 5503 12222 5537
rect 12260 5503 12284 5537
rect 12284 5503 12294 5537
rect 12332 5503 12352 5537
rect 12352 5503 12366 5537
rect 12404 5503 12420 5537
rect 12420 5503 12438 5537
rect 12476 5503 12488 5537
rect 12488 5503 12510 5537
rect 11370 5449 11404 5462
rect 11370 5428 11404 5449
rect 11370 5381 11404 5390
rect 11370 5356 11404 5381
rect 11370 5313 11404 5318
rect 11370 5284 11404 5313
rect 12522 5449 12556 5462
rect 12522 5428 12556 5449
rect 12522 5381 12556 5390
rect 12522 5356 12556 5381
rect 11370 5245 11404 5246
rect 11370 5212 11404 5245
rect 11370 5143 11404 5174
rect 11370 5140 11404 5143
rect 11370 5075 11404 5102
rect 11370 5068 11404 5075
rect 11370 5007 11404 5030
rect 11370 4996 11404 5007
rect 11370 4939 11404 4958
rect 11370 4924 11404 4939
rect 11370 4871 11404 4886
rect 11370 4852 11404 4871
rect 11370 4803 11404 4814
rect 11370 4780 11404 4803
rect 11370 4735 11404 4742
rect 11370 4708 11404 4735
rect 2402 4616 10428 4648
rect 10467 4616 10501 4648
rect 10540 4616 10574 4648
rect 10613 4616 10647 4648
rect 10686 4616 10720 4648
rect 10759 4616 10793 4648
rect 10832 4616 10866 4648
rect 10904 4618 10938 4652
rect 10976 4619 11006 4653
rect 11006 4619 11010 4653
rect 2402 4582 2404 4616
rect 2404 4582 2438 4616
rect 2438 4582 2472 4616
rect 2330 4548 2364 4576
rect 2402 4548 2472 4582
rect 2472 4576 10428 4616
rect 10467 4614 10501 4616
rect 10540 4614 10574 4616
rect 10613 4614 10647 4616
rect 10686 4614 10720 4616
rect 10759 4614 10793 4616
rect 10832 4614 10866 4616
rect 2330 4542 2334 4548
rect 2334 4542 2364 4548
rect 2402 4542 2436 4548
rect 2436 4542 2472 4548
rect 2472 4542 10500 4576
rect 10539 4542 10573 4576
rect 10612 4542 10646 4576
rect 10685 4542 10719 4576
rect 10758 4542 10792 4576
rect 10831 4542 10865 4576
rect 10904 4548 10938 4576
rect 10976 4568 11010 4578
rect 10904 4542 10938 4548
rect 2474 4514 10500 4542
rect 2330 4469 2334 4503
rect 2334 4469 2364 4503
rect 2402 4469 2436 4503
rect 2474 4480 2540 4514
rect 2474 4470 2504 4480
rect 2504 4470 2540 4480
rect 2540 4470 10500 4514
rect 10976 4544 11006 4568
rect 11006 4544 11010 4568
rect 10539 4470 10573 4504
rect 10612 4470 10646 4504
rect 10685 4470 10719 4504
rect 10758 4470 10792 4504
rect 10831 4470 10865 4504
rect 10904 4470 10938 4504
rect 11517 5212 11551 5246
rect 11517 5140 11551 5174
rect 11517 5068 11551 5102
rect 11517 4996 11551 5030
rect 11517 4924 11551 4958
rect 11517 4852 11551 4886
rect 11517 4780 11551 4814
rect 11517 4708 11551 4742
rect 12376 5212 12410 5246
rect 12376 5140 12410 5174
rect 12376 5068 12410 5102
rect 12376 4996 12410 5030
rect 12376 4924 12410 4958
rect 12376 4852 12410 4886
rect 12376 4780 12410 4814
rect 12376 4708 12410 4742
rect 12522 5313 12556 5318
rect 12522 5284 12556 5313
rect 12522 5245 12556 5246
rect 12522 5212 12556 5245
rect 12522 5143 12556 5174
rect 12522 5140 12556 5143
rect 12522 5075 12556 5102
rect 12522 5068 12556 5075
rect 12522 5007 12556 5030
rect 12522 4996 12556 5007
rect 12522 4939 12556 4958
rect 12522 4924 12556 4939
rect 12522 4871 12556 4886
rect 12522 4852 12556 4871
rect 12522 4803 12556 4814
rect 12522 4780 12556 4803
rect 12522 4735 12556 4742
rect 12522 4708 12556 4735
rect 2330 4396 2334 4430
rect 2334 4396 2364 4430
rect 2402 4396 2436 4430
rect 2474 4397 2504 4431
rect 2504 4397 2508 4431
rect 2330 4323 2334 4357
rect 2334 4323 2364 4357
rect 2402 4323 2436 4357
rect 2474 4324 2504 4358
rect 2504 4324 2508 4358
rect 13948 5453 13956 5610
rect 13956 5453 14126 5610
rect 13948 5380 13956 5414
rect 13956 5380 13982 5414
rect 14020 5380 14054 5414
rect 14092 5380 14126 5414
rect 13948 5307 13956 5341
rect 13956 5307 13982 5341
rect 14020 5307 14054 5341
rect 14092 5307 14126 5341
rect 13948 5234 13956 5268
rect 13956 5234 13982 5268
rect 14020 5234 14054 5268
rect 14092 5234 14126 5268
rect 13948 5161 13956 5195
rect 13956 5161 13982 5195
rect 14020 5161 14054 5195
rect 14092 5161 14126 5195
rect 13948 5088 13956 5122
rect 13956 5088 13982 5122
rect 14020 5088 14054 5122
rect 14092 5088 14126 5122
rect 13948 5015 13956 5049
rect 13956 5015 13982 5049
rect 14020 5015 14054 5049
rect 14092 5015 14126 5049
rect 13948 4942 13956 4976
rect 13956 4942 13982 4976
rect 14020 4942 14054 4976
rect 14092 4942 14126 4976
rect 13948 4869 13956 4903
rect 13956 4869 13982 4903
rect 14020 4869 14054 4903
rect 14092 4869 14126 4903
rect 13948 4796 13956 4830
rect 13956 4796 13982 4830
rect 14020 4796 14054 4830
rect 14092 4796 14126 4830
rect 13948 4723 13956 4757
rect 13956 4723 13982 4757
rect 14020 4723 14054 4757
rect 14092 4723 14126 4757
rect 13948 4650 13956 4684
rect 13956 4650 13982 4684
rect 14020 4650 14054 4684
rect 14092 4650 14126 4684
rect 13948 4577 13956 4611
rect 13956 4577 13982 4611
rect 14020 4577 14054 4611
rect 14092 4577 14126 4611
rect 13948 4504 13956 4538
rect 13956 4504 13982 4538
rect 14020 4504 14054 4538
rect 14092 4504 14126 4538
rect 11597 4353 11629 4387
rect 11629 4353 11631 4387
rect 11669 4353 11697 4387
rect 11697 4353 11703 4387
rect 11741 4353 11765 4387
rect 11765 4353 11775 4387
rect 11813 4353 11833 4387
rect 11833 4353 11847 4387
rect 11885 4353 11901 4387
rect 11901 4353 11919 4387
rect 11957 4353 11969 4387
rect 11969 4353 11991 4387
rect 12029 4353 12037 4387
rect 12037 4353 12063 4387
rect 12101 4353 12105 4387
rect 12105 4353 12135 4387
rect 12173 4353 12207 4387
rect 12245 4353 12275 4387
rect 12275 4353 12279 4387
rect 12317 4353 12343 4387
rect 12343 4353 12351 4387
rect 2330 4250 2334 4284
rect 2334 4250 2364 4284
rect 2402 4250 2436 4284
rect 2474 4251 2504 4285
rect 2504 4251 2508 4285
rect 2330 4177 2334 4211
rect 2334 4177 2364 4211
rect 2402 4177 2436 4211
rect 2474 4178 2504 4212
rect 2504 4178 2508 4212
rect 2330 4104 2334 4138
rect 2334 4104 2364 4138
rect 2402 4104 2436 4138
rect 2474 4105 2504 4139
rect 2504 4105 2508 4139
rect 2330 4031 2334 4065
rect 2334 4031 2364 4065
rect 2402 4031 2436 4065
rect 2474 4032 2504 4066
rect 2504 4032 2508 4066
rect 2330 3958 2334 3992
rect 2334 3958 2364 3992
rect 2402 3958 2436 3992
rect 2474 3959 2504 3993
rect 2504 3959 2508 3993
rect 2330 3885 2334 3919
rect 2334 3885 2364 3919
rect 2402 3885 2436 3919
rect 2474 3886 2504 3920
rect 2504 3886 2508 3920
rect 2330 3812 2334 3846
rect 2334 3812 2364 3846
rect 2402 3812 2436 3846
rect 2474 3813 2504 3847
rect 2504 3813 2508 3847
rect 2330 3739 2334 3773
rect 2334 3739 2364 3773
rect 2402 3739 2436 3773
rect 2474 3740 2504 3774
rect 2504 3740 2508 3774
rect 2330 3666 2334 3700
rect 2334 3666 2364 3700
rect 2402 3666 2436 3700
rect 2474 3667 2504 3701
rect 2504 3667 2508 3701
rect 2330 3593 2334 3627
rect 2334 3593 2364 3627
rect 2402 3593 2436 3627
rect 2474 3594 2504 3628
rect 2504 3594 2508 3628
rect 2330 3520 2334 3554
rect 2334 3520 2364 3554
rect 2402 3520 2436 3554
rect 2474 3521 2504 3555
rect 2504 3521 2508 3555
rect 2330 3447 2334 3481
rect 2334 3447 2364 3481
rect 2402 3447 2436 3481
rect 2474 3448 2504 3482
rect 2504 3448 2508 3482
rect 2330 3374 2334 3408
rect 2334 3374 2364 3408
rect 2402 3374 2436 3408
rect 2474 3375 2504 3409
rect 2504 3375 2508 3409
rect 2330 3301 2334 3335
rect 2334 3301 2364 3335
rect 2402 3301 2436 3335
rect 2474 3302 2504 3336
rect 2504 3302 2508 3336
rect 2330 3228 2334 3262
rect 2334 3228 2364 3262
rect 2402 3228 2436 3262
rect 2474 3229 2504 3263
rect 2504 3229 2508 3263
rect 13953 4213 13956 4247
rect 13956 4213 13987 4247
rect 14091 4213 14125 4247
rect 13953 4138 13956 4172
rect 13956 4138 13987 4172
rect 14091 4138 14125 4172
rect 13953 4063 13956 4097
rect 13956 4063 13987 4097
rect 14091 4063 14125 4097
rect 13953 3988 13956 4022
rect 13956 3988 13987 4022
rect 14091 3988 14125 4022
rect 13953 3913 13956 3947
rect 13956 3913 13987 3947
rect 14091 3913 14125 3947
rect 13953 3838 13956 3872
rect 13956 3838 13987 3872
rect 14091 3838 14125 3872
rect 13953 3763 13956 3797
rect 13956 3763 13987 3797
rect 14091 3763 14125 3797
rect 13953 3688 13956 3722
rect 13956 3688 13987 3722
rect 14091 3688 14125 3722
rect 13953 3613 13956 3647
rect 13956 3613 13987 3647
rect 14091 3613 14125 3647
rect 13953 3537 13956 3571
rect 13956 3537 13987 3571
rect 14091 3537 14125 3571
rect 13953 3461 13956 3495
rect 13956 3461 13987 3495
rect 14091 3461 14125 3495
rect 13953 3385 13956 3419
rect 13956 3385 13987 3419
rect 14091 3385 14125 3419
rect 13953 3309 13956 3343
rect 13956 3309 13987 3343
rect 14091 3309 14125 3343
rect 13953 3233 13956 3267
rect 13956 3233 13987 3267
rect 14091 3233 14125 3267
rect 2330 3155 2334 3189
rect 2334 3155 2364 3189
rect 2402 3155 2436 3189
rect 2474 3156 2504 3190
rect 2504 3156 2508 3190
rect 2330 3082 2334 3116
rect 2334 3082 2364 3116
rect 2402 3082 2436 3116
rect 2474 3083 2504 3117
rect 2504 3083 2508 3117
rect 2330 3009 2334 3043
rect 2334 3009 2364 3043
rect 2402 3009 2436 3043
rect 2474 3010 2504 3044
rect 2504 3010 2508 3044
rect 2330 502 2334 2970
rect 2334 2898 2436 2970
rect 2474 2937 2504 2971
rect 2504 2937 2508 2971
rect 2334 502 2504 2898
rect 2504 502 2508 2898
rect 13953 2949 13956 2983
rect 13956 2949 13987 2983
rect 14091 2949 14125 2983
rect 13953 2874 13956 2908
rect 13956 2874 13987 2908
rect 14091 2874 14125 2908
rect 13953 2799 13956 2833
rect 13956 2799 13987 2833
rect 14091 2799 14125 2833
rect 13953 2724 13956 2758
rect 13956 2724 13987 2758
rect 14091 2724 14125 2758
rect 13953 2649 13956 2683
rect 13956 2649 13987 2683
rect 14091 2649 14125 2683
rect 13953 2574 13956 2608
rect 13956 2574 13987 2608
rect 14091 2574 14125 2608
rect 13953 2499 13956 2533
rect 13956 2499 13987 2533
rect 14091 2499 14125 2533
rect 13953 2424 13956 2458
rect 13956 2424 13987 2458
rect 14091 2424 14125 2458
rect 13953 2349 13956 2383
rect 13956 2349 13987 2383
rect 14091 2349 14125 2383
rect 13953 2273 13956 2307
rect 13956 2273 13987 2307
rect 14091 2273 14125 2307
rect 13953 2197 13956 2231
rect 13956 2197 13987 2231
rect 14091 2197 14125 2231
rect 13953 2121 13956 2155
rect 13956 2121 13987 2155
rect 14091 2121 14125 2155
rect 13953 2045 13956 2079
rect 13956 2045 13987 2079
rect 14091 2045 14125 2079
rect 13953 1969 13956 2003
rect 13956 1969 13987 2003
rect 14091 1969 14125 2003
rect 13953 1749 13956 1783
rect 13956 1749 13987 1783
rect 14091 1749 14125 1783
rect 13953 1674 13956 1708
rect 13956 1674 13987 1708
rect 14091 1674 14125 1708
rect 13953 1599 13956 1633
rect 13956 1599 13987 1633
rect 14091 1599 14125 1633
rect 13953 1524 13956 1558
rect 13956 1524 13987 1558
rect 14091 1524 14125 1558
rect 13953 1449 13956 1483
rect 13956 1449 13987 1483
rect 14091 1449 14125 1483
rect 13953 1374 13956 1408
rect 13956 1374 13987 1408
rect 14091 1374 14125 1408
rect 13953 1299 13956 1333
rect 13956 1299 13987 1333
rect 14091 1299 14125 1333
rect 13953 1224 13956 1258
rect 13956 1224 13987 1258
rect 14091 1224 14125 1258
rect 13953 1149 13956 1183
rect 13956 1149 13987 1183
rect 14091 1149 14125 1183
rect 13953 1073 13956 1107
rect 13956 1073 13987 1107
rect 14091 1073 14125 1107
rect 13953 997 13956 1031
rect 13956 997 13987 1031
rect 14091 997 14125 1031
rect 13953 921 13956 955
rect 13956 921 13987 955
rect 14091 921 14125 955
rect 13953 845 13956 879
rect 13956 845 13987 879
rect 14091 845 14125 879
rect 13953 769 13956 803
rect 13956 769 13987 803
rect 14091 769 14125 803
rect 2330 390 2508 502
rect 2330 356 2334 390
rect 2334 356 2368 390
rect 2368 356 2402 390
rect 2402 356 2436 390
rect 2436 374 2508 390
rect 13952 520 13956 554
rect 13956 520 13986 554
rect 14024 520 14058 554
rect 14096 520 14126 554
rect 14126 520 14130 554
rect 13952 432 13956 466
rect 13956 432 13986 466
rect 14024 438 14058 472
rect 14096 438 14126 472
rect 14126 438 14130 472
rect 2547 374 2581 378
rect 2620 374 2654 378
rect 2693 374 2727 378
rect 2766 374 2800 378
rect 2839 374 2873 378
rect 2912 374 2946 378
rect 2985 374 3019 378
rect 3058 374 3092 378
rect 3131 374 3165 378
rect 3204 374 3238 378
rect 3277 374 3311 378
rect 3350 374 3384 378
rect 3423 374 3457 378
rect 3496 374 3530 378
rect 3569 374 3603 378
rect 3642 374 3676 378
rect 3715 374 3749 378
rect 3788 374 3822 378
rect 3861 374 3895 378
rect 3934 374 3968 378
rect 4007 374 4041 378
rect 4080 374 4114 378
rect 4153 374 4187 378
rect 4226 374 4260 378
rect 4299 374 4333 378
rect 4372 374 4406 378
rect 4445 374 4479 378
rect 4518 374 4552 378
rect 4591 374 4625 378
rect 4664 374 13956 378
rect 2436 356 2470 374
rect 2330 344 2470 356
rect 2470 344 2508 374
rect 2547 344 2581 374
rect 2620 344 2654 374
rect 2693 344 2727 374
rect 2766 344 2800 374
rect 2839 344 2873 374
rect 2912 344 2946 374
rect 2985 344 3019 374
rect 3058 344 3092 374
rect 3131 344 3165 374
rect 3204 344 3238 374
rect 3277 344 3311 374
rect 3350 344 3384 374
rect 3423 344 3457 374
rect 3496 344 3530 374
rect 3569 344 3603 374
rect 3642 344 3676 374
rect 3715 344 3749 374
rect 3788 344 3822 374
rect 3861 344 3895 374
rect 3934 344 3968 374
rect 4007 344 4041 374
rect 4080 344 4114 374
rect 4153 344 4187 374
rect 4226 344 4260 374
rect 4299 344 4333 374
rect 4372 344 4406 374
rect 4445 344 4479 374
rect 4518 344 4552 374
rect 4591 344 4625 374
rect 2330 322 2436 344
rect 2330 288 2334 322
rect 2334 288 2368 322
rect 2368 306 2436 322
rect 4664 306 13860 374
rect 13860 340 13956 374
rect 13956 340 13986 378
rect 14024 355 14058 389
rect 14096 355 14126 389
rect 14126 355 14130 389
rect 13860 306 13986 340
rect 2368 288 2402 306
rect 2330 272 2402 288
rect 2402 272 2436 306
rect 2475 272 2509 306
rect 2548 272 2582 306
rect 2621 272 2655 306
rect 2694 272 2728 306
rect 2767 272 2801 306
rect 2840 272 2874 306
rect 2913 272 2947 306
rect 2986 272 3020 306
rect 3059 272 3093 306
rect 3132 272 3166 306
rect 3205 272 3239 306
rect 3278 272 3312 306
rect 3351 272 3385 306
rect 3424 272 3458 306
rect 3497 272 3531 306
rect 3570 272 3604 306
rect 3643 272 3677 306
rect 3716 272 3750 306
rect 3789 272 3823 306
rect 3862 272 3896 306
rect 3935 272 3969 306
rect 4008 272 4042 306
rect 4081 272 4115 306
rect 4154 272 4188 306
rect 4227 272 4261 306
rect 4300 272 4334 306
rect 4373 272 4407 306
rect 4446 272 4480 306
rect 4519 272 4553 306
rect 2402 204 2436 234
rect 2475 204 2509 234
rect 2548 204 2582 234
rect 2621 204 2655 234
rect 2694 204 2728 234
rect 2767 204 2801 234
rect 2840 204 2874 234
rect 2913 204 2947 234
rect 2986 204 3020 234
rect 3059 204 3093 234
rect 3132 204 3166 234
rect 3205 204 3239 234
rect 3278 204 3312 234
rect 3351 204 3385 234
rect 3424 204 3458 234
rect 3497 204 3531 234
rect 3570 204 3604 234
rect 3643 204 3677 234
rect 3716 204 3750 234
rect 3789 204 3823 234
rect 3862 204 3896 234
rect 3935 204 3969 234
rect 4008 204 4042 234
rect 4081 204 4115 234
rect 4154 204 4188 234
rect 4227 204 4261 234
rect 4300 204 4334 234
rect 4373 204 4407 234
rect 4446 204 4480 234
rect 4519 204 4553 234
rect 4592 204 13928 306
rect 13928 272 14024 306
rect 14024 272 14058 306
rect 14096 272 14126 306
rect 14126 272 14130 306
rect 13928 238 14058 272
rect 13928 204 13962 238
rect 13962 204 13996 238
rect 13996 204 14058 238
rect 2402 200 2436 204
rect 2475 200 2509 204
rect 2548 200 2582 204
rect 2621 200 2655 204
rect 2694 200 2728 204
rect 2767 200 2801 204
rect 2840 200 2874 204
rect 2913 200 2947 204
rect 2986 200 3020 204
rect 3059 200 3093 204
rect 3132 200 3166 204
rect 3205 200 3239 204
rect 3278 200 3312 204
rect 3351 200 3385 204
rect 3424 200 3458 204
rect 3497 200 3531 204
rect 3570 200 3604 204
rect 3643 200 3677 204
rect 3716 200 3750 204
rect 3789 200 3823 204
rect 3862 200 3896 204
rect 3935 200 3969 204
rect 4008 200 4042 204
rect 4081 200 4115 204
rect 4154 200 4188 204
rect 4227 200 4261 204
rect 4300 200 4334 204
rect 4373 200 4407 204
rect 4446 200 4480 204
rect 4519 200 4553 204
rect 4592 200 14058 204
<< metal1 >>
rect 1824 39939 14031 39945
rect 1824 39905 1902 39939
rect 1936 39905 1975 39939
rect 2009 39905 2048 39939
rect 2082 39905 2121 39939
rect 2155 39905 2194 39939
rect 2228 39905 2267 39939
rect 2301 39905 2340 39939
rect 2374 39905 2413 39939
rect 2447 39905 2486 39939
rect 2520 39905 2559 39939
rect 2593 39905 2632 39939
rect 2666 39905 2705 39939
rect 2739 39905 2778 39939
rect 2812 39905 2851 39939
rect 2885 39905 2924 39939
rect 2958 39905 2997 39939
rect 3031 39905 3070 39939
rect 3104 39905 3143 39939
rect 3177 39905 3216 39939
rect 3250 39905 3289 39939
rect 3323 39905 3362 39939
rect 3396 39905 3435 39939
rect 3469 39905 3508 39939
rect 3542 39905 3581 39939
rect 3615 39905 3654 39939
rect 3688 39905 3727 39939
rect 3761 39905 3800 39939
rect 3834 39905 3873 39939
rect 3907 39905 3946 39939
rect 3980 39905 4019 39939
rect 4053 39905 4092 39939
rect 4126 39905 4165 39939
rect 4199 39905 4238 39939
rect 4272 39905 4311 39939
rect 4345 39905 4384 39939
rect 4418 39905 4457 39939
rect 4491 39905 4530 39939
rect 4564 39905 4603 39939
rect 4637 39905 4676 39939
rect 4710 39905 4749 39939
rect 4783 39905 4822 39939
rect 4856 39905 4895 39939
rect 4929 39905 4968 39939
rect 5002 39905 5041 39939
rect 5075 39905 5114 39939
rect 5148 39905 5187 39939
rect 5221 39905 5260 39939
rect 5294 39905 5333 39939
rect 5367 39905 5406 39939
rect 5440 39905 5479 39939
rect 5513 39905 5552 39939
rect 5586 39905 5625 39939
rect 5659 39905 5698 39939
rect 5732 39905 5771 39939
rect 5805 39905 5844 39939
rect 5878 39905 5917 39939
rect 5951 39905 5990 39939
rect 6024 39905 6063 39939
rect 6097 39905 6136 39939
rect 6170 39905 6209 39939
rect 6243 39905 6282 39939
rect 6316 39905 6355 39939
rect 6389 39905 6428 39939
rect 6462 39905 6501 39939
rect 6535 39905 6574 39939
rect 6608 39905 6647 39939
rect 1824 39867 6647 39905
rect 1824 35873 1830 39867
rect 1936 39833 1975 39867
rect 2009 39833 2048 39867
rect 2082 39833 2121 39867
rect 2155 39833 2194 39867
rect 2228 39833 2267 39867
rect 2301 39833 2340 39867
rect 2374 39833 2413 39867
rect 2447 39833 2486 39867
rect 2520 39833 2559 39867
rect 2593 39833 2632 39867
rect 2666 39833 2705 39867
rect 2739 39833 2778 39867
rect 2812 39833 2851 39867
rect 2885 39833 2924 39867
rect 2958 39833 2997 39867
rect 3031 39833 3070 39867
rect 3104 39833 3143 39867
rect 3177 39833 3216 39867
rect 3250 39833 3289 39867
rect 3323 39833 3362 39867
rect 3396 39833 3435 39867
rect 3469 39833 3508 39867
rect 3542 39833 3581 39867
rect 3615 39833 3654 39867
rect 3688 39833 3727 39867
rect 3761 39833 3800 39867
rect 3834 39833 3873 39867
rect 3907 39833 3946 39867
rect 3980 39833 4019 39867
rect 4053 39833 4092 39867
rect 4126 39833 4165 39867
rect 4199 39833 4238 39867
rect 4272 39833 4311 39867
rect 4345 39833 4384 39867
rect 4418 39833 4457 39867
rect 4491 39833 4530 39867
rect 4564 39833 4603 39867
rect 4637 39833 4676 39867
rect 4710 39833 4749 39867
rect 4783 39833 4822 39867
rect 4856 39833 4895 39867
rect 4929 39833 4968 39867
rect 5002 39833 5041 39867
rect 5075 39833 5114 39867
rect 5148 39833 5187 39867
rect 5221 39833 5260 39867
rect 5294 39833 5333 39867
rect 5367 39833 5406 39867
rect 5440 39833 5479 39867
rect 5513 39833 5552 39867
rect 5586 39833 5625 39867
rect 5659 39833 5698 39867
rect 5732 39833 5771 39867
rect 5805 39833 5844 39867
rect 5878 39833 5917 39867
rect 5951 39833 5990 39867
rect 6024 39833 6063 39867
rect 6097 39833 6136 39867
rect 6170 39833 6209 39867
rect 6243 39833 6282 39867
rect 6316 39833 6355 39867
rect 6389 39833 6428 39867
rect 6462 39833 6501 39867
rect 6535 39833 6574 39867
rect 6608 39833 6647 39867
rect 13953 39867 14031 39939
rect 13953 39833 13991 39867
rect 14025 39833 14031 39867
rect 14437 39876 14567 39882
rect 14437 39842 14449 39876
rect 14483 39842 14521 39876
rect 14555 39842 14567 39876
rect 14437 39836 14567 39842
rect 1936 39795 6719 39833
rect 2008 39761 2047 39795
rect 2081 39761 2120 39795
rect 2154 39761 2193 39795
rect 2227 39761 2266 39795
rect 2300 39761 2339 39795
rect 2373 39761 2412 39795
rect 2446 39761 2485 39795
rect 2519 39761 2558 39795
rect 2592 39761 2631 39795
rect 2665 39761 2704 39795
rect 2738 39761 2777 39795
rect 2811 39761 2850 39795
rect 2884 39761 2923 39795
rect 2957 39761 2996 39795
rect 3030 39761 3069 39795
rect 3103 39761 3142 39795
rect 3176 39761 3215 39795
rect 3249 39761 3288 39795
rect 3322 39761 3361 39795
rect 3395 39761 3434 39795
rect 3468 39761 3507 39795
rect 3541 39761 3580 39795
rect 3614 39761 3653 39795
rect 3687 39761 3726 39795
rect 3760 39761 3799 39795
rect 3833 39761 3872 39795
rect 3906 39761 3945 39795
rect 3979 39761 4018 39795
rect 4052 39761 4091 39795
rect 4125 39761 4164 39795
rect 4198 39761 4237 39795
rect 4271 39761 4310 39795
rect 4344 39761 4383 39795
rect 4417 39761 4456 39795
rect 4490 39761 4529 39795
rect 4563 39761 4602 39795
rect 4636 39761 4675 39795
rect 4709 39761 4748 39795
rect 4782 39761 4821 39795
rect 4855 39761 4894 39795
rect 4928 39761 4967 39795
rect 5001 39761 5040 39795
rect 5074 39761 5113 39795
rect 5147 39761 5186 39795
rect 5220 39761 5259 39795
rect 5293 39761 5332 39795
rect 5366 39761 5405 39795
rect 5439 39761 5478 39795
rect 5512 39761 5551 39795
rect 5585 39761 5624 39795
rect 5658 39761 5697 39795
rect 5731 39761 5770 39795
rect 5804 39761 5843 39795
rect 5877 39761 5916 39795
rect 5950 39761 5989 39795
rect 6023 39761 6062 39795
rect 6096 39761 6135 39795
rect 6169 39761 6208 39795
rect 6242 39761 6281 39795
rect 6315 39761 6354 39795
rect 6388 39761 6427 39795
rect 6461 39761 6500 39795
rect 6534 39761 6573 39795
rect 6607 39761 6646 39795
rect 6680 39761 6719 39795
rect 13881 39794 14031 39833
tri 14442 39802 14476 39836 ne
rect 13881 39761 13919 39794
rect 2008 39723 6791 39761
rect 2080 39689 2119 39723
rect 2153 39689 2192 39723
rect 2226 39689 2265 39723
rect 2299 39689 2338 39723
rect 2372 39689 2411 39723
rect 2445 39689 2484 39723
rect 2518 39689 2557 39723
rect 2591 39689 2630 39723
rect 2664 39689 2703 39723
rect 2737 39689 2776 39723
rect 2810 39689 2849 39723
rect 2883 39689 2922 39723
rect 2956 39689 2995 39723
rect 3029 39689 3068 39723
rect 3102 39689 3141 39723
rect 3175 39689 3214 39723
rect 3248 39689 3287 39723
rect 3321 39689 3360 39723
rect 3394 39689 3433 39723
rect 3467 39689 3506 39723
rect 3540 39689 3579 39723
rect 3613 39689 3652 39723
rect 3686 39689 3725 39723
rect 3759 39689 3798 39723
rect 3832 39689 3871 39723
rect 3905 39689 3944 39723
rect 3978 39689 4017 39723
rect 4051 39689 4090 39723
rect 4124 39689 4163 39723
rect 4197 39689 4236 39723
rect 4270 39689 4309 39723
rect 4343 39689 4382 39723
rect 4416 39689 4455 39723
rect 4489 39689 4528 39723
rect 4562 39689 4601 39723
rect 4635 39689 4674 39723
rect 4708 39689 4747 39723
rect 4781 39689 4820 39723
rect 4854 39689 4893 39723
rect 4927 39689 4966 39723
rect 5000 39689 5039 39723
rect 5073 39689 5112 39723
rect 5146 39689 5185 39723
rect 5219 39689 5258 39723
rect 5292 39689 5331 39723
rect 5365 39689 5404 39723
rect 5438 39689 5477 39723
rect 5511 39689 5550 39723
rect 5584 39689 5623 39723
rect 5657 39689 5696 39723
rect 5730 39689 5769 39723
rect 5803 39689 5842 39723
rect 5876 39689 5915 39723
rect 5949 39689 5988 39723
rect 6022 39689 6061 39723
rect 6095 39689 6134 39723
rect 6168 39689 6207 39723
rect 6241 39689 6280 39723
rect 6314 39689 6353 39723
rect 6387 39689 6426 39723
rect 6460 39689 6499 39723
rect 6533 39689 6572 39723
rect 6606 39689 6645 39723
rect 6679 39689 6718 39723
rect 6752 39689 6791 39723
rect 13809 39760 13919 39761
rect 13953 39760 13991 39794
rect 14025 39760 14031 39794
rect 13809 39722 14031 39760
rect 13809 39689 13847 39722
rect 2080 39688 13847 39689
rect 13881 39721 14031 39722
rect 13881 39688 13919 39721
rect 2080 39687 13919 39688
rect 13953 39687 13991 39721
rect 14025 39687 14031 39721
rect 2080 39683 14031 39687
rect 2080 39650 2197 39683
tri 2197 39650 2230 39683 nw
tri 13601 39650 13634 39683 ne
rect 13634 39650 14031 39683
rect 2080 39616 2163 39650
tri 2163 39616 2197 39650 nw
tri 13634 39616 13668 39650 ne
rect 13668 39616 13775 39650
rect 13809 39649 14031 39650
rect 13809 39616 13847 39649
rect 2080 39615 2162 39616
tri 2162 39615 2163 39616 nw
tri 13668 39615 13669 39616 ne
rect 13669 39615 13847 39616
rect 13881 39648 14031 39649
rect 13881 39615 13919 39648
rect 2080 39614 2161 39615
tri 2161 39614 2162 39615 nw
tri 13669 39614 13670 39615 ne
rect 13670 39614 13919 39615
rect 13953 39614 13991 39648
rect 14025 39614 14031 39648
rect 2080 39577 2124 39614
tri 2124 39577 2161 39614 nw
tri 13670 39577 13707 39614 ne
rect 13707 39577 14031 39614
rect 2080 39551 2098 39577
tri 2098 39551 2124 39577 nw
tri 13707 39551 13733 39577 ne
rect 13733 39551 13775 39577
rect 2080 39545 2092 39551
tri 2092 39545 2098 39551 nw
rect 2214 39545 13637 39551
rect 2080 35873 2086 39545
tri 2086 39539 2092 39545 nw
rect 1824 35834 2086 35873
rect 1824 35800 1830 35834
rect 1864 35800 1902 35834
rect 1936 35800 1974 35834
rect 2008 35800 2046 35834
rect 2080 35800 2086 35834
rect 1824 35761 2086 35800
rect 1824 35727 1830 35761
rect 1864 35727 1902 35761
rect 1936 35727 1974 35761
rect 2008 35727 2046 35761
rect 2080 35727 2086 35761
rect 1824 35688 2086 35727
rect 1824 35654 1830 35688
rect 1864 35654 1902 35688
rect 1936 35654 1974 35688
rect 2008 35654 2046 35688
rect 2080 35654 2086 35688
rect 1824 35615 2086 35654
rect 1824 35581 1830 35615
rect 1864 35581 1902 35615
rect 1936 35581 1974 35615
rect 2008 35581 2046 35615
rect 2080 35581 2086 35615
rect 1824 35542 2086 35581
rect 1824 35508 1830 35542
rect 1864 35508 1902 35542
rect 1936 35508 1974 35542
rect 2008 35508 2046 35542
rect 2080 35508 2086 35542
rect 1824 35469 2086 35508
rect 1824 35435 1830 35469
rect 1864 35435 1902 35469
rect 1936 35435 1974 35469
rect 2008 35435 2046 35469
rect 2080 35435 2086 35469
rect 1824 35396 2086 35435
rect 1824 35362 1830 35396
rect 1864 35362 1902 35396
rect 1936 35362 1974 35396
rect 2008 35362 2046 35396
rect 2080 35362 2086 35396
rect 1824 35323 2086 35362
rect 1824 35289 1830 35323
rect 1864 35289 1902 35323
rect 1936 35289 1974 35323
rect 2008 35289 2046 35323
rect 2080 35289 2086 35323
rect 1824 35250 2086 35289
rect 1824 35216 1830 35250
rect 1864 35216 1902 35250
rect 1936 35216 1974 35250
rect 2008 35216 2046 35250
rect 2080 35216 2086 35250
rect 1824 35177 2086 35216
rect 1824 35143 1830 35177
rect 1864 35143 1902 35177
rect 1936 35143 1974 35177
rect 2008 35143 2046 35177
rect 2080 35143 2086 35177
rect 1824 35104 2086 35143
rect 1824 35070 1830 35104
rect 1864 35070 1902 35104
rect 1936 35070 1974 35104
rect 2008 35070 2046 35104
rect 2080 35070 2086 35104
rect 1824 35031 2086 35070
rect 1824 34997 1830 35031
rect 1864 34997 1902 35031
rect 1936 34997 1974 35031
rect 2008 34997 2046 35031
rect 2080 34997 2086 35031
rect 1824 34958 2086 34997
rect 1824 34924 1830 34958
rect 1864 34924 1902 34958
rect 1936 34924 1974 34958
rect 2008 34924 2046 34958
rect 2080 34924 2086 34958
rect 1824 34885 2086 34924
rect 1824 34851 1830 34885
rect 1864 34851 1902 34885
rect 1936 34851 1974 34885
rect 2008 34851 2046 34885
rect 2080 34851 2086 34885
rect 1824 34812 2086 34851
rect 1824 34778 1830 34812
rect 1864 34778 1902 34812
rect 1936 34778 1974 34812
rect 2008 34778 2046 34812
rect 2080 34778 2086 34812
rect 1824 34739 2086 34778
rect 1824 34705 1830 34739
rect 1864 34705 1902 34739
rect 1936 34705 1974 34739
rect 2008 34705 2046 34739
rect 2080 34705 2086 34739
rect 1824 34666 2086 34705
rect 1824 34632 1830 34666
rect 1864 34632 1902 34666
rect 1936 34632 1974 34666
rect 2008 34632 2046 34666
rect 2080 34632 2086 34666
rect 1824 34593 2086 34632
rect 1824 34559 1830 34593
rect 1864 34559 1902 34593
rect 1936 34559 1974 34593
rect 2008 34559 2046 34593
rect 2080 34559 2086 34593
rect 1824 34520 2086 34559
rect 1824 34486 1830 34520
rect 1864 34486 1902 34520
rect 1936 34486 1974 34520
rect 2008 34486 2046 34520
rect 2080 34486 2086 34520
rect 1824 34447 2086 34486
rect 1824 34413 1830 34447
rect 1864 34413 1902 34447
rect 1936 34413 1974 34447
rect 2008 34413 2046 34447
rect 2080 34413 2086 34447
rect 1824 34374 2086 34413
rect 1824 34340 1830 34374
rect 1864 34340 1902 34374
rect 1936 34340 1974 34374
rect 2008 34340 2046 34374
rect 2080 34340 2086 34374
rect 1824 34301 2086 34340
tri 1792 34267 1824 34299 se
rect 1824 34267 1830 34301
rect 1864 34267 1902 34301
rect 1936 34267 1974 34301
rect 2008 34267 2046 34301
rect 2080 34267 2086 34301
tri 1765 34240 1792 34267 se
rect 1792 34240 2086 34267
tri 1764 34239 1765 34240 se
rect 1765 34239 2086 34240
tri 1753 34228 1764 34239 se
rect 1764 34228 2086 34239
tri 1719 34194 1753 34228 se
rect 1753 34194 1830 34228
rect 1864 34194 1902 34228
rect 1936 34194 1974 34228
rect 2008 34194 2046 34228
rect 2080 34194 2086 34228
tri 1707 34182 1719 34194 se
rect 1719 34182 2086 34194
rect 2214 39511 2292 39545
rect 2326 39511 2365 39545
rect 2214 39473 2365 39511
rect 2214 37855 2220 39473
rect 2326 39439 2365 39473
rect 13559 39473 13637 39545
tri 13733 39543 13741 39551 ne
rect 13741 39543 13775 39551
rect 13809 39576 14031 39577
rect 13809 39543 13847 39576
tri 13741 39542 13742 39543 ne
rect 13742 39542 13847 39543
rect 13881 39575 14031 39576
rect 13881 39542 13919 39575
tri 13742 39541 13743 39542 ne
rect 13743 39541 13919 39542
rect 13953 39541 13991 39575
rect 14025 39541 14031 39575
tri 13743 39515 13769 39541 ne
rect 13559 39439 13597 39473
rect 13631 39439 13637 39473
rect 2326 39401 2437 39439
rect 2398 39367 2437 39401
rect 13487 39400 13637 39439
rect 13487 39367 13525 39400
rect 2398 39366 13525 39367
rect 13559 39366 13597 39400
rect 13631 39366 13637 39400
rect 2398 39361 13637 39366
rect 2398 39358 2467 39361
tri 2467 39358 2470 39361 nw
tri 13381 39358 13384 39361 ne
rect 13384 39358 13637 39361
rect 2398 39328 2437 39358
tri 2437 39328 2467 39358 nw
tri 13384 39328 13414 39358 ne
rect 13414 39328 13637 39358
rect 2398 37855 2404 39328
tri 2404 39295 2437 39328 nw
tri 13414 39295 13447 39328 ne
rect 13447 39294 13453 39328
rect 13487 39327 13637 39328
rect 13487 39294 13525 39327
rect 13447 39293 13525 39294
rect 13559 39293 13597 39327
rect 13631 39293 13637 39327
rect 13447 39255 13637 39293
rect 13447 39221 13453 39255
rect 13487 39254 13637 39255
rect 13487 39221 13525 39254
rect 13447 39220 13525 39221
rect 13559 39220 13597 39254
rect 13631 39220 13637 39254
rect 13447 39182 13637 39220
rect 13447 39148 13453 39182
rect 13487 39181 13637 39182
rect 13487 39148 13525 39181
rect 13447 39147 13525 39148
rect 13559 39147 13597 39181
rect 13631 39147 13637 39181
rect 2214 37816 2231 37855
rect 2283 37816 2335 37855
rect 2387 37816 2404 37855
rect 2214 37782 2220 37816
rect 2283 37813 2292 37816
rect 2254 37801 2292 37813
rect 2283 37782 2292 37801
rect 2326 37813 2335 37816
rect 2326 37801 2364 37813
rect 2326 37782 2335 37801
rect 2398 37782 2404 37816
rect 2214 37749 2231 37782
rect 2283 37749 2335 37782
rect 2387 37749 2404 37782
rect 2214 37743 2404 37749
rect 2214 37709 2220 37743
rect 2254 37737 2292 37743
rect 2283 37709 2292 37737
rect 2326 37737 2364 37743
rect 2326 37709 2335 37737
rect 2398 37709 2404 37743
rect 2214 37685 2231 37709
rect 2283 37685 2335 37709
rect 2387 37685 2404 37709
rect 2214 37673 2404 37685
rect 2214 37670 2231 37673
rect 2283 37670 2335 37673
rect 2387 37670 2404 37673
rect 2214 37636 2220 37670
rect 2283 37636 2292 37670
rect 2326 37636 2335 37670
rect 2398 37636 2404 37670
rect 2214 37621 2231 37636
rect 2283 37621 2335 37636
rect 2387 37621 2404 37636
rect 2214 37609 2404 37621
rect 2214 37597 2231 37609
rect 2283 37597 2335 37609
rect 2387 37597 2404 37609
rect 2214 37563 2220 37597
rect 2283 37563 2292 37597
rect 2326 37563 2335 37597
rect 2398 37563 2404 37597
rect 2214 37557 2231 37563
rect 2283 37557 2335 37563
rect 2387 37557 2404 37563
rect 2214 37545 2404 37557
rect 2214 37524 2231 37545
rect 2283 37524 2335 37545
rect 2387 37524 2404 37545
rect 2214 37490 2220 37524
rect 2283 37493 2292 37524
rect 2254 37490 2292 37493
rect 2326 37493 2335 37524
rect 2326 37490 2364 37493
rect 2398 37490 2404 37524
rect 2214 37481 2404 37490
rect 2214 37451 2231 37481
rect 2283 37451 2335 37481
rect 2387 37451 2404 37481
rect 2214 37417 2220 37451
rect 2283 37429 2292 37451
rect 2254 37417 2292 37429
rect 2326 37429 2335 37451
rect 2326 37417 2364 37429
rect 2398 37417 2404 37451
rect 2214 37378 2231 37417
rect 2283 37378 2335 37417
rect 2387 37378 2404 37417
rect 2214 37344 2220 37378
rect 2283 37365 2292 37378
rect 2254 37353 2292 37365
rect 2283 37344 2292 37353
rect 2326 37365 2335 37378
rect 2326 37353 2364 37365
rect 2326 37344 2335 37353
rect 2398 37344 2404 37378
rect 2214 37305 2231 37344
rect 2283 37305 2335 37344
rect 2387 37305 2404 37344
rect 2214 37271 2220 37305
rect 2283 37301 2292 37305
rect 2254 37289 2292 37301
rect 2283 37271 2292 37289
rect 2326 37301 2335 37305
rect 2326 37289 2364 37301
rect 2326 37271 2335 37289
rect 2398 37271 2404 37305
rect 2214 37237 2231 37271
rect 2283 37237 2335 37271
rect 2387 37237 2404 37271
rect 2214 37232 2404 37237
rect 2214 37198 2220 37232
rect 2254 37225 2292 37232
rect 2283 37198 2292 37225
rect 2326 37225 2364 37232
rect 2326 37198 2335 37225
rect 2398 37198 2404 37232
rect 2214 37173 2231 37198
rect 2283 37173 2335 37198
rect 2387 37173 2404 37198
rect 2214 37161 2404 37173
rect 2214 37159 2231 37161
rect 2283 37159 2335 37161
rect 2387 37159 2404 37161
rect 2214 37125 2220 37159
rect 2283 37125 2292 37159
rect 2326 37125 2335 37159
rect 2398 37125 2404 37159
rect 2214 37109 2231 37125
rect 2283 37109 2335 37125
rect 2387 37109 2404 37125
rect 2214 37097 2404 37109
rect 2214 37086 2231 37097
rect 2283 37086 2335 37097
rect 2387 37086 2404 37097
rect 2214 37052 2220 37086
rect 2283 37052 2292 37086
rect 2326 37052 2335 37086
rect 2398 37052 2404 37086
rect 2214 37045 2231 37052
rect 2283 37045 2335 37052
rect 2387 37045 2404 37052
rect 2214 37033 2404 37045
rect 2214 37013 2231 37033
rect 2283 37013 2335 37033
rect 2387 37013 2404 37033
rect 2214 36979 2220 37013
rect 2283 36981 2292 37013
rect 2254 36979 2292 36981
rect 2326 36981 2335 37013
rect 2326 36979 2364 36981
rect 2398 36979 2404 37013
rect 2214 36969 2404 36979
rect 2214 36940 2231 36969
rect 2283 36940 2335 36969
rect 2387 36940 2404 36969
rect 2214 36906 2220 36940
rect 2283 36917 2292 36940
rect 2254 36906 2292 36917
rect 2326 36917 2335 36940
rect 2326 36906 2364 36917
rect 2398 36906 2404 36940
rect 2214 36905 2404 36906
rect 2214 36867 2231 36905
rect 2283 36867 2335 36905
rect 2387 36867 2404 36905
rect 2214 36833 2220 36867
rect 2283 36853 2292 36867
rect 2254 36841 2292 36853
rect 2283 36833 2292 36841
rect 2326 36853 2335 36867
rect 2326 36841 2364 36853
rect 2326 36833 2335 36841
rect 2398 36833 2404 36867
rect 2214 36794 2231 36833
rect 2283 36794 2335 36833
rect 2387 36794 2404 36833
rect 2214 36760 2220 36794
rect 2283 36789 2292 36794
rect 2254 36777 2292 36789
rect 2283 36760 2292 36777
rect 2326 36789 2335 36794
rect 2326 36777 2364 36789
rect 2326 36760 2335 36777
rect 2398 36760 2404 36794
rect 2214 36725 2231 36760
rect 2283 36725 2335 36760
rect 2387 36725 2404 36760
rect 2214 36721 2404 36725
rect 2214 36687 2220 36721
rect 2254 36713 2292 36721
rect 2283 36687 2292 36713
rect 2326 36713 2364 36721
rect 2326 36687 2335 36713
rect 2398 36687 2404 36721
rect 2214 36661 2231 36687
rect 2283 36661 2335 36687
rect 2387 36661 2404 36687
rect 2214 36649 2404 36661
rect 2214 36648 2231 36649
rect 2283 36648 2335 36649
rect 2387 36648 2404 36649
rect 2214 36614 2220 36648
rect 2283 36614 2292 36648
rect 2326 36614 2335 36648
rect 2398 36614 2404 36648
rect 2214 36597 2231 36614
rect 2283 36597 2335 36614
rect 2387 36597 2404 36614
rect 2214 36585 2404 36597
rect 2214 36575 2231 36585
rect 2283 36575 2335 36585
rect 2387 36575 2404 36585
rect 2214 36541 2220 36575
rect 2283 36541 2292 36575
rect 2326 36541 2335 36575
rect 2398 36541 2404 36575
rect 2214 36533 2231 36541
rect 2283 36533 2335 36541
rect 2387 36533 2404 36541
rect 2214 36521 2404 36533
rect 2214 36502 2231 36521
rect 2283 36502 2335 36521
rect 2387 36502 2404 36521
rect 2214 36468 2220 36502
rect 2283 36469 2292 36502
rect 2254 36468 2292 36469
rect 2326 36469 2335 36502
rect 2326 36468 2364 36469
rect 2398 36468 2404 36502
rect 2214 36457 2404 36468
rect 2214 36429 2231 36457
rect 2283 36429 2335 36457
rect 2387 36429 2404 36457
rect 2214 36395 2220 36429
rect 2283 36405 2292 36429
rect 2254 36395 2292 36405
rect 2326 36405 2335 36429
rect 2326 36395 2364 36405
rect 2398 36395 2404 36429
rect 2214 36393 2404 36395
rect 2214 36356 2231 36393
rect 2283 36356 2335 36393
rect 2387 36356 2404 36393
rect 2214 36322 2220 36356
rect 2283 36341 2292 36356
rect 2254 36329 2292 36341
rect 2283 36322 2292 36329
rect 2326 36341 2335 36356
rect 2326 36329 2364 36341
rect 2326 36322 2335 36329
rect 2398 36322 2404 36356
rect 2214 36283 2231 36322
rect 2283 36283 2335 36322
rect 2387 36283 2404 36322
rect 2214 36249 2220 36283
rect 2283 36277 2292 36283
rect 2254 36265 2292 36277
rect 2283 36249 2292 36265
rect 2326 36277 2335 36283
rect 2326 36265 2364 36277
rect 2326 36249 2335 36265
rect 2398 36249 2404 36283
rect 2214 36213 2231 36249
rect 2283 36213 2335 36249
rect 2387 36213 2404 36249
rect 2214 36210 2404 36213
rect 2214 36176 2220 36210
rect 2254 36201 2292 36210
rect 2283 36176 2292 36201
rect 2326 36201 2364 36210
rect 2326 36176 2335 36201
rect 2398 36176 2404 36210
rect 2214 36149 2231 36176
rect 2283 36149 2335 36176
rect 2387 36149 2404 36176
rect 2214 36137 2404 36149
rect 2214 36103 2220 36137
rect 2283 36103 2292 36137
rect 2326 36103 2335 36137
rect 2398 36103 2404 36137
rect 2214 36085 2231 36103
rect 2283 36085 2335 36103
rect 2387 36085 2404 36103
rect 2214 36073 2404 36085
rect 2214 36064 2231 36073
rect 2283 36064 2335 36073
rect 2387 36064 2404 36073
rect 2214 36030 2220 36064
rect 2283 36030 2292 36064
rect 2326 36030 2335 36064
rect 2398 36030 2404 36064
rect 2214 36021 2231 36030
rect 2283 36021 2335 36030
rect 2387 36021 2404 36030
rect 2214 36009 2404 36021
rect 2214 35991 2231 36009
rect 2283 35991 2335 36009
rect 2387 35991 2404 36009
rect 2214 35957 2220 35991
rect 2283 35957 2292 35991
rect 2326 35957 2335 35991
rect 2398 35957 2404 35991
rect 2214 35945 2404 35957
rect 2214 35918 2231 35945
rect 2283 35918 2335 35945
rect 2387 35918 2404 35945
rect 2214 35884 2220 35918
rect 2283 35893 2292 35918
rect 2254 35884 2292 35893
rect 2326 35893 2335 35918
rect 2326 35884 2364 35893
rect 2398 35884 2404 35918
rect 2214 35881 2404 35884
rect 2214 35845 2231 35881
rect 2283 35845 2335 35881
rect 2387 35845 2404 35881
rect 2214 35811 2220 35845
rect 2283 35829 2292 35845
rect 2254 35817 2292 35829
rect 2283 35811 2292 35817
rect 2326 35829 2335 35845
rect 2326 35817 2364 35829
rect 2326 35811 2335 35817
rect 2398 35811 2404 35845
rect 2214 35772 2231 35811
rect 2283 35772 2335 35811
rect 2387 35772 2404 35811
rect 2214 35738 2220 35772
rect 2283 35765 2292 35772
rect 2254 35753 2292 35765
rect 2283 35738 2292 35753
rect 2326 35765 2335 35772
rect 2326 35753 2364 35765
rect 2326 35738 2335 35753
rect 2398 35738 2404 35772
rect 2214 35701 2231 35738
rect 2283 35701 2335 35738
rect 2387 35701 2404 35738
rect 2214 35699 2404 35701
rect 2214 35665 2220 35699
rect 2254 35689 2292 35699
rect 2283 35665 2292 35689
rect 2326 35689 2364 35699
rect 2326 35665 2335 35689
rect 2398 35665 2404 35699
rect 2214 35637 2231 35665
rect 2283 35637 2335 35665
rect 2387 35637 2404 35665
rect 2214 35626 2404 35637
rect 2214 35592 2220 35626
rect 2254 35625 2292 35626
rect 2283 35592 2292 35625
rect 2326 35625 2364 35626
rect 2326 35592 2335 35625
rect 2398 35592 2404 35626
rect 2214 35573 2231 35592
rect 2283 35573 2335 35592
rect 2387 35573 2404 35592
rect 2214 35561 2404 35573
rect 2214 35553 2231 35561
rect 2283 35553 2335 35561
rect 2387 35553 2404 35561
rect 2214 35519 2220 35553
rect 2283 35519 2292 35553
rect 2326 35519 2335 35553
rect 2398 35519 2404 35553
rect 2214 35509 2231 35519
rect 2283 35509 2335 35519
rect 2387 35509 2404 35519
rect 2214 35497 2404 35509
rect 2214 35480 2231 35497
rect 2283 35480 2335 35497
rect 2387 35480 2404 35497
rect 2214 35446 2220 35480
rect 2283 35446 2292 35480
rect 2326 35446 2335 35480
rect 2398 35446 2404 35480
rect 2214 35445 2231 35446
rect 2283 35445 2335 35446
rect 2387 35445 2404 35446
rect 2214 35433 2404 35445
rect 2214 35407 2231 35433
rect 2283 35407 2335 35433
rect 2387 35407 2404 35433
rect 2214 35373 2220 35407
rect 2283 35381 2292 35407
rect 2254 35373 2292 35381
rect 2326 35381 2335 35407
rect 2326 35373 2364 35381
rect 2398 35373 2404 35407
rect 2214 35369 2404 35373
rect 2214 35334 2231 35369
rect 2283 35334 2335 35369
rect 2387 35334 2404 35369
rect 2214 35300 2220 35334
rect 2283 35317 2292 35334
rect 2254 35305 2292 35317
rect 2283 35300 2292 35305
rect 2326 35317 2335 35334
rect 2326 35305 2364 35317
rect 2326 35300 2335 35305
rect 2398 35300 2404 35334
rect 2214 35261 2231 35300
rect 2283 35261 2335 35300
rect 2387 35261 2404 35300
rect 2214 35227 2220 35261
rect 2283 35253 2292 35261
rect 2254 35241 2292 35253
rect 2283 35227 2292 35241
rect 2326 35253 2335 35261
rect 2326 35241 2364 35253
rect 2326 35227 2335 35241
rect 2398 35227 2404 35261
rect 2214 35189 2231 35227
rect 2283 35189 2335 35227
rect 2387 35189 2404 35227
rect 2214 35188 2404 35189
rect 2214 35154 2220 35188
rect 2254 35176 2292 35188
rect 2283 35154 2292 35176
rect 2326 35176 2364 35188
rect 2326 35154 2335 35176
rect 2398 35154 2404 35188
rect 2214 35124 2231 35154
rect 2283 35124 2335 35154
rect 2387 35124 2404 35154
rect 2214 35115 2404 35124
rect 2214 35081 2220 35115
rect 2254 35111 2292 35115
rect 2283 35081 2292 35111
rect 2326 35111 2364 35115
rect 2326 35081 2335 35111
rect 2398 35081 2404 35115
rect 2214 35059 2231 35081
rect 2283 35059 2335 35081
rect 2387 35059 2404 35081
rect 2214 35046 2404 35059
rect 2214 35042 2231 35046
rect 2283 35042 2335 35046
rect 2387 35042 2404 35046
rect 2214 35008 2220 35042
rect 2283 35008 2292 35042
rect 2326 35008 2335 35042
rect 2398 35008 2404 35042
rect 2214 34994 2231 35008
rect 2283 34994 2335 35008
rect 2387 34994 2404 35008
rect 2214 34981 2404 34994
rect 2214 34969 2231 34981
rect 2283 34969 2335 34981
rect 2387 34969 2404 34981
rect 2214 34935 2220 34969
rect 2283 34935 2292 34969
rect 2326 34935 2335 34969
rect 2398 34935 2404 34969
rect 2214 34929 2231 34935
rect 2283 34929 2335 34935
rect 2387 34929 2404 34935
rect 2214 34916 2404 34929
rect 2214 34896 2231 34916
rect 2283 34896 2335 34916
rect 2387 34896 2404 34916
rect 2214 34862 2220 34896
rect 2283 34864 2292 34896
rect 2254 34862 2292 34864
rect 2326 34864 2335 34896
rect 2326 34862 2364 34864
rect 2398 34862 2404 34896
rect 2214 34851 2404 34862
rect 2214 34823 2231 34851
rect 2283 34823 2335 34851
rect 2387 34823 2404 34851
rect 2214 34789 2220 34823
rect 2283 34799 2292 34823
rect 2254 34789 2292 34799
rect 2326 34799 2335 34823
rect 2326 34789 2364 34799
rect 2398 34789 2404 34823
rect 2214 34786 2404 34789
rect 2214 34750 2231 34786
rect 2283 34750 2335 34786
rect 2387 34750 2404 34786
rect 2214 34716 2220 34750
rect 2283 34734 2292 34750
rect 2254 34721 2292 34734
rect 2283 34716 2292 34721
rect 2326 34734 2335 34750
rect 2326 34721 2364 34734
rect 2326 34716 2335 34721
rect 2398 34716 2404 34750
rect 2214 34677 2231 34716
rect 2283 34677 2335 34716
rect 2387 34677 2404 34716
rect 2214 34643 2220 34677
rect 2283 34669 2292 34677
rect 2254 34656 2292 34669
rect 2283 34643 2292 34656
rect 2326 34669 2335 34677
rect 2326 34656 2364 34669
rect 2326 34643 2335 34656
rect 2398 34643 2404 34677
rect 2214 34604 2231 34643
rect 2283 34604 2335 34643
rect 2387 34604 2404 34643
rect 2214 34570 2220 34604
rect 2254 34591 2292 34604
rect 2283 34570 2292 34591
rect 2326 34591 2364 34604
rect 2326 34570 2335 34591
rect 2398 34570 2404 34604
rect 2214 34539 2231 34570
rect 2283 34539 2335 34570
rect 2387 34539 2404 34570
rect 2214 34531 2404 34539
rect 2214 34497 2220 34531
rect 2254 34526 2292 34531
rect 2283 34497 2292 34526
rect 2326 34526 2364 34531
rect 2326 34497 2335 34526
rect 2398 34497 2404 34531
rect 2214 34474 2231 34497
rect 2283 34474 2335 34497
rect 2387 34474 2404 34497
rect 2214 34461 2404 34474
rect 2214 34458 2231 34461
rect 2283 34458 2335 34461
rect 2387 34458 2404 34461
rect 2214 34424 2220 34458
rect 2283 34424 2292 34458
rect 2326 34424 2335 34458
rect 2398 34424 2404 34458
rect 2214 34409 2231 34424
rect 2283 34409 2335 34424
rect 2387 34409 2404 34424
rect 2214 34396 2404 34409
rect 2214 34385 2231 34396
rect 2283 34385 2335 34396
rect 2387 34385 2404 34396
rect 2214 34351 2220 34385
rect 2283 34351 2292 34385
rect 2326 34351 2335 34385
rect 2398 34351 2404 34385
rect 2214 34344 2231 34351
rect 2283 34344 2335 34351
rect 2387 34344 2404 34351
rect 2214 34331 2404 34344
rect 2214 34312 2231 34331
rect 2283 34312 2335 34331
rect 2387 34312 2404 34331
rect 2214 34278 2220 34312
rect 2283 34279 2292 34312
rect 2254 34278 2292 34279
rect 2326 34279 2335 34312
rect 2326 34278 2364 34279
rect 2398 34278 2404 34312
rect 2214 34266 2404 34278
rect 2214 34239 2231 34266
rect 2283 34239 2335 34266
rect 2387 34239 2404 34266
rect 2214 34205 2220 34239
rect 2283 34214 2292 34239
rect 2254 34205 2292 34214
rect 2326 34214 2335 34239
rect 2326 34205 2364 34214
rect 2398 34205 2404 34239
rect 2214 34193 2404 34205
rect 2214 34192 2403 34193
tri 2403 34192 2404 34193 nw
rect 2566 39108 12896 39114
rect 2566 39074 3176 39108
rect 3210 39074 3248 39108
rect 3282 39074 3578 39108
rect 3612 39074 3650 39108
rect 3684 39074 4096 39108
rect 4130 39074 4168 39108
rect 4202 39074 4498 39108
rect 4532 39074 4570 39108
rect 4604 39074 5016 39108
rect 5050 39074 5088 39108
rect 5122 39074 5418 39108
rect 5452 39074 5490 39108
rect 5524 39074 5936 39108
rect 5970 39074 6008 39108
rect 6042 39074 6338 39108
rect 6372 39074 6410 39108
rect 6444 39074 6856 39108
rect 6890 39074 6928 39108
rect 6962 39074 7258 39108
rect 7292 39074 7330 39108
rect 7364 39074 7776 39108
rect 7810 39074 7848 39108
rect 7882 39074 8178 39108
rect 8212 39074 8250 39108
rect 8284 39074 8696 39108
rect 8730 39074 8768 39108
rect 8802 39074 9098 39108
rect 9132 39074 9170 39108
rect 9204 39074 9616 39108
rect 9650 39074 9688 39108
rect 9722 39074 10018 39108
rect 10052 39074 10090 39108
rect 10124 39074 10536 39108
rect 10570 39074 10608 39108
rect 10642 39074 10938 39108
rect 10972 39074 11010 39108
rect 11044 39074 11456 39108
rect 11490 39074 11528 39108
rect 11562 39074 11858 39108
rect 11892 39074 11930 39108
rect 11964 39074 12376 39108
rect 12410 39074 12448 39108
rect 12482 39074 12778 39108
rect 12812 39074 12850 39108
rect 12884 39074 12896 39108
rect 2566 39068 12896 39074
rect 13447 39109 13637 39147
rect 13447 39075 13453 39109
rect 13487 39108 13637 39109
rect 13487 39075 13525 39108
rect 13447 39074 13525 39075
rect 13559 39074 13597 39108
rect 13631 39074 13637 39108
rect 2566 39066 2685 39068
tri 2685 39066 2687 39068 nw
rect 2566 39036 2655 39066
tri 2655 39036 2685 39066 nw
rect 2566 39028 2647 39036
tri 2647 39028 2655 39036 nw
rect 11151 39028 11341 39040
rect 2566 39015 2634 39028
tri 2634 39015 2647 39028 nw
rect 2871 39015 3061 39027
rect 2566 36986 2633 39015
tri 2633 39014 2634 39015 nw
rect 2566 36952 2583 36986
rect 2617 36952 2633 36986
rect 2566 36901 2633 36952
rect 2566 36867 2583 36901
rect 2617 36867 2633 36901
rect 2566 36816 2633 36867
rect 2566 36782 2583 36816
rect 2617 36782 2633 36816
rect 2566 36731 2633 36782
rect 2566 36697 2583 36731
rect 2617 36697 2633 36731
rect 2566 36646 2633 36697
rect 2566 36612 2583 36646
rect 2617 36612 2633 36646
rect 2566 36560 2633 36612
rect 2566 36526 2583 36560
rect 2617 36526 2633 36560
tri 2204 34182 2214 34192 se
rect 2214 34182 2379 34192
tri 1696 34171 1707 34182 se
rect 1707 34171 2074 34182
tri 2074 34171 2085 34182 nw
tri 2193 34171 2204 34182 se
rect 2204 34171 2379 34182
rect 1696 34168 2071 34171
tri 2071 34168 2074 34171 nw
tri 2190 34168 2193 34171 se
rect 2193 34168 2379 34171
tri 2379 34168 2403 34192 nw
rect 1696 34156 2059 34168
tri 2059 34156 2071 34168 nw
tri 2178 34156 2190 34168 se
rect 2190 34156 2341 34168
rect 1696 34144 2033 34156
rect 1696 34110 1702 34144
rect 1736 34110 1808 34144
rect 1842 34130 2033 34144
tri 2033 34130 2059 34156 nw
tri 2152 34130 2178 34156 se
rect 2178 34130 2341 34156
tri 2341 34130 2379 34168 nw
rect 1842 34115 2018 34130
tri 2018 34115 2033 34130 nw
tri 2148 34126 2152 34130 se
rect 2152 34126 2337 34130
tri 2337 34126 2341 34130 nw
rect 2148 34115 2326 34126
tri 2326 34115 2337 34126 nw
rect 1842 34110 2006 34115
rect 1696 34103 2006 34110
tri 2006 34103 2018 34115 nw
rect 2148 34103 2307 34115
rect 1696 34069 1972 34103
tri 1972 34069 2006 34103 nw
rect 2148 34069 2154 34103
rect 2188 34069 2226 34103
rect 2260 34096 2307 34103
tri 2307 34096 2326 34115 nw
rect 2260 34069 2269 34096
rect 1696 34035 1702 34069
rect 1736 34035 1808 34069
rect 1842 34058 1961 34069
tri 1961 34058 1972 34069 nw
rect 2148 34058 2269 34069
tri 2269 34058 2307 34096 nw
rect 1842 34035 1933 34058
rect 1696 34030 1933 34035
tri 1933 34030 1961 34058 nw
rect 2148 34030 2266 34058
tri 2266 34055 2269 34058 nw
rect 1696 33996 1899 34030
tri 1899 33996 1933 34030 nw
rect 2148 33996 2154 34030
rect 2188 33996 2226 34030
rect 2260 33996 2266 34030
rect 1696 33994 1889 33996
rect 1696 33960 1702 33994
rect 1736 33960 1808 33994
rect 1842 33986 1889 33994
tri 1889 33986 1899 33996 nw
rect 1842 33960 1860 33986
rect 1696 33957 1860 33960
tri 1860 33957 1889 33986 nw
rect 2148 33957 2266 33996
rect 1696 33919 1848 33957
tri 1848 33945 1860 33957 nw
rect 1696 33885 1702 33919
rect 1736 33885 1808 33919
rect 1842 33885 1848 33919
rect 1696 33844 1848 33885
rect 1696 33810 1702 33844
rect 1736 33810 1808 33844
rect 1842 33810 1848 33844
rect 1696 33769 1848 33810
rect 1696 33735 1702 33769
rect 1736 33735 1808 33769
rect 1842 33735 1848 33769
rect 1696 33694 1848 33735
rect 1696 33660 1702 33694
rect 1736 33660 1808 33694
rect 1842 33660 1848 33694
rect 1696 33619 1848 33660
rect 1696 33585 1702 33619
rect 1736 33585 1808 33619
rect 1842 33585 1848 33619
rect 1696 33544 1848 33585
rect 1696 33510 1702 33544
rect 1736 33510 1808 33544
rect 1842 33510 1848 33544
rect 1696 33469 1848 33510
rect 1696 33435 1702 33469
rect 1736 33435 1808 33469
rect 1842 33435 1848 33469
rect 1696 33394 1848 33435
rect 1696 33360 1702 33394
rect 1736 33360 1808 33394
rect 1842 33360 1848 33394
rect 1696 33319 1848 33360
rect 1696 33285 1702 33319
rect 1736 33285 1808 33319
rect 1842 33285 1848 33319
rect 1696 33244 1848 33285
rect 1696 33210 1702 33244
rect 1736 33210 1808 33244
rect 1842 33210 1848 33244
rect 1696 33169 1848 33210
rect 1696 33135 1702 33169
rect 1736 33135 1808 33169
rect 1842 33135 1848 33169
rect 1696 33094 1848 33135
rect 1696 33060 1702 33094
rect 1736 33060 1808 33094
rect 1842 33060 1848 33094
rect 1696 33019 1848 33060
rect 1696 32985 1702 33019
rect 1736 32985 1808 33019
rect 1842 32985 1848 33019
rect 1696 32944 1848 32985
rect 1696 32910 1702 32944
rect 1736 32910 1808 32944
rect 1842 32910 1848 32944
rect 1696 32869 1848 32910
rect 1696 32835 1702 32869
rect 1736 32835 1808 32869
rect 1842 32835 1848 32869
rect 1696 32793 1848 32835
rect 1696 32759 1702 32793
rect 1736 32759 1808 32793
rect 1842 32759 1848 32793
rect 1696 32717 1848 32759
rect 1696 32683 1702 32717
rect 1736 32683 1808 32717
rect 1842 32683 1848 32717
rect 1696 32641 1848 32683
rect 1696 32607 1702 32641
rect 1736 32607 1808 32641
rect 1842 32607 1848 32641
rect 1696 32565 1848 32607
rect 1696 32531 1702 32565
rect 1736 32531 1808 32565
rect 1842 32531 1848 32565
rect 1696 32519 1848 32531
rect 2148 33923 2154 33957
rect 2188 33923 2226 33957
rect 2260 33923 2266 33957
rect 2148 33884 2266 33923
rect 2148 33850 2154 33884
rect 2188 33850 2226 33884
rect 2260 33850 2266 33884
rect 2148 33811 2266 33850
rect 2148 33777 2154 33811
rect 2188 33777 2226 33811
rect 2260 33777 2266 33811
rect 2148 33738 2266 33777
rect 2148 33704 2154 33738
rect 2188 33704 2226 33738
rect 2260 33704 2266 33738
rect 2148 33665 2266 33704
rect 2148 33631 2154 33665
rect 2188 33631 2226 33665
rect 2260 33631 2266 33665
rect 2148 33592 2266 33631
rect 2148 33558 2154 33592
rect 2188 33558 2226 33592
rect 2260 33558 2266 33592
rect 2148 33519 2266 33558
rect 2148 33485 2154 33519
rect 2188 33485 2226 33519
rect 2260 33485 2266 33519
rect 2148 33446 2266 33485
rect 2148 33412 2154 33446
rect 2188 33412 2226 33446
rect 2260 33412 2266 33446
rect 2148 33373 2266 33412
rect 2148 33339 2154 33373
rect 2188 33339 2226 33373
rect 2260 33339 2266 33373
rect 2148 33300 2266 33339
rect 2148 33266 2154 33300
rect 2188 33266 2226 33300
rect 2260 33266 2266 33300
rect 2148 33227 2266 33266
rect 2148 33193 2154 33227
rect 2188 33193 2226 33227
rect 2260 33193 2266 33227
rect 2148 33154 2266 33193
rect 2148 33120 2154 33154
rect 2188 33120 2226 33154
rect 2260 33120 2266 33154
rect 2148 33081 2266 33120
rect 2148 33047 2154 33081
rect 2188 33047 2226 33081
rect 2260 33047 2266 33081
rect 2148 33008 2266 33047
rect 2148 32974 2154 33008
rect 2188 32974 2226 33008
rect 2260 32974 2266 33008
rect 2148 32935 2266 32974
rect 2148 32901 2154 32935
rect 2188 32901 2226 32935
rect 2260 32901 2266 32935
rect 2148 32861 2266 32901
rect 2148 32827 2154 32861
rect 2188 32827 2226 32861
rect 2260 32827 2266 32861
rect 2148 32787 2266 32827
rect 2148 32753 2154 32787
rect 2188 32753 2226 32787
rect 2260 32753 2266 32787
rect 2148 32713 2266 32753
rect 2148 32679 2154 32713
rect 2188 32679 2226 32713
rect 2260 32679 2266 32713
rect 2148 32639 2266 32679
rect 2148 32605 2154 32639
rect 2188 32605 2226 32639
rect 2260 32605 2266 32639
rect 2148 32565 2266 32605
rect 2148 32531 2154 32565
rect 2188 32531 2226 32565
rect 2260 32531 2266 32565
rect 2148 32519 2266 32531
tri 2564 32292 2566 32294 se
rect 2566 32292 2633 36526
rect 2871 39009 2877 39015
rect 3055 39009 3061 39015
rect 2871 38957 2872 39009
rect 3060 38957 3061 39009
rect 2871 38944 2877 38957
rect 3055 38944 3061 38957
rect 2871 38892 2872 38944
rect 3060 38892 3061 38944
rect 2871 38879 2877 38892
rect 3055 38879 3061 38892
rect 2871 38827 2872 38879
rect 3060 38827 3061 38879
rect 2871 38814 2877 38827
rect 3055 38814 3061 38827
rect 2871 38762 2872 38814
rect 3060 38762 3061 38814
rect 2871 38749 2877 38762
rect 3055 38749 3061 38762
rect 2871 38697 2872 38749
rect 3060 38697 3061 38749
rect 2871 38684 2877 38697
rect 3055 38684 3061 38697
rect 2871 38632 2872 38684
rect 3060 38632 3061 38684
rect 2871 38619 2877 38632
rect 3055 38619 3061 38632
rect 2871 38567 2872 38619
rect 3060 38567 3061 38619
rect 2871 38554 2877 38567
rect 3055 38554 3061 38567
rect 2871 38502 2872 38554
rect 3060 38502 3061 38554
rect 2871 38490 2877 38502
rect 3055 38490 3061 38502
rect 2871 38438 2872 38490
rect 3060 38438 3061 38490
rect 2871 38426 2877 38438
rect 3055 38426 3061 38438
rect 2871 38374 2872 38426
rect 3060 38374 3061 38426
rect 2871 38362 2877 38374
rect 3055 38362 3061 38374
rect 2871 38310 2872 38362
rect 3060 38310 3061 38362
rect 2871 38298 2877 38310
rect 3055 38298 3061 38310
rect 2871 38246 2872 38298
rect 3060 38246 3061 38298
rect 2871 38234 2877 38246
rect 3055 38234 3061 38246
rect 2871 38182 2872 38234
rect 3060 38182 3061 38234
rect 2871 38170 2877 38182
rect 3055 38170 3061 38182
rect 2871 38118 2872 38170
rect 3060 38118 3061 38170
rect 2871 37541 2877 38118
rect 3055 37541 3061 38118
rect 3791 39015 3981 39027
rect 3791 39009 3797 39015
rect 3975 39009 3981 39015
rect 3791 38957 3792 39009
rect 3980 38957 3981 39009
rect 3791 38944 3797 38957
rect 3975 38944 3981 38957
rect 3791 38892 3792 38944
rect 3980 38892 3981 38944
rect 3791 38879 3797 38892
rect 3975 38879 3981 38892
rect 3791 38827 3792 38879
rect 3980 38827 3981 38879
rect 3791 38814 3797 38827
rect 3975 38814 3981 38827
rect 3791 38762 3792 38814
rect 3980 38762 3981 38814
rect 3791 38749 3797 38762
rect 3975 38749 3981 38762
rect 3791 38697 3792 38749
rect 3980 38697 3981 38749
rect 3791 38684 3797 38697
rect 3975 38684 3981 38697
rect 3791 38632 3792 38684
rect 3980 38632 3981 38684
rect 3791 38619 3797 38632
rect 3975 38619 3981 38632
rect 3791 38567 3792 38619
rect 3980 38567 3981 38619
rect 3791 38554 3797 38567
rect 3975 38554 3981 38567
rect 3791 38502 3792 38554
rect 3980 38502 3981 38554
rect 3791 38490 3797 38502
rect 3975 38490 3981 38502
rect 3791 38438 3792 38490
rect 3980 38438 3981 38490
rect 3791 38426 3797 38438
rect 3975 38426 3981 38438
rect 3791 38374 3792 38426
rect 3980 38374 3981 38426
rect 3791 38362 3797 38374
rect 3975 38362 3981 38374
rect 3791 38310 3792 38362
rect 3980 38310 3981 38362
rect 3791 38298 3797 38310
rect 3975 38298 3981 38310
rect 3791 38246 3792 38298
rect 3980 38246 3981 38298
rect 3791 38234 3797 38246
rect 3975 38234 3981 38246
rect 3791 38182 3792 38234
rect 3980 38182 3981 38234
rect 3791 38170 3797 38182
rect 3975 38170 3981 38182
rect 3791 38118 3792 38170
rect 3980 38118 3981 38170
rect 2871 37502 3061 37541
rect 2871 37468 2877 37502
rect 2911 37468 2949 37502
rect 2983 37468 3021 37502
rect 3055 37468 3061 37502
rect 2871 37429 3061 37468
rect 2871 37395 2877 37429
rect 2911 37395 2949 37429
rect 2983 37395 3021 37429
rect 3055 37395 3061 37429
rect 2871 37356 3061 37395
rect 2871 37322 2877 37356
rect 2911 37322 2949 37356
rect 2983 37322 3021 37356
rect 3055 37322 3061 37356
rect 2871 37283 3061 37322
rect 2871 37249 2877 37283
rect 2911 37249 2949 37283
rect 2983 37249 3021 37283
rect 3055 37249 3061 37283
rect 2871 37210 3061 37249
rect 2871 37176 2877 37210
rect 2911 37176 2949 37210
rect 2983 37176 3021 37210
rect 3055 37176 3061 37210
rect 2871 37137 3061 37176
rect 2871 37103 2877 37137
rect 2911 37103 2949 37137
rect 2983 37103 3021 37137
rect 3055 37103 3061 37137
rect 2871 36368 3061 37103
rect 2871 36316 2872 36368
rect 2924 36316 2940 36368
rect 2992 36316 3008 36368
rect 3060 36316 3061 36368
rect 2871 36304 3061 36316
rect 2871 36252 2872 36304
rect 2924 36252 2940 36304
rect 2992 36252 3008 36304
rect 3060 36252 3061 36304
rect 2871 36239 3061 36252
rect 2871 36187 2872 36239
rect 2924 36187 2940 36239
rect 2992 36187 3008 36239
rect 3060 36187 3061 36239
rect 2871 36184 2943 36187
rect 2977 36184 3021 36187
rect 3055 36184 3061 36187
rect 2871 36174 3061 36184
rect 2871 36122 2872 36174
rect 2924 36122 2940 36174
rect 2992 36122 3008 36174
rect 3060 36122 3061 36174
rect 2871 36112 2943 36122
rect 2977 36112 3021 36122
rect 3055 36112 3061 36122
rect 2871 36109 3061 36112
rect 2871 36057 2872 36109
rect 2924 36057 2940 36109
rect 2992 36057 3008 36109
rect 3060 36057 3061 36109
rect 2871 36044 2943 36057
rect 2977 36044 3021 36057
rect 3055 36044 3061 36057
rect 2871 35992 2872 36044
rect 2924 35992 2940 36044
rect 2992 35992 3008 36044
rect 3060 35992 3061 36044
rect 2871 35979 2943 35992
rect 2977 35979 3021 35992
rect 3055 35979 3061 35992
rect 2871 35927 2872 35979
rect 2924 35927 2940 35979
rect 2992 35927 3008 35979
rect 3060 35927 3061 35979
rect 2871 35914 2943 35927
rect 2977 35914 3021 35927
rect 3055 35914 3061 35927
rect 2871 35862 2872 35914
rect 2924 35862 2940 35914
rect 2992 35862 3008 35914
rect 3060 35862 3061 35914
rect 2871 35858 3061 35862
rect 2871 35849 2943 35858
rect 2977 35849 3021 35858
rect 3055 35849 3061 35858
rect 2871 35797 2872 35849
rect 2924 35797 2940 35849
rect 2992 35797 3008 35849
rect 3060 35797 3061 35849
rect 2871 35786 3061 35797
rect 2871 35784 2943 35786
rect 2977 35784 3021 35786
rect 3055 35784 3061 35786
rect 2871 35732 2872 35784
rect 2924 35732 2940 35784
rect 2992 35732 3008 35784
rect 3060 35732 3061 35784
rect 2871 35719 3061 35732
rect 2871 35667 2872 35719
rect 2924 35667 2940 35719
rect 2992 35667 3008 35719
rect 3060 35667 3061 35719
rect 2871 35654 3061 35667
rect 2871 35602 2872 35654
rect 2924 35602 2940 35654
rect 2992 35602 3008 35654
rect 3060 35602 3061 35654
rect 2871 35589 3061 35602
rect 2871 35537 2872 35589
rect 2924 35537 2940 35589
rect 2992 35537 3008 35589
rect 3060 35537 3061 35589
rect 2871 35536 2943 35537
rect 2977 35536 3021 35537
rect 3055 35536 3061 35537
rect 2871 35524 3061 35536
rect 2871 35472 2872 35524
rect 2924 35472 2940 35524
rect 2992 35472 3008 35524
rect 3060 35472 3061 35524
rect 2871 35464 2943 35472
rect 2977 35464 3021 35472
rect 3055 35464 3061 35472
rect 2871 35459 3061 35464
rect 2871 35407 2872 35459
rect 2924 35407 2940 35459
rect 2992 35407 3008 35459
rect 3060 35407 3061 35459
rect 2871 35394 2943 35407
rect 2977 35394 3021 35407
rect 3055 35394 3061 35407
rect 2871 35342 2872 35394
rect 2924 35342 2940 35394
rect 2992 35342 3008 35394
rect 3060 35342 3061 35394
rect 2871 35329 2943 35342
rect 2977 35329 3021 35342
rect 3055 35329 3061 35342
rect 2871 35277 2872 35329
rect 2924 35277 2940 35329
rect 2992 35277 3008 35329
rect 3060 35277 3061 35329
rect 2871 35264 2943 35277
rect 2977 35264 3021 35277
rect 3055 35264 3061 35277
rect 2871 35212 2872 35264
rect 2924 35212 2940 35264
rect 2992 35212 3008 35264
rect 3060 35212 3061 35264
rect 2871 35210 3061 35212
rect 2871 35199 2943 35210
rect 2977 35199 3021 35210
rect 3055 35199 3061 35210
rect 2871 35147 2872 35199
rect 2924 35147 2940 35199
rect 2992 35147 3008 35199
rect 3060 35147 3061 35199
rect 2871 35138 3061 35147
rect 2871 35134 2943 35138
rect 2977 35134 3021 35138
rect 3055 35134 3061 35138
rect 2871 35082 2872 35134
rect 2924 35082 2940 35134
rect 2992 35082 3008 35134
rect 3060 35082 3061 35134
rect 2871 35069 3061 35082
rect 2871 35017 2872 35069
rect 2924 35017 2940 35069
rect 2992 35017 3008 35069
rect 3060 35017 3061 35069
rect 2871 35004 3061 35017
rect 2871 34952 2872 35004
rect 2924 34952 2940 35004
rect 2992 34952 3008 35004
rect 3060 34952 3061 35004
rect 2871 34939 3061 34952
rect 2871 34887 2872 34939
rect 2924 34887 2940 34939
rect 2992 34887 3008 34939
rect 3060 34887 3061 34939
rect 2871 34874 3061 34887
rect 2871 34822 2872 34874
rect 2924 34822 2940 34874
rect 2992 34822 3008 34874
rect 3060 34822 3061 34874
rect 2871 34816 2943 34822
rect 2977 34816 3021 34822
rect 3055 34816 3061 34822
rect 2871 34809 3061 34816
rect 2871 34757 2872 34809
rect 2924 34757 2940 34809
rect 2992 34757 3008 34809
rect 3060 34757 3061 34809
rect 2871 34744 2943 34757
rect 2977 34744 3021 34757
rect 3055 34744 3061 34757
rect 2871 34692 2872 34744
rect 2924 34692 2940 34744
rect 2992 34692 3008 34744
rect 3060 34692 3061 34744
rect 2871 34679 2943 34692
rect 2977 34679 3021 34692
rect 3055 34679 3061 34692
rect 2871 34627 2872 34679
rect 2924 34627 2940 34679
rect 2992 34627 3008 34679
rect 3060 34627 3061 34679
rect 2871 34614 2943 34627
rect 2977 34614 3021 34627
rect 3055 34614 3061 34627
rect 2871 34562 2872 34614
rect 2924 34562 2940 34614
rect 2992 34562 3008 34614
rect 3060 34562 3061 34614
rect 2871 34528 2943 34562
rect 2977 34528 3021 34562
rect 3055 34528 3061 34562
rect 2871 34490 3061 34528
rect 2871 34456 2943 34490
rect 2977 34456 3021 34490
rect 3055 34456 3061 34490
rect 2871 34418 3061 34456
rect 2871 34384 2943 34418
rect 2977 34384 3021 34418
rect 3055 34384 3061 34418
rect 2871 34346 3061 34384
rect 2871 34312 2943 34346
rect 2977 34312 3021 34346
rect 3055 34312 3061 34346
rect 2871 34274 3061 34312
rect 2871 34240 2943 34274
rect 2977 34240 3021 34274
rect 3055 34240 3061 34274
rect 2871 34202 3061 34240
rect 2871 34177 2943 34202
tri 2871 34168 2880 34177 ne
rect 2880 34168 2943 34177
rect 2977 34168 3021 34202
rect 3055 34168 3061 34202
tri 2880 34130 2918 34168 ne
rect 2918 34130 3061 34168
tri 2918 34111 2937 34130 ne
rect 2937 34096 2943 34130
rect 2977 34096 3021 34130
rect 3055 34096 3061 34130
rect 2937 34058 3061 34096
rect 2937 34024 2943 34058
rect 2977 34024 3021 34058
rect 3055 34024 3061 34058
rect 2937 33986 3061 34024
rect 2937 33952 2943 33986
rect 2977 33952 3021 33986
rect 3055 33952 3061 33986
rect 2937 33914 3061 33952
rect 2937 33880 2943 33914
rect 2977 33880 3021 33914
rect 3055 33880 3061 33914
rect 2937 33842 3061 33880
rect 2937 33808 2943 33842
rect 2977 33808 3021 33842
rect 3055 33808 3061 33842
rect 2937 33770 3061 33808
rect 2937 33736 2943 33770
rect 2977 33736 3021 33770
rect 3055 33736 3061 33770
rect 2937 33698 3061 33736
rect 2937 33664 2943 33698
rect 2977 33664 3021 33698
rect 3055 33664 3061 33698
rect 2937 33626 3061 33664
rect 2937 33592 2943 33626
rect 2977 33592 3021 33626
rect 3055 33592 3061 33626
rect 2937 33554 3061 33592
rect 2937 33520 2943 33554
rect 2977 33520 3021 33554
rect 3055 33520 3061 33554
rect 2937 33482 3061 33520
rect 2937 33448 2943 33482
rect 2977 33448 3021 33482
rect 3055 33448 3061 33482
rect 2937 33410 3061 33448
rect 2937 33376 2943 33410
rect 2977 33376 3021 33410
rect 3055 33376 3061 33410
rect 2937 33338 3061 33376
rect 2937 33304 2943 33338
rect 2977 33304 3021 33338
rect 3055 33304 3061 33338
rect 2937 33266 3061 33304
rect 2937 33232 2943 33266
rect 2977 33232 3021 33266
rect 3055 33232 3061 33266
rect 2937 33194 3061 33232
rect 2937 33160 2943 33194
rect 2977 33160 3021 33194
rect 3055 33160 3061 33194
rect 2937 33121 3061 33160
rect 2937 33087 2943 33121
rect 2977 33087 3021 33121
rect 3055 33087 3061 33121
rect 2937 33048 3061 33087
rect 2937 33014 2943 33048
rect 2977 33014 3021 33048
rect 3055 33014 3061 33048
rect 2937 32975 3061 33014
rect 2937 32941 2943 32975
rect 2977 32941 3021 32975
rect 3055 32941 3061 32975
rect 2937 32902 3061 32941
rect 2937 32868 2943 32902
rect 2977 32868 3021 32902
rect 3055 32868 3061 32902
rect 2937 32829 3061 32868
rect 2937 32795 2943 32829
rect 2977 32795 3021 32829
rect 3055 32795 3061 32829
rect 2937 32756 3061 32795
rect 2937 32722 2943 32756
rect 2977 32722 3021 32756
rect 3055 32722 3061 32756
rect 2937 32683 3061 32722
rect 2937 32649 2943 32683
rect 2977 32649 3021 32683
rect 3055 32649 3061 32683
rect 2937 32610 3061 32649
rect 2937 32576 2943 32610
rect 2977 32576 3021 32610
rect 3055 32576 3061 32610
rect 2937 32537 3061 32576
rect 2937 32503 2943 32537
rect 2977 32503 3021 32537
rect 3055 32503 3061 32537
rect 2937 32491 3061 32503
rect 3361 37997 3491 38003
rect 3413 37945 3439 37997
rect 3361 37929 3491 37945
rect 3413 37877 3439 37929
rect 3361 37861 3491 37877
rect 3413 37809 3439 37861
rect 3361 37793 3491 37809
rect 3413 37741 3439 37793
rect 3361 37725 3491 37741
rect 3413 37673 3439 37725
rect 3361 37657 3491 37673
rect 3413 37605 3439 37657
rect 3361 37589 3491 37605
rect 3413 37537 3439 37589
rect 3361 37521 3491 37537
rect 3413 37469 3439 37521
rect 3361 37453 3491 37469
rect 3413 37401 3439 37453
rect 3361 37385 3491 37401
rect 3413 37333 3439 37385
rect 3361 37318 3491 37333
rect 3413 37266 3439 37318
rect 3361 37251 3491 37266
rect 3413 37199 3439 37251
rect 3361 37184 3491 37199
rect 3413 37132 3439 37184
rect 3361 37117 3491 37132
rect 3413 37065 3439 37117
rect 3361 34225 3491 37065
rect 3413 34173 3439 34225
rect 3361 34161 3491 34173
rect 3413 34109 3439 34161
rect 3361 34097 3491 34109
rect 3413 34045 3439 34097
rect 3361 34033 3491 34045
rect 3413 33981 3439 34033
rect 3361 33969 3491 33981
rect 3413 33917 3439 33969
rect 3361 33905 3491 33917
rect 3413 33853 3439 33905
rect 3361 33841 3491 33853
rect 3413 33789 3439 33841
rect 3361 33777 3491 33789
rect 3413 33725 3439 33777
rect 3361 33713 3491 33725
rect 3413 33661 3439 33713
rect 3361 33649 3491 33661
rect 3413 33597 3439 33649
rect 3361 33585 3491 33597
rect 3413 33533 3439 33585
rect 3361 33521 3491 33533
rect 3413 33469 3439 33521
rect 3361 33457 3491 33469
rect 3413 33405 3439 33457
rect 3361 33393 3491 33405
rect 3413 33341 3439 33393
rect 3361 33329 3491 33341
rect 3413 33277 3439 33329
rect 3361 33264 3491 33277
rect 3413 33212 3439 33264
rect 3361 33199 3491 33212
rect 3413 33147 3439 33199
rect 3361 33134 3491 33147
rect 3413 33082 3439 33134
rect 3361 33069 3491 33082
rect 3413 33017 3439 33069
rect 3361 33004 3491 33017
rect 3413 32952 3439 33004
rect 3361 32939 3491 32952
rect 3413 32887 3439 32939
rect 3361 32874 3491 32887
rect 3413 32822 3439 32874
rect 3361 32809 3491 32822
rect 3413 32757 3439 32809
rect 3361 32744 3491 32757
rect 3413 32692 3439 32744
rect 3361 32679 3491 32692
rect 3413 32627 3439 32679
rect 3361 32614 3491 32627
rect 3413 32562 3439 32614
rect 3361 32549 3491 32562
rect 3413 32497 3439 32549
tri 2633 32292 2634 32293 sw
tri 2530 32258 2564 32292 se
rect 2564 32258 2634 32292
tri 2634 32258 2668 32292 sw
tri 2526 32254 2530 32258 se
rect 2530 32254 2668 32258
tri 2668 32254 2672 32258 sw
tri 2522 32250 2526 32254 se
rect 2526 32250 2672 32254
rect 1418 32220 1498 32250
tri 1498 32220 1528 32250 sw
tri 2492 32220 2522 32250 se
rect 2522 32220 2672 32250
tri 2672 32220 2706 32254 sw
rect 1418 32219 1528 32220
tri 1528 32219 1529 32220 sw
tri 2491 32219 2492 32220 se
rect 2492 32219 2706 32220
tri 2706 32219 2707 32220 sw
rect 1418 32216 1529 32219
tri 1529 32216 1532 32219 sw
tri 2488 32216 2491 32219 se
rect 2491 32216 2707 32219
tri 2707 32216 2710 32219 sw
rect 1418 32210 2710 32216
rect 1418 32176 2494 32210
rect 2528 32176 2579 32210
rect 2613 32176 2664 32210
rect 2698 32176 2710 32210
rect 1418 32138 2710 32176
rect 1418 32104 2494 32138
rect 2528 32104 2579 32138
rect 2613 32104 2664 32138
rect 2698 32104 2710 32138
rect 1418 32098 2710 32104
rect 1418 32076 1510 32098
tri 1510 32076 1532 32098 nw
rect 1418 32073 1507 32076
tri 1507 32073 1510 32076 nw
rect 1418 26341 1498 32073
tri 1498 32064 1507 32073 nw
rect 1834 31783 1986 31795
rect 1834 31749 1840 31783
rect 1874 31749 1946 31783
rect 1980 31749 1986 31783
rect 1834 31711 1986 31749
rect 1834 31677 1840 31711
rect 1874 31677 1946 31711
rect 1980 31677 1986 31711
rect 1834 31639 1986 31677
rect 1834 31638 1946 31639
rect 1834 31604 1840 31638
rect 1874 31605 1946 31638
rect 1980 31605 1986 31639
rect 1874 31604 1986 31605
rect 1834 31567 1986 31604
rect 1834 31565 1946 31567
rect 1834 31531 1840 31565
rect 1874 31533 1946 31565
rect 1980 31533 1986 31567
rect 1874 31531 1986 31533
rect 1834 31495 1986 31531
rect 1834 31492 1946 31495
rect 1834 31458 1840 31492
rect 1874 31461 1946 31492
rect 1980 31461 1986 31495
rect 1874 31458 1986 31461
rect 1834 31423 1986 31458
rect 1834 31419 1946 31423
rect 1834 31385 1840 31419
rect 1874 31389 1946 31419
rect 1980 31389 1986 31423
rect 1874 31385 1986 31389
rect 1834 31351 1986 31385
rect 1834 31346 1946 31351
rect 1834 31312 1840 31346
rect 1874 31317 1946 31346
rect 1980 31317 1986 31351
rect 1874 31312 1986 31317
rect 1834 31279 1986 31312
rect 1834 31273 1946 31279
rect 1834 31239 1840 31273
rect 1874 31245 1946 31273
rect 1980 31245 1986 31279
rect 1874 31239 1986 31245
rect 1834 31207 1986 31239
rect 1834 31200 1946 31207
rect 1834 31166 1840 31200
rect 1874 31173 1946 31200
rect 1980 31173 1986 31207
rect 1874 31166 1986 31173
rect 1834 31135 1986 31166
rect 1834 31127 1946 31135
rect 1834 31093 1840 31127
rect 1874 31101 1946 31127
rect 1980 31101 1986 31135
rect 1874 31093 1986 31101
rect 1834 31063 1986 31093
rect 1834 31054 1946 31063
rect 1834 31020 1840 31054
rect 1874 31029 1946 31054
rect 1980 31029 1986 31063
rect 1874 31020 1986 31029
rect 1834 30991 1986 31020
rect 1834 30981 1946 30991
rect 1834 30947 1840 30981
rect 1874 30957 1946 30981
rect 1980 30957 1986 30991
rect 1874 30947 1986 30957
rect 1834 30919 1986 30947
rect 1834 30908 1946 30919
rect 1834 30874 1840 30908
rect 1874 30885 1946 30908
rect 1980 30885 1986 30919
rect 1874 30874 1986 30885
rect 1834 30847 1986 30874
rect 1834 30835 1946 30847
rect 1834 30801 1840 30835
rect 1874 30813 1946 30835
rect 1980 30813 1986 30847
rect 1874 30801 1986 30813
rect 1834 30775 1986 30801
rect 1834 30762 1946 30775
rect 1834 30728 1840 30762
rect 1874 30741 1946 30762
rect 1980 30741 1986 30775
rect 1874 30728 1986 30741
rect 1834 30703 1986 30728
rect 1834 30689 1946 30703
rect 1834 30655 1840 30689
rect 1874 30669 1946 30689
rect 1980 30669 1986 30703
rect 1874 30655 1986 30669
rect 1834 30631 1986 30655
rect 1834 30616 1946 30631
rect 1834 30582 1840 30616
rect 1874 30597 1946 30616
rect 1980 30597 1986 30631
rect 1874 30582 1986 30597
rect 1834 30559 1986 30582
rect 1834 30543 1946 30559
rect 1834 30509 1840 30543
rect 1874 30525 1946 30543
rect 1980 30525 1986 30559
rect 1874 30509 1986 30525
rect 1834 30487 1986 30509
rect 1834 30470 1946 30487
rect 1834 30436 1840 30470
rect 1874 30453 1946 30470
rect 1980 30453 1986 30487
rect 1874 30436 1986 30453
rect 1834 30415 1986 30436
rect 1834 30397 1946 30415
rect 1834 30363 1840 30397
rect 1874 30381 1946 30397
rect 1980 30381 1986 30415
rect 1874 30363 1986 30381
rect 1834 30343 1986 30363
rect 1834 30324 1946 30343
rect 1834 30290 1840 30324
rect 1874 30309 1946 30324
rect 1980 30309 1986 30343
rect 1874 30290 1986 30309
rect 1834 30271 1986 30290
rect 1834 30251 1946 30271
rect 1834 30217 1840 30251
rect 1874 30237 1946 30251
rect 1980 30237 1986 30271
rect 1874 30217 1986 30237
rect 1834 30199 1986 30217
rect 1834 30178 1946 30199
rect 1834 30144 1840 30178
rect 1874 30165 1946 30178
rect 1980 30165 1986 30199
rect 1874 30144 1986 30165
rect 1834 30127 1986 30144
rect 1834 30105 1946 30127
rect 1834 30071 1840 30105
rect 1874 30093 1946 30105
rect 1980 30093 1986 30127
rect 1874 30071 1986 30093
rect 1834 30055 1986 30071
rect 1834 30032 1946 30055
rect 1834 29998 1840 30032
rect 1874 30021 1946 30032
rect 1980 30021 1986 30055
rect 1874 29998 1986 30021
rect 1834 29983 1986 29998
rect 1834 29959 1946 29983
rect 1834 29925 1840 29959
rect 1874 29949 1946 29959
rect 1980 29949 1986 29983
rect 1874 29925 1986 29949
rect 1834 29911 1986 29925
rect 1834 29886 1946 29911
rect 1834 29852 1840 29886
rect 1874 29877 1946 29886
rect 1980 29877 1986 29911
rect 1874 29852 1986 29877
rect 1834 29839 1986 29852
rect 1834 29813 1946 29839
rect 1834 29779 1840 29813
rect 1874 29805 1946 29813
rect 1980 29805 1986 29839
rect 1874 29779 1986 29805
rect 1834 29767 1986 29779
rect 1834 29740 1946 29767
rect 1834 29706 1840 29740
rect 1874 29733 1946 29740
rect 1980 29733 1986 29767
rect 1874 29706 1986 29733
rect 1834 29695 1986 29706
rect 1834 29667 1946 29695
rect 1834 29633 1840 29667
rect 1874 29661 1946 29667
rect 1980 29661 1986 29695
rect 1874 29633 1986 29661
rect 1834 29623 1986 29633
rect 1834 29594 1946 29623
rect 1834 29560 1840 29594
rect 1874 29589 1946 29594
rect 1980 29589 1986 29623
rect 1874 29560 1986 29589
rect 1834 29551 1986 29560
rect 1834 29521 1946 29551
rect 1834 29487 1840 29521
rect 1874 29517 1946 29521
rect 1980 29517 1986 29551
rect 1874 29487 1986 29517
rect 1834 29479 1986 29487
rect 1834 29448 1946 29479
rect 1834 29414 1840 29448
rect 1874 29445 1946 29448
rect 1980 29445 1986 29479
rect 1874 29414 1986 29445
rect 1834 29407 1986 29414
rect 1834 29375 1946 29407
rect 1834 29341 1840 29375
rect 1874 29373 1946 29375
rect 1980 29373 1986 29407
rect 1874 29341 1986 29373
rect 1834 29335 1986 29341
rect 1834 29302 1946 29335
rect 1834 29268 1840 29302
rect 1874 29301 1946 29302
rect 1980 29301 1986 29335
rect 1874 29268 1986 29301
rect 1834 29263 1986 29268
rect 1834 29229 1946 29263
rect 1980 29229 1986 29263
rect 1834 29195 1840 29229
rect 1874 29195 1986 29229
rect 1834 29190 1986 29195
rect 1834 29156 1946 29190
rect 1980 29156 1986 29190
rect 1834 29122 1840 29156
rect 1874 29122 1986 29156
rect 1834 29117 1986 29122
rect 1834 29083 1946 29117
rect 1980 29083 1986 29117
rect 1834 29049 1840 29083
rect 1874 29049 1986 29083
rect 1834 29044 1986 29049
rect 1834 29010 1946 29044
rect 1980 29010 1986 29044
rect 1834 28976 1840 29010
rect 1874 28976 1986 29010
rect 1834 28971 1986 28976
rect 1834 28937 1946 28971
rect 1980 28937 1986 28971
rect 1834 28903 1840 28937
rect 1874 28903 1986 28937
rect 1834 28898 1986 28903
rect 1834 28864 1946 28898
rect 1980 28864 1986 28898
rect 1834 28830 1840 28864
rect 1874 28830 1986 28864
rect 1834 28825 1986 28830
rect 1834 28791 1946 28825
rect 1980 28791 1986 28825
rect 1834 28757 1840 28791
rect 1874 28757 1986 28791
rect 1834 28752 1986 28757
rect 1834 28718 1946 28752
rect 1980 28718 1986 28752
rect 1834 28684 1840 28718
rect 1874 28684 1986 28718
rect 1834 28679 1986 28684
rect 1834 28645 1946 28679
rect 1980 28645 1986 28679
rect 1834 28611 1840 28645
rect 1874 28611 1986 28645
rect 1834 28606 1986 28611
rect 1834 28572 1946 28606
rect 1980 28572 1986 28606
rect 1834 28538 1840 28572
rect 1874 28538 1986 28572
rect 1834 28533 1986 28538
rect 1834 28499 1946 28533
rect 1980 28499 1986 28533
rect 1834 28465 1840 28499
rect 1874 28465 1986 28499
rect 1834 28460 1986 28465
rect 1834 28426 1946 28460
rect 1980 28426 1986 28460
rect 1834 28392 1840 28426
rect 1874 28392 1986 28426
rect 1834 28387 1986 28392
rect 1834 28353 1946 28387
rect 1980 28353 1986 28387
rect 1834 28319 1840 28353
rect 1874 28319 1986 28353
rect 1834 28314 1986 28319
rect 1834 28280 1946 28314
rect 1980 28280 1986 28314
rect 1834 28246 1840 28280
rect 1874 28246 1986 28280
rect 1834 28241 1986 28246
rect 1834 28207 1946 28241
rect 1980 28207 1986 28241
rect 1834 28173 1840 28207
rect 1874 28173 1986 28207
rect 1834 28168 1986 28173
rect 1834 28134 1946 28168
rect 1980 28134 1986 28168
rect 1834 28100 1840 28134
rect 1874 28100 1986 28134
rect 1834 28095 1986 28100
rect 1834 28061 1946 28095
rect 1980 28061 1986 28095
rect 1834 28027 1840 28061
rect 1874 28027 1986 28061
rect 1834 28022 1986 28027
rect 1834 27988 1946 28022
rect 1980 27988 1986 28022
rect 1834 27954 1840 27988
rect 1874 27954 1986 27988
rect 1834 27949 1986 27954
rect 1834 27915 1946 27949
rect 1980 27915 1986 27949
rect 1834 27881 1840 27915
rect 1874 27881 1986 27915
rect 1834 27876 1986 27881
rect 1834 27842 1946 27876
rect 1980 27842 1986 27876
rect 1834 27808 1840 27842
rect 1874 27808 1986 27842
rect 1834 27803 1986 27808
rect 1834 27769 1946 27803
rect 1980 27769 1986 27803
rect 1834 27735 1840 27769
rect 1874 27735 1986 27769
rect 1834 27730 1986 27735
rect 1834 27696 1946 27730
rect 1980 27696 1986 27730
rect 1834 27662 1840 27696
rect 1874 27662 1986 27696
rect 1834 27657 1986 27662
rect 1834 27623 1946 27657
rect 1980 27623 1986 27657
rect 1834 27589 1840 27623
rect 1874 27589 1986 27623
rect 1834 27584 1986 27589
rect 1834 27550 1946 27584
rect 1980 27550 1986 27584
rect 1834 27516 1840 27550
rect 1874 27516 1986 27550
rect 1834 27511 1986 27516
rect 1834 27477 1946 27511
rect 1980 27477 1986 27511
rect 1834 27443 1840 27477
rect 1874 27443 1986 27477
rect 1834 27438 1986 27443
rect 1834 27404 1946 27438
rect 1980 27404 1986 27438
rect 1834 27370 1840 27404
rect 1874 27370 1986 27404
rect 1834 27365 1986 27370
rect 1834 27331 1946 27365
rect 1980 27331 1986 27365
rect 1834 27297 1840 27331
rect 1874 27297 1986 27331
rect 1834 27292 1986 27297
rect 1834 27258 1946 27292
rect 1980 27258 1986 27292
rect 1834 27224 1840 27258
rect 1874 27224 1986 27258
rect 1834 27219 1986 27224
rect 1834 27185 1946 27219
rect 1980 27185 1986 27219
rect 1834 27151 1840 27185
rect 1874 27151 1986 27185
rect 1834 27146 1986 27151
rect 1834 27112 1946 27146
rect 1980 27112 1986 27146
rect 1834 27078 1840 27112
rect 1874 27078 1986 27112
rect 2308 31783 2426 31795
rect 2308 30381 2314 31783
rect 2420 30381 2426 31783
rect 2308 30342 2426 30381
rect 2308 30308 2314 30342
rect 2348 30308 2386 30342
rect 2420 30308 2426 30342
rect 2308 30269 2426 30308
rect 2308 30235 2314 30269
rect 2348 30235 2386 30269
rect 2420 30235 2426 30269
rect 2308 30196 2426 30235
rect 2308 30162 2314 30196
rect 2348 30162 2386 30196
rect 2420 30162 2426 30196
rect 2308 30123 2426 30162
rect 2308 30089 2314 30123
rect 2348 30089 2386 30123
rect 2420 30089 2426 30123
rect 2308 30050 2426 30089
rect 2308 30016 2314 30050
rect 2348 30016 2386 30050
rect 2420 30016 2426 30050
rect 2308 29977 2426 30016
rect 2308 29943 2314 29977
rect 2348 29943 2386 29977
rect 2420 29943 2426 29977
rect 2308 29904 2426 29943
rect 2308 29870 2314 29904
rect 2348 29870 2386 29904
rect 2420 29870 2426 29904
rect 2308 29831 2426 29870
rect 2308 29797 2314 29831
rect 2348 29797 2386 29831
rect 2420 29797 2426 29831
rect 2308 29758 2426 29797
rect 2308 29724 2314 29758
rect 2348 29724 2386 29758
rect 2420 29724 2426 29758
rect 2308 29685 2426 29724
rect 2308 29651 2314 29685
rect 2348 29651 2386 29685
rect 2420 29651 2426 29685
rect 2308 29612 2426 29651
rect 2308 29578 2314 29612
rect 2348 29578 2386 29612
rect 2420 29578 2426 29612
rect 2308 29539 2426 29578
rect 2308 29505 2314 29539
rect 2348 29505 2386 29539
rect 2420 29505 2426 29539
rect 2308 29466 2426 29505
rect 2308 29432 2314 29466
rect 2348 29432 2386 29466
rect 2420 29432 2426 29466
rect 2308 29393 2426 29432
rect 2308 29359 2314 29393
rect 2348 29359 2386 29393
rect 2420 29359 2426 29393
rect 2308 29320 2426 29359
rect 2308 29286 2314 29320
rect 2348 29286 2386 29320
rect 2420 29286 2426 29320
rect 2308 29247 2426 29286
rect 2308 29213 2314 29247
rect 2348 29213 2386 29247
rect 2420 29213 2426 29247
rect 2308 29174 2426 29213
rect 2308 29140 2314 29174
rect 2348 29140 2386 29174
rect 2420 29140 2426 29174
rect 2308 29101 2426 29140
rect 2308 29067 2314 29101
rect 2348 29067 2386 29101
rect 2420 29067 2426 29101
rect 2308 29028 2426 29067
rect 2308 28994 2314 29028
rect 2348 28994 2386 29028
rect 2420 28994 2426 29028
rect 2308 28955 2426 28994
rect 2308 28921 2314 28955
rect 2348 28921 2386 28955
rect 2420 28921 2426 28955
rect 2308 28882 2426 28921
rect 2308 28848 2314 28882
rect 2348 28848 2386 28882
rect 2420 28848 2426 28882
rect 2308 28809 2426 28848
rect 2308 28775 2314 28809
rect 2348 28775 2386 28809
rect 2420 28775 2426 28809
rect 2308 28736 2426 28775
rect 2308 28702 2314 28736
rect 2348 28702 2386 28736
rect 2420 28702 2426 28736
rect 2308 28663 2426 28702
rect 2308 28629 2314 28663
rect 2348 28629 2386 28663
rect 2420 28629 2426 28663
rect 2308 28590 2426 28629
rect 2308 28556 2314 28590
rect 2348 28556 2386 28590
rect 2420 28556 2426 28590
rect 2308 28517 2426 28556
rect 2308 28483 2314 28517
rect 2348 28483 2386 28517
rect 2420 28483 2426 28517
rect 2308 28444 2426 28483
rect 2308 28410 2314 28444
rect 2348 28410 2386 28444
rect 2420 28410 2426 28444
rect 2308 28371 2426 28410
rect 2308 28337 2314 28371
rect 2348 28337 2386 28371
rect 2420 28337 2426 28371
rect 2308 28298 2426 28337
rect 2308 28264 2314 28298
rect 2348 28264 2386 28298
rect 2420 28264 2426 28298
rect 2308 28225 2426 28264
rect 2308 28191 2314 28225
rect 2348 28191 2386 28225
rect 2420 28191 2426 28225
rect 2308 28152 2426 28191
rect 2308 28118 2314 28152
rect 2348 28118 2386 28152
rect 2420 28118 2426 28152
rect 2308 28079 2426 28118
rect 2308 28045 2314 28079
rect 2348 28045 2386 28079
rect 2420 28045 2426 28079
rect 2308 28006 2426 28045
rect 2308 27972 2314 28006
rect 2348 27972 2386 28006
rect 2420 27972 2426 28006
rect 2308 27933 2426 27972
rect 2308 27899 2314 27933
rect 2348 27899 2386 27933
rect 2420 27899 2426 27933
rect 2308 27860 2426 27899
rect 2871 31768 3061 31786
rect 2871 31716 2872 31768
rect 2924 31762 2940 31768
rect 2992 31762 3008 31768
rect 3060 31716 3061 31768
rect 2871 31704 2877 31716
rect 3055 31704 3061 31716
rect 2871 31652 2872 31704
rect 3060 31652 3061 31704
rect 2871 31639 2877 31652
rect 3055 31639 3061 31652
rect 2871 31587 2872 31639
rect 3060 31587 3061 31639
rect 2871 31574 2877 31587
rect 3055 31574 3061 31587
rect 2871 31522 2872 31574
rect 3060 31522 3061 31574
rect 2871 31509 2877 31522
rect 3055 31509 3061 31522
rect 2871 31457 2872 31509
rect 3060 31457 3061 31509
rect 2871 31444 2877 31457
rect 3055 31444 3061 31457
rect 2871 31392 2872 31444
rect 3060 31392 3061 31444
rect 2871 31379 2877 31392
rect 3055 31379 3061 31392
rect 2871 31327 2872 31379
rect 3060 31327 3061 31379
rect 2871 31314 2877 31327
rect 3055 31314 3061 31327
rect 2871 31262 2872 31314
rect 3060 31262 3061 31314
rect 2871 31249 2877 31262
rect 3055 31249 3061 31262
rect 2871 31197 2872 31249
rect 3060 31197 3061 31249
rect 2871 31184 2877 31197
rect 3055 31184 3061 31197
rect 2871 31132 2872 31184
rect 3060 31132 3061 31184
rect 2871 31119 2877 31132
rect 3055 31119 3061 31132
rect 2871 31067 2872 31119
rect 3060 31067 3061 31119
rect 2871 31054 2877 31067
rect 3055 31054 3061 31067
rect 2871 31002 2872 31054
rect 3060 31002 3061 31054
rect 2871 30989 2877 31002
rect 3055 30989 3061 31002
rect 2871 30937 2872 30989
rect 3060 30937 3061 30989
rect 2871 30924 2877 30937
rect 3055 30924 3061 30937
rect 2871 30872 2872 30924
rect 3060 30872 3061 30924
rect 2871 30859 2877 30872
rect 3055 30859 3061 30872
rect 2871 30807 2872 30859
rect 3060 30807 3061 30859
rect 2871 30794 2877 30807
rect 3055 30794 3061 30807
rect 2871 30742 2872 30794
rect 3060 30742 3061 30794
rect 2871 30729 2877 30742
rect 3055 30729 3061 30742
rect 2871 30677 2872 30729
rect 3060 30677 3061 30729
rect 2871 30664 2877 30677
rect 3055 30664 3061 30677
rect 2871 30612 2872 30664
rect 3060 30612 3061 30664
rect 2871 30599 2877 30612
rect 3055 30599 3061 30612
rect 2871 30547 2872 30599
rect 3060 30547 3061 30599
rect 2871 30534 2877 30547
rect 3055 30534 3061 30547
rect 2871 30482 2872 30534
rect 3060 30482 3061 30534
rect 2871 30469 2877 30482
rect 3055 30469 3061 30482
rect 2871 30417 2872 30469
rect 3060 30417 3061 30469
rect 2871 30404 2877 30417
rect 3055 30404 3061 30417
rect 2871 30352 2872 30404
rect 3060 30352 3061 30404
rect 2871 30339 2877 30352
rect 3055 30339 3061 30352
rect 2871 30287 2872 30339
rect 3060 30287 3061 30339
rect 2871 30274 2877 30287
rect 3055 30274 3061 30287
rect 2871 30222 2872 30274
rect 3060 30222 3061 30274
rect 2871 30209 2877 30222
rect 3055 30209 3061 30222
rect 2871 30157 2872 30209
rect 3060 30157 3061 30209
rect 2871 30144 2877 30157
rect 3055 30144 3061 30157
rect 2871 30092 2872 30144
rect 3060 30092 3061 30144
rect 2871 30079 2877 30092
rect 3055 30079 3061 30092
rect 2871 30027 2872 30079
rect 3060 30027 3061 30079
rect 2871 30014 2877 30027
rect 3055 30014 3061 30027
rect 2871 29962 2872 30014
rect 3060 29962 3061 30014
rect 2871 28560 2877 29962
rect 3055 28560 3061 29962
rect 2871 28521 3061 28560
rect 2871 28487 2877 28521
rect 2911 28487 2949 28521
rect 2983 28487 3021 28521
rect 3055 28487 3061 28521
rect 2871 28448 3061 28487
rect 2871 28414 2877 28448
rect 2911 28414 2949 28448
rect 2983 28414 3021 28448
rect 3055 28414 3061 28448
rect 2871 28375 3061 28414
rect 2871 28341 2877 28375
rect 2911 28341 2949 28375
rect 2983 28341 3021 28375
rect 3055 28341 3061 28375
rect 2871 28302 3061 28341
rect 2871 28268 2877 28302
rect 2911 28268 2949 28302
rect 2983 28268 3021 28302
rect 3055 28268 3061 28302
rect 2871 28229 3061 28268
rect 2871 28195 2877 28229
rect 2911 28195 2949 28229
rect 2983 28195 3021 28229
rect 3055 28195 3061 28229
rect 2871 28156 3061 28195
rect 2871 28122 2877 28156
rect 2911 28122 2949 28156
rect 2983 28122 3021 28156
rect 3055 28122 3061 28156
rect 2871 28083 3061 28122
rect 2871 28049 2877 28083
rect 2911 28049 2949 28083
rect 2983 28049 3021 28083
rect 3055 28049 3061 28083
rect 2871 28010 3061 28049
rect 2871 27976 2877 28010
rect 2911 27976 2949 28010
rect 2983 27976 3021 28010
rect 3055 27976 3061 28010
rect 2871 27937 3061 27976
rect 2871 27903 2877 27937
rect 2911 27903 2949 27937
rect 2983 27903 3021 27937
rect 3055 27903 3061 27937
rect 2871 27891 3061 27903
rect 3361 29336 3491 32497
rect 3413 29284 3439 29336
rect 3361 29270 3491 29284
rect 3413 29218 3439 29270
rect 3361 29204 3491 29218
rect 3413 29152 3439 29204
rect 3361 29138 3491 29152
rect 3413 29086 3439 29138
rect 3361 29072 3491 29086
rect 3413 29020 3439 29072
rect 3361 29006 3491 29020
rect 3413 28954 3439 29006
rect 3361 28940 3491 28954
rect 3413 28888 3439 28940
rect 3361 28874 3491 28888
rect 3413 28822 3439 28874
rect 3361 28808 3491 28822
rect 3413 28756 3439 28808
rect 3361 28742 3491 28756
rect 3413 28690 3439 28742
rect 3361 28676 3491 28690
rect 3413 28624 3439 28676
rect 3361 28610 3491 28624
rect 3413 28558 3439 28610
rect 3361 28544 3491 28558
rect 3413 28492 3439 28544
rect 3361 28478 3491 28492
rect 3413 28426 3439 28478
rect 3361 28412 3491 28426
rect 3413 28360 3439 28412
rect 3361 28346 3491 28360
rect 3413 28294 3439 28346
rect 3361 28280 3491 28294
rect 3413 28228 3439 28280
rect 3361 28214 3491 28228
rect 3413 28162 3439 28214
rect 3361 28148 3491 28162
rect 3413 28096 3439 28148
rect 3361 28082 3491 28096
rect 3413 28030 3439 28082
rect 3361 28016 3491 28030
rect 3413 27964 3439 28016
rect 3361 27949 3491 27964
rect 3413 27897 3439 27949
rect 3361 27891 3491 27897
rect 3791 37541 3797 38118
rect 3975 37541 3981 38118
rect 4711 39009 4901 39018
rect 4711 38957 4712 39009
rect 4764 38957 4780 39009
rect 4832 38957 4848 39009
rect 4900 38957 4901 39009
rect 4711 38944 4901 38957
rect 4711 38892 4712 38944
rect 4764 38892 4780 38944
rect 4832 38892 4848 38944
rect 4900 38892 4901 38944
rect 4711 38879 4901 38892
rect 4711 38827 4712 38879
rect 4764 38827 4780 38879
rect 4832 38827 4848 38879
rect 4900 38827 4901 38879
rect 4711 38824 4717 38827
rect 4751 38824 4789 38827
rect 4823 38824 4861 38827
rect 4895 38824 4901 38827
rect 4711 38814 4901 38824
rect 4711 38762 4712 38814
rect 4764 38762 4780 38814
rect 4832 38762 4848 38814
rect 4900 38762 4901 38814
rect 4711 38750 4717 38762
rect 4751 38750 4789 38762
rect 4823 38750 4861 38762
rect 4895 38750 4901 38762
rect 4711 38749 4901 38750
rect 4711 38697 4712 38749
rect 4764 38697 4780 38749
rect 4832 38697 4848 38749
rect 4900 38697 4901 38749
rect 4711 38684 4717 38697
rect 4751 38684 4789 38697
rect 4823 38684 4861 38697
rect 4895 38684 4901 38697
rect 4711 38632 4712 38684
rect 4764 38632 4780 38684
rect 4832 38632 4848 38684
rect 4900 38632 4901 38684
rect 4711 38619 4717 38632
rect 4751 38619 4789 38632
rect 4823 38619 4861 38632
rect 4895 38619 4901 38632
rect 4711 38567 4712 38619
rect 4764 38567 4780 38619
rect 4832 38567 4848 38619
rect 4900 38567 4901 38619
rect 4711 38562 4901 38567
rect 4711 38554 4717 38562
rect 4751 38554 4789 38562
rect 4823 38554 4861 38562
rect 4895 38554 4901 38562
rect 4711 38502 4712 38554
rect 4764 38502 4780 38554
rect 4832 38502 4848 38554
rect 4900 38502 4901 38554
rect 4711 38490 4901 38502
rect 4711 38438 4712 38490
rect 4764 38438 4780 38490
rect 4832 38438 4848 38490
rect 4900 38438 4901 38490
rect 4711 38426 4901 38438
rect 4711 38374 4712 38426
rect 4764 38374 4780 38426
rect 4832 38374 4848 38426
rect 4900 38374 4901 38426
rect 4711 38362 4901 38374
rect 4711 38310 4712 38362
rect 4764 38310 4780 38362
rect 4832 38310 4848 38362
rect 4900 38310 4901 38362
rect 4711 38303 4717 38310
rect 4751 38303 4789 38310
rect 4823 38303 4861 38310
rect 4895 38303 4901 38310
rect 4711 38298 4901 38303
rect 4711 38246 4712 38298
rect 4764 38246 4780 38298
rect 4832 38246 4848 38298
rect 4900 38246 4901 38298
rect 4711 38234 4717 38246
rect 4751 38234 4789 38246
rect 4823 38234 4861 38246
rect 4895 38234 4901 38246
rect 4711 38182 4712 38234
rect 4764 38182 4780 38234
rect 4832 38182 4848 38234
rect 4900 38182 4901 38234
rect 4711 38170 4717 38182
rect 4751 38170 4789 38182
rect 4823 38170 4861 38182
rect 4895 38170 4901 38182
rect 4711 38118 4712 38170
rect 4764 38118 4780 38170
rect 4832 38118 4848 38170
rect 4900 38118 4901 38170
rect 4711 38112 4901 38118
rect 4711 38078 4717 38112
rect 4751 38078 4789 38112
rect 4823 38078 4861 38112
rect 4895 38078 4901 38112
rect 4711 38037 4901 38078
rect 4711 38003 4717 38037
rect 4751 38003 4789 38037
rect 4823 38003 4861 38037
rect 4895 38003 4901 38037
rect 5631 39009 5821 39018
rect 5631 38957 5632 39009
rect 5684 38957 5700 39009
rect 5752 38957 5768 39009
rect 5820 38957 5821 39009
rect 5631 38944 5821 38957
rect 5631 38892 5632 38944
rect 5684 38892 5700 38944
rect 5752 38892 5768 38944
rect 5820 38892 5821 38944
rect 5631 38879 5821 38892
rect 5631 38827 5632 38879
rect 5684 38827 5700 38879
rect 5752 38827 5768 38879
rect 5820 38827 5821 38879
rect 5631 38824 5637 38827
rect 5671 38824 5709 38827
rect 5743 38824 5781 38827
rect 5815 38824 5821 38827
rect 5631 38814 5821 38824
rect 5631 38762 5632 38814
rect 5684 38762 5700 38814
rect 5752 38762 5768 38814
rect 5820 38762 5821 38814
rect 5631 38750 5637 38762
rect 5671 38750 5709 38762
rect 5743 38750 5781 38762
rect 5815 38750 5821 38762
rect 5631 38749 5821 38750
rect 5631 38697 5632 38749
rect 5684 38697 5700 38749
rect 5752 38697 5768 38749
rect 5820 38697 5821 38749
rect 5631 38684 5637 38697
rect 5671 38684 5709 38697
rect 5743 38684 5781 38697
rect 5815 38684 5821 38697
rect 5631 38632 5632 38684
rect 5684 38632 5700 38684
rect 5752 38632 5768 38684
rect 5820 38632 5821 38684
rect 5631 38619 5637 38632
rect 5671 38619 5709 38632
rect 5743 38619 5781 38632
rect 5815 38619 5821 38632
rect 5631 38567 5632 38619
rect 5684 38567 5700 38619
rect 5752 38567 5768 38619
rect 5820 38567 5821 38619
rect 5631 38562 5821 38567
rect 5631 38554 5637 38562
rect 5671 38554 5709 38562
rect 5743 38554 5781 38562
rect 5815 38554 5821 38562
rect 5631 38502 5632 38554
rect 5684 38502 5700 38554
rect 5752 38502 5768 38554
rect 5820 38502 5821 38554
rect 5631 38490 5821 38502
rect 5631 38438 5632 38490
rect 5684 38438 5700 38490
rect 5752 38438 5768 38490
rect 5820 38438 5821 38490
rect 5631 38426 5821 38438
rect 5631 38374 5632 38426
rect 5684 38374 5700 38426
rect 5752 38374 5768 38426
rect 5820 38374 5821 38426
rect 5631 38362 5821 38374
rect 5631 38310 5632 38362
rect 5684 38310 5700 38362
rect 5752 38310 5768 38362
rect 5820 38310 5821 38362
rect 5631 38303 5637 38310
rect 5671 38303 5709 38310
rect 5743 38303 5781 38310
rect 5815 38303 5821 38310
rect 5631 38298 5821 38303
rect 5631 38246 5632 38298
rect 5684 38246 5700 38298
rect 5752 38246 5768 38298
rect 5820 38246 5821 38298
rect 5631 38234 5637 38246
rect 5671 38234 5709 38246
rect 5743 38234 5781 38246
rect 5815 38234 5821 38246
rect 5631 38182 5632 38234
rect 5684 38182 5700 38234
rect 5752 38182 5768 38234
rect 5820 38182 5821 38234
rect 5631 38170 5637 38182
rect 5671 38170 5709 38182
rect 5743 38170 5781 38182
rect 5815 38170 5821 38182
rect 5631 38118 5632 38170
rect 5684 38118 5700 38170
rect 5752 38118 5768 38170
rect 5820 38118 5821 38170
rect 5631 38112 5821 38118
rect 5631 38078 5637 38112
rect 5671 38078 5709 38112
rect 5743 38078 5781 38112
rect 5815 38078 5821 38112
rect 5631 38037 5821 38078
rect 5631 38003 5637 38037
rect 5671 38003 5709 38037
rect 5743 38003 5781 38037
rect 5815 38003 5821 38037
rect 6551 39009 6741 39018
rect 6551 38957 6552 39009
rect 6604 38957 6620 39009
rect 6672 38957 6688 39009
rect 6740 38957 6741 39009
rect 6551 38944 6741 38957
rect 6551 38892 6552 38944
rect 6604 38892 6620 38944
rect 6672 38892 6688 38944
rect 6740 38892 6741 38944
rect 6551 38879 6741 38892
rect 6551 38827 6552 38879
rect 6604 38827 6620 38879
rect 6672 38827 6688 38879
rect 6740 38827 6741 38879
rect 6551 38824 6557 38827
rect 6591 38824 6629 38827
rect 6663 38824 6701 38827
rect 6735 38824 6741 38827
rect 6551 38814 6741 38824
rect 6551 38762 6552 38814
rect 6604 38762 6620 38814
rect 6672 38762 6688 38814
rect 6740 38762 6741 38814
rect 6551 38750 6557 38762
rect 6591 38750 6629 38762
rect 6663 38750 6701 38762
rect 6735 38750 6741 38762
rect 6551 38749 6741 38750
rect 6551 38697 6552 38749
rect 6604 38697 6620 38749
rect 6672 38697 6688 38749
rect 6740 38697 6741 38749
rect 6551 38684 6557 38697
rect 6591 38684 6629 38697
rect 6663 38684 6701 38697
rect 6735 38684 6741 38697
rect 6551 38632 6552 38684
rect 6604 38632 6620 38684
rect 6672 38632 6688 38684
rect 6740 38632 6741 38684
rect 6551 38619 6557 38632
rect 6591 38619 6629 38632
rect 6663 38619 6701 38632
rect 6735 38619 6741 38632
rect 6551 38567 6552 38619
rect 6604 38567 6620 38619
rect 6672 38567 6688 38619
rect 6740 38567 6741 38619
rect 6551 38562 6741 38567
rect 6551 38554 6557 38562
rect 6591 38554 6629 38562
rect 6663 38554 6701 38562
rect 6735 38554 6741 38562
rect 6551 38502 6552 38554
rect 6604 38502 6620 38554
rect 6672 38502 6688 38554
rect 6740 38502 6741 38554
rect 6551 38490 6741 38502
rect 6551 38438 6552 38490
rect 6604 38438 6620 38490
rect 6672 38438 6688 38490
rect 6740 38438 6741 38490
rect 6551 38426 6741 38438
rect 6551 38374 6552 38426
rect 6604 38374 6620 38426
rect 6672 38374 6688 38426
rect 6740 38374 6741 38426
rect 6551 38362 6741 38374
rect 6551 38310 6552 38362
rect 6604 38310 6620 38362
rect 6672 38310 6688 38362
rect 6740 38310 6741 38362
rect 6551 38303 6557 38310
rect 6591 38303 6629 38310
rect 6663 38303 6701 38310
rect 6735 38303 6741 38310
rect 6551 38298 6741 38303
rect 6551 38246 6552 38298
rect 6604 38246 6620 38298
rect 6672 38246 6688 38298
rect 6740 38246 6741 38298
rect 6551 38234 6557 38246
rect 6591 38234 6629 38246
rect 6663 38234 6701 38246
rect 6735 38234 6741 38246
rect 6551 38182 6552 38234
rect 6604 38182 6620 38234
rect 6672 38182 6688 38234
rect 6740 38182 6741 38234
rect 6551 38170 6557 38182
rect 6591 38170 6629 38182
rect 6663 38170 6701 38182
rect 6735 38170 6741 38182
rect 6551 38118 6552 38170
rect 6604 38118 6620 38170
rect 6672 38118 6688 38170
rect 6740 38118 6741 38170
rect 6551 38112 6741 38118
rect 6551 38078 6557 38112
rect 6591 38078 6629 38112
rect 6663 38078 6701 38112
rect 6735 38078 6741 38112
rect 6551 38037 6741 38078
rect 6551 38003 6557 38037
rect 6591 38003 6629 38037
rect 6663 38003 6701 38037
rect 6735 38003 6741 38037
rect 7471 39009 7661 39018
rect 7471 38957 7472 39009
rect 7524 38957 7540 39009
rect 7592 38957 7608 39009
rect 7660 38957 7661 39009
rect 7471 38944 7661 38957
rect 7471 38892 7472 38944
rect 7524 38892 7540 38944
rect 7592 38892 7608 38944
rect 7660 38892 7661 38944
rect 7471 38879 7661 38892
rect 7471 38827 7472 38879
rect 7524 38827 7540 38879
rect 7592 38827 7608 38879
rect 7660 38827 7661 38879
rect 7471 38824 7477 38827
rect 7511 38824 7549 38827
rect 7583 38824 7621 38827
rect 7655 38824 7661 38827
rect 7471 38814 7661 38824
rect 7471 38762 7472 38814
rect 7524 38762 7540 38814
rect 7592 38762 7608 38814
rect 7660 38762 7661 38814
rect 7471 38750 7477 38762
rect 7511 38750 7549 38762
rect 7583 38750 7621 38762
rect 7655 38750 7661 38762
rect 7471 38749 7661 38750
rect 7471 38697 7472 38749
rect 7524 38697 7540 38749
rect 7592 38697 7608 38749
rect 7660 38697 7661 38749
rect 7471 38684 7477 38697
rect 7511 38684 7549 38697
rect 7583 38684 7621 38697
rect 7655 38684 7661 38697
rect 7471 38632 7472 38684
rect 7524 38632 7540 38684
rect 7592 38632 7608 38684
rect 7660 38632 7661 38684
rect 7471 38619 7477 38632
rect 7511 38619 7549 38632
rect 7583 38619 7621 38632
rect 7655 38619 7661 38632
rect 7471 38567 7472 38619
rect 7524 38567 7540 38619
rect 7592 38567 7608 38619
rect 7660 38567 7661 38619
rect 7471 38562 7661 38567
rect 7471 38554 7477 38562
rect 7511 38554 7549 38562
rect 7583 38554 7621 38562
rect 7655 38554 7661 38562
rect 7471 38502 7472 38554
rect 7524 38502 7540 38554
rect 7592 38502 7608 38554
rect 7660 38502 7661 38554
rect 7471 38490 7661 38502
rect 7471 38438 7472 38490
rect 7524 38438 7540 38490
rect 7592 38438 7608 38490
rect 7660 38438 7661 38490
rect 7471 38426 7661 38438
rect 7471 38374 7472 38426
rect 7524 38374 7540 38426
rect 7592 38374 7608 38426
rect 7660 38374 7661 38426
rect 7471 38362 7661 38374
rect 7471 38310 7472 38362
rect 7524 38310 7540 38362
rect 7592 38310 7608 38362
rect 7660 38310 7661 38362
rect 7471 38303 7477 38310
rect 7511 38303 7549 38310
rect 7583 38303 7621 38310
rect 7655 38303 7661 38310
rect 7471 38298 7661 38303
rect 7471 38246 7472 38298
rect 7524 38246 7540 38298
rect 7592 38246 7608 38298
rect 7660 38246 7661 38298
rect 7471 38234 7477 38246
rect 7511 38234 7549 38246
rect 7583 38234 7621 38246
rect 7655 38234 7661 38246
rect 7471 38182 7472 38234
rect 7524 38182 7540 38234
rect 7592 38182 7608 38234
rect 7660 38182 7661 38234
rect 7471 38170 7477 38182
rect 7511 38170 7549 38182
rect 7583 38170 7621 38182
rect 7655 38170 7661 38182
rect 7471 38118 7472 38170
rect 7524 38118 7540 38170
rect 7592 38118 7608 38170
rect 7660 38118 7661 38170
rect 7471 38112 7661 38118
rect 7471 38078 7477 38112
rect 7511 38078 7549 38112
rect 7583 38078 7621 38112
rect 7655 38078 7661 38112
rect 7471 38037 7661 38078
rect 7471 38003 7477 38037
rect 7511 38003 7549 38037
rect 7583 38003 7621 38037
rect 7655 38003 7661 38037
rect 8391 39009 8581 39018
rect 8391 38957 8392 39009
rect 8444 38957 8460 39009
rect 8512 38957 8528 39009
rect 8580 38957 8581 39009
rect 8391 38944 8581 38957
rect 8391 38892 8392 38944
rect 8444 38892 8460 38944
rect 8512 38892 8528 38944
rect 8580 38892 8581 38944
rect 8391 38879 8581 38892
rect 8391 38827 8392 38879
rect 8444 38827 8460 38879
rect 8512 38827 8528 38879
rect 8580 38827 8581 38879
rect 8391 38824 8397 38827
rect 8431 38824 8469 38827
rect 8503 38824 8541 38827
rect 8575 38824 8581 38827
rect 8391 38814 8581 38824
rect 8391 38762 8392 38814
rect 8444 38762 8460 38814
rect 8512 38762 8528 38814
rect 8580 38762 8581 38814
rect 8391 38750 8397 38762
rect 8431 38750 8469 38762
rect 8503 38750 8541 38762
rect 8575 38750 8581 38762
rect 8391 38749 8581 38750
rect 8391 38697 8392 38749
rect 8444 38697 8460 38749
rect 8512 38697 8528 38749
rect 8580 38697 8581 38749
rect 8391 38684 8397 38697
rect 8431 38684 8469 38697
rect 8503 38684 8541 38697
rect 8575 38684 8581 38697
rect 8391 38632 8392 38684
rect 8444 38632 8460 38684
rect 8512 38632 8528 38684
rect 8580 38632 8581 38684
rect 8391 38619 8397 38632
rect 8431 38619 8469 38632
rect 8503 38619 8541 38632
rect 8575 38619 8581 38632
rect 8391 38567 8392 38619
rect 8444 38567 8460 38619
rect 8512 38567 8528 38619
rect 8580 38567 8581 38619
rect 8391 38562 8581 38567
rect 8391 38554 8397 38562
rect 8431 38554 8469 38562
rect 8503 38554 8541 38562
rect 8575 38554 8581 38562
rect 8391 38502 8392 38554
rect 8444 38502 8460 38554
rect 8512 38502 8528 38554
rect 8580 38502 8581 38554
rect 8391 38490 8581 38502
rect 8391 38438 8392 38490
rect 8444 38438 8460 38490
rect 8512 38438 8528 38490
rect 8580 38438 8581 38490
rect 8391 38426 8581 38438
rect 8391 38374 8392 38426
rect 8444 38374 8460 38426
rect 8512 38374 8528 38426
rect 8580 38374 8581 38426
rect 8391 38362 8581 38374
rect 8391 38310 8392 38362
rect 8444 38310 8460 38362
rect 8512 38310 8528 38362
rect 8580 38310 8581 38362
rect 8391 38303 8397 38310
rect 8431 38303 8469 38310
rect 8503 38303 8541 38310
rect 8575 38303 8581 38310
rect 8391 38298 8581 38303
rect 8391 38246 8392 38298
rect 8444 38246 8460 38298
rect 8512 38246 8528 38298
rect 8580 38246 8581 38298
rect 8391 38234 8397 38246
rect 8431 38234 8469 38246
rect 8503 38234 8541 38246
rect 8575 38234 8581 38246
rect 8391 38182 8392 38234
rect 8444 38182 8460 38234
rect 8512 38182 8528 38234
rect 8580 38182 8581 38234
rect 8391 38170 8397 38182
rect 8431 38170 8469 38182
rect 8503 38170 8541 38182
rect 8575 38170 8581 38182
rect 8391 38118 8392 38170
rect 8444 38118 8460 38170
rect 8512 38118 8528 38170
rect 8580 38118 8581 38170
rect 8391 38112 8581 38118
rect 8391 38078 8397 38112
rect 8431 38078 8469 38112
rect 8503 38078 8541 38112
rect 8575 38078 8581 38112
rect 8391 38037 8581 38078
rect 8391 38003 8397 38037
rect 8431 38003 8469 38037
rect 8503 38003 8541 38037
rect 8575 38003 8581 38037
rect 9311 39009 9501 39018
rect 9311 38957 9312 39009
rect 9364 38957 9380 39009
rect 9432 38957 9448 39009
rect 9500 38957 9501 39009
rect 9311 38944 9501 38957
rect 9311 38892 9312 38944
rect 9364 38892 9380 38944
rect 9432 38892 9448 38944
rect 9500 38892 9501 38944
rect 9311 38879 9501 38892
rect 9311 38827 9312 38879
rect 9364 38827 9380 38879
rect 9432 38827 9448 38879
rect 9500 38827 9501 38879
rect 9311 38824 9317 38827
rect 9351 38824 9389 38827
rect 9423 38824 9461 38827
rect 9495 38824 9501 38827
rect 9311 38814 9501 38824
rect 9311 38762 9312 38814
rect 9364 38762 9380 38814
rect 9432 38762 9448 38814
rect 9500 38762 9501 38814
rect 9311 38750 9317 38762
rect 9351 38750 9389 38762
rect 9423 38750 9461 38762
rect 9495 38750 9501 38762
rect 9311 38749 9501 38750
rect 9311 38697 9312 38749
rect 9364 38697 9380 38749
rect 9432 38697 9448 38749
rect 9500 38697 9501 38749
rect 9311 38684 9317 38697
rect 9351 38684 9389 38697
rect 9423 38684 9461 38697
rect 9495 38684 9501 38697
rect 9311 38632 9312 38684
rect 9364 38632 9380 38684
rect 9432 38632 9448 38684
rect 9500 38632 9501 38684
rect 9311 38619 9317 38632
rect 9351 38619 9389 38632
rect 9423 38619 9461 38632
rect 9495 38619 9501 38632
rect 9311 38567 9312 38619
rect 9364 38567 9380 38619
rect 9432 38567 9448 38619
rect 9500 38567 9501 38619
rect 9311 38562 9501 38567
rect 9311 38554 9317 38562
rect 9351 38554 9389 38562
rect 9423 38554 9461 38562
rect 9495 38554 9501 38562
rect 9311 38502 9312 38554
rect 9364 38502 9380 38554
rect 9432 38502 9448 38554
rect 9500 38502 9501 38554
rect 9311 38490 9501 38502
rect 9311 38438 9312 38490
rect 9364 38438 9380 38490
rect 9432 38438 9448 38490
rect 9500 38438 9501 38490
rect 9311 38426 9501 38438
rect 9311 38374 9312 38426
rect 9364 38374 9380 38426
rect 9432 38374 9448 38426
rect 9500 38374 9501 38426
rect 9311 38362 9501 38374
rect 9311 38310 9312 38362
rect 9364 38310 9380 38362
rect 9432 38310 9448 38362
rect 9500 38310 9501 38362
rect 9311 38303 9317 38310
rect 9351 38303 9389 38310
rect 9423 38303 9461 38310
rect 9495 38303 9501 38310
rect 9311 38298 9501 38303
rect 9311 38246 9312 38298
rect 9364 38246 9380 38298
rect 9432 38246 9448 38298
rect 9500 38246 9501 38298
rect 9311 38234 9317 38246
rect 9351 38234 9389 38246
rect 9423 38234 9461 38246
rect 9495 38234 9501 38246
rect 9311 38182 9312 38234
rect 9364 38182 9380 38234
rect 9432 38182 9448 38234
rect 9500 38182 9501 38234
rect 9311 38170 9317 38182
rect 9351 38170 9389 38182
rect 9423 38170 9461 38182
rect 9495 38170 9501 38182
rect 9311 38118 9312 38170
rect 9364 38118 9380 38170
rect 9432 38118 9448 38170
rect 9500 38118 9501 38170
rect 9311 38112 9501 38118
rect 9311 38078 9317 38112
rect 9351 38078 9389 38112
rect 9423 38078 9461 38112
rect 9495 38078 9501 38112
rect 9311 38037 9501 38078
rect 9311 38003 9317 38037
rect 9351 38003 9389 38037
rect 9423 38003 9461 38037
rect 9495 38003 9501 38037
rect 10231 39009 10421 39018
rect 10231 38957 10232 39009
rect 10284 38957 10300 39009
rect 10352 38957 10368 39009
rect 10420 38957 10421 39009
rect 10231 38944 10421 38957
rect 10231 38892 10232 38944
rect 10284 38892 10300 38944
rect 10352 38892 10368 38944
rect 10420 38892 10421 38944
rect 10231 38879 10421 38892
rect 10231 38827 10232 38879
rect 10284 38827 10300 38879
rect 10352 38827 10368 38879
rect 10420 38827 10421 38879
rect 10231 38824 10237 38827
rect 10271 38824 10309 38827
rect 10343 38824 10381 38827
rect 10415 38824 10421 38827
rect 10231 38814 10421 38824
rect 10231 38762 10232 38814
rect 10284 38762 10300 38814
rect 10352 38762 10368 38814
rect 10420 38762 10421 38814
rect 10231 38750 10237 38762
rect 10271 38750 10309 38762
rect 10343 38750 10381 38762
rect 10415 38750 10421 38762
rect 10231 38749 10421 38750
rect 10231 38697 10232 38749
rect 10284 38697 10300 38749
rect 10352 38697 10368 38749
rect 10420 38697 10421 38749
rect 10231 38684 10237 38697
rect 10271 38684 10309 38697
rect 10343 38684 10381 38697
rect 10415 38684 10421 38697
rect 10231 38632 10232 38684
rect 10284 38632 10300 38684
rect 10352 38632 10368 38684
rect 10420 38632 10421 38684
rect 10231 38619 10237 38632
rect 10271 38619 10309 38632
rect 10343 38619 10381 38632
rect 10415 38619 10421 38632
rect 10231 38567 10232 38619
rect 10284 38567 10300 38619
rect 10352 38567 10368 38619
rect 10420 38567 10421 38619
rect 10231 38562 10421 38567
rect 10231 38554 10237 38562
rect 10271 38554 10309 38562
rect 10343 38554 10381 38562
rect 10415 38554 10421 38562
rect 10231 38502 10232 38554
rect 10284 38502 10300 38554
rect 10352 38502 10368 38554
rect 10420 38502 10421 38554
rect 10231 38490 10421 38502
rect 10231 38438 10232 38490
rect 10284 38438 10300 38490
rect 10352 38438 10368 38490
rect 10420 38438 10421 38490
rect 10231 38426 10421 38438
rect 10231 38374 10232 38426
rect 10284 38374 10300 38426
rect 10352 38374 10368 38426
rect 10420 38374 10421 38426
rect 10231 38362 10421 38374
rect 10231 38310 10232 38362
rect 10284 38310 10300 38362
rect 10352 38310 10368 38362
rect 10420 38310 10421 38362
rect 10231 38303 10237 38310
rect 10271 38303 10309 38310
rect 10343 38303 10381 38310
rect 10415 38303 10421 38310
rect 10231 38298 10421 38303
rect 10231 38246 10232 38298
rect 10284 38246 10300 38298
rect 10352 38246 10368 38298
rect 10420 38246 10421 38298
rect 10231 38234 10237 38246
rect 10271 38234 10309 38246
rect 10343 38234 10381 38246
rect 10415 38234 10421 38246
rect 10231 38182 10232 38234
rect 10284 38182 10300 38234
rect 10352 38182 10368 38234
rect 10420 38182 10421 38234
rect 10231 38170 10237 38182
rect 10271 38170 10309 38182
rect 10343 38170 10381 38182
rect 10415 38170 10421 38182
rect 10231 38118 10232 38170
rect 10284 38118 10300 38170
rect 10352 38118 10368 38170
rect 10420 38118 10421 38170
rect 10231 38112 10421 38118
rect 10231 38078 10237 38112
rect 10271 38078 10309 38112
rect 10343 38078 10381 38112
rect 10415 38078 10421 38112
rect 10231 38037 10421 38078
rect 10231 38003 10237 38037
rect 10271 38003 10309 38037
rect 10343 38003 10381 38037
rect 10415 38003 10421 38037
rect 11151 39009 11157 39028
rect 11335 39009 11341 39028
rect 11151 38957 11152 39009
rect 11340 38957 11341 39009
rect 11151 38944 11157 38957
rect 11335 38944 11341 38957
rect 11151 38892 11152 38944
rect 11340 38892 11341 38944
rect 11151 38879 11157 38892
rect 11335 38879 11341 38892
rect 11151 38827 11152 38879
rect 11340 38827 11341 38879
rect 11151 38814 11157 38827
rect 11335 38814 11341 38827
rect 11151 38762 11152 38814
rect 11340 38762 11341 38814
rect 11151 38749 11157 38762
rect 11335 38749 11341 38762
rect 11151 38697 11152 38749
rect 11340 38697 11341 38749
rect 11151 38684 11157 38697
rect 11335 38684 11341 38697
rect 11151 38632 11152 38684
rect 11340 38632 11341 38684
rect 11151 38619 11157 38632
rect 11335 38619 11341 38632
rect 11151 38567 11152 38619
rect 11340 38567 11341 38619
rect 11151 38554 11157 38567
rect 11335 38554 11341 38567
rect 11151 38502 11152 38554
rect 11340 38502 11341 38554
rect 11151 38490 11157 38502
rect 11335 38490 11341 38502
rect 11151 38438 11152 38490
rect 11204 38438 11220 38490
rect 11272 38438 11288 38490
rect 11340 38438 11341 38490
rect 11151 38426 11157 38438
rect 11191 38426 11229 38438
rect 11263 38426 11301 38438
rect 11335 38426 11341 38438
rect 11151 38374 11152 38426
rect 11204 38374 11220 38426
rect 11272 38374 11288 38426
rect 11340 38374 11341 38426
rect 11151 38362 11157 38374
rect 11191 38362 11229 38374
rect 11263 38362 11301 38374
rect 11335 38362 11341 38374
rect 11151 38310 11152 38362
rect 11204 38310 11220 38362
rect 11272 38310 11288 38362
rect 11340 38310 11341 38362
rect 11151 38305 11341 38310
rect 11151 38298 11157 38305
rect 11191 38298 11229 38305
rect 11263 38298 11301 38305
rect 11335 38298 11341 38305
rect 11151 38246 11152 38298
rect 11204 38246 11220 38298
rect 11272 38246 11288 38298
rect 11340 38246 11341 38298
rect 11151 38234 11341 38246
rect 11151 38182 11152 38234
rect 11204 38182 11220 38234
rect 11272 38182 11288 38234
rect 11340 38182 11341 38234
rect 11151 38170 11341 38182
rect 11151 38118 11152 38170
rect 11204 38118 11220 38170
rect 11272 38118 11288 38170
rect 11340 38118 11341 38170
rect 11151 38086 11341 38118
rect 11151 38052 11157 38086
rect 11191 38052 11229 38086
rect 11263 38052 11301 38086
rect 11335 38052 11341 38086
rect 11151 38013 11341 38052
rect 3791 37502 3981 37541
rect 3791 37468 3797 37502
rect 3831 37468 3869 37502
rect 3903 37468 3941 37502
rect 3975 37468 3981 37502
rect 3791 37429 3981 37468
rect 3791 37395 3797 37429
rect 3831 37395 3869 37429
rect 3903 37395 3941 37429
rect 3975 37395 3981 37429
rect 3791 37356 3981 37395
rect 3791 37322 3797 37356
rect 3831 37322 3869 37356
rect 3903 37322 3941 37356
rect 3975 37322 3981 37356
rect 3791 37283 3981 37322
rect 3791 37249 3797 37283
rect 3831 37249 3869 37283
rect 3903 37249 3941 37283
rect 3975 37249 3981 37283
rect 3791 37210 3981 37249
rect 3791 37176 3797 37210
rect 3831 37176 3869 37210
rect 3903 37176 3941 37210
rect 3975 37176 3981 37210
rect 3791 37137 3981 37176
rect 3791 37103 3797 37137
rect 3831 37103 3869 37137
rect 3903 37103 3941 37137
rect 3975 37103 3981 37137
rect 3791 36362 3981 37103
rect 3791 36290 3797 36362
rect 3975 36290 3981 36362
rect 3791 36238 3792 36290
rect 3980 36238 3981 36290
rect 3791 36226 3797 36238
rect 3975 36226 3981 36238
rect 3791 36174 3792 36226
rect 3980 36174 3981 36226
rect 3791 36162 3797 36174
rect 3975 36162 3981 36174
rect 3791 36110 3792 36162
rect 3980 36110 3981 36162
rect 3791 36098 3797 36110
rect 3975 36098 3981 36110
rect 3791 36046 3792 36098
rect 3980 36046 3981 36098
rect 3791 36034 3797 36046
rect 3975 36034 3981 36046
rect 3791 35982 3792 36034
rect 3980 35982 3981 36034
rect 3791 35970 3797 35982
rect 3975 35970 3981 35982
rect 3791 35918 3792 35970
rect 3980 35918 3981 35970
rect 3791 35906 3797 35918
rect 3975 35906 3981 35918
rect 3791 35854 3792 35906
rect 3980 35854 3981 35906
rect 3791 35842 3797 35854
rect 3975 35842 3981 35854
rect 3791 35790 3792 35842
rect 3980 35790 3981 35842
rect 3791 35778 3797 35790
rect 3975 35778 3981 35790
rect 3791 35726 3792 35778
rect 3980 35726 3981 35778
rect 3791 35714 3797 35726
rect 3975 35714 3981 35726
rect 3791 35662 3792 35714
rect 3980 35662 3981 35714
rect 3791 35650 3797 35662
rect 3975 35650 3981 35662
rect 3791 35598 3792 35650
rect 3980 35598 3981 35650
rect 3791 35586 3797 35598
rect 3975 35586 3981 35598
rect 3791 35534 3792 35586
rect 3980 35534 3981 35586
rect 3791 35522 3797 35534
rect 3975 35522 3981 35534
rect 3791 35470 3792 35522
rect 3980 35470 3981 35522
rect 3791 35458 3797 35470
rect 3975 35458 3981 35470
rect 3791 35406 3792 35458
rect 3980 35406 3981 35458
rect 3791 35394 3797 35406
rect 3975 35394 3981 35406
rect 3791 35342 3792 35394
rect 3980 35342 3981 35394
rect 3791 35329 3797 35342
rect 3975 35329 3981 35342
rect 3791 35277 3792 35329
rect 3980 35277 3981 35329
rect 3791 35264 3797 35277
rect 3975 35264 3981 35277
rect 3791 35212 3792 35264
rect 3980 35212 3981 35264
rect 3791 35199 3797 35212
rect 3975 35199 3981 35212
rect 3791 35147 3792 35199
rect 3980 35147 3981 35199
rect 3791 35134 3797 35147
rect 3975 35134 3981 35147
rect 3791 35082 3792 35134
rect 3980 35082 3981 35134
rect 3791 35069 3797 35082
rect 3975 35069 3981 35082
rect 3791 35017 3792 35069
rect 3980 35017 3981 35069
rect 3791 35004 3797 35017
rect 3975 35004 3981 35017
rect 3791 34952 3792 35004
rect 3980 34952 3981 35004
rect 3791 34939 3797 34952
rect 3975 34939 3981 34952
rect 3791 34887 3792 34939
rect 3980 34887 3981 34939
rect 3791 34874 3797 34887
rect 3975 34874 3981 34887
rect 3791 34822 3792 34874
rect 3980 34822 3981 34874
rect 3791 34809 3797 34822
rect 3975 34809 3981 34822
rect 3791 34757 3792 34809
rect 3980 34757 3981 34809
rect 3791 34744 3797 34757
rect 3975 34744 3981 34757
rect 3791 34692 3792 34744
rect 3980 34692 3981 34744
rect 3791 34679 3797 34692
rect 3975 34679 3981 34692
rect 3791 34627 3792 34679
rect 3980 34627 3981 34679
rect 3791 34614 3797 34627
rect 3975 34614 3981 34627
rect 3791 34562 3792 34614
rect 3980 34562 3981 34614
rect 3791 33160 3797 34562
rect 3975 33160 3981 34562
rect 3791 33121 3981 33160
rect 3791 33087 3797 33121
rect 3831 33087 3869 33121
rect 3903 33087 3941 33121
rect 3975 33087 3981 33121
rect 3791 33048 3981 33087
rect 3791 33014 3797 33048
rect 3831 33014 3869 33048
rect 3903 33014 3941 33048
rect 3975 33014 3981 33048
rect 3791 32975 3981 33014
rect 3791 32941 3797 32975
rect 3831 32941 3869 32975
rect 3903 32941 3941 32975
rect 3975 32941 3981 32975
rect 3791 32902 3981 32941
rect 3791 32868 3797 32902
rect 3831 32868 3869 32902
rect 3903 32868 3941 32902
rect 3975 32868 3981 32902
rect 3791 32829 3981 32868
rect 3791 32795 3797 32829
rect 3831 32795 3869 32829
rect 3903 32795 3941 32829
rect 3975 32795 3981 32829
rect 3791 32756 3981 32795
rect 3791 32722 3797 32756
rect 3831 32722 3869 32756
rect 3903 32722 3941 32756
rect 3975 32722 3981 32756
rect 3791 32683 3981 32722
rect 3791 32649 3797 32683
rect 3831 32649 3869 32683
rect 3903 32649 3941 32683
rect 3975 32649 3981 32683
rect 3791 32610 3981 32649
rect 3791 32576 3797 32610
rect 3831 32576 3869 32610
rect 3903 32576 3941 32610
rect 3975 32576 3981 32610
rect 3791 32537 3981 32576
rect 3791 32503 3797 32537
rect 3831 32503 3869 32537
rect 3903 32503 3941 32537
rect 3975 32503 3981 32537
rect 3791 31762 3981 32503
rect 3791 31690 3797 31762
rect 3975 31690 3981 31762
rect 3791 31638 3792 31690
rect 3980 31638 3981 31690
rect 3791 31626 3797 31638
rect 3975 31626 3981 31638
rect 3791 31574 3792 31626
rect 3980 31574 3981 31626
rect 3791 31562 3797 31574
rect 3975 31562 3981 31574
rect 3791 31510 3792 31562
rect 3980 31510 3981 31562
rect 3791 31498 3797 31510
rect 3975 31498 3981 31510
rect 3791 31446 3792 31498
rect 3980 31446 3981 31498
rect 3791 31434 3797 31446
rect 3975 31434 3981 31446
rect 3791 31382 3792 31434
rect 3980 31382 3981 31434
rect 3791 31370 3797 31382
rect 3975 31370 3981 31382
rect 3791 31318 3792 31370
rect 3980 31318 3981 31370
rect 3791 31306 3797 31318
rect 3975 31306 3981 31318
rect 3791 31254 3792 31306
rect 3980 31254 3981 31306
rect 3791 31242 3797 31254
rect 3975 31242 3981 31254
rect 3791 31190 3792 31242
rect 3980 31190 3981 31242
rect 3791 31178 3797 31190
rect 3975 31178 3981 31190
rect 3791 31126 3792 31178
rect 3980 31126 3981 31178
rect 3791 31114 3797 31126
rect 3975 31114 3981 31126
rect 3791 31062 3792 31114
rect 3980 31062 3981 31114
rect 3791 31050 3797 31062
rect 3975 31050 3981 31062
rect 3791 30998 3792 31050
rect 3980 30998 3981 31050
rect 3791 30986 3797 30998
rect 3975 30986 3981 30998
rect 3791 30934 3792 30986
rect 3980 30934 3981 30986
rect 3791 30922 3797 30934
rect 3975 30922 3981 30934
rect 3791 30870 3792 30922
rect 3980 30870 3981 30922
rect 3791 30858 3797 30870
rect 3975 30858 3981 30870
rect 3791 30806 3792 30858
rect 3980 30806 3981 30858
rect 3791 30794 3797 30806
rect 3975 30794 3981 30806
rect 3791 30742 3792 30794
rect 3980 30742 3981 30794
rect 3791 30729 3797 30742
rect 3975 30729 3981 30742
rect 3791 30677 3792 30729
rect 3980 30677 3981 30729
rect 3791 30664 3797 30677
rect 3975 30664 3981 30677
rect 3791 30612 3792 30664
rect 3980 30612 3981 30664
rect 3791 30599 3797 30612
rect 3975 30599 3981 30612
rect 3791 30547 3792 30599
rect 3980 30547 3981 30599
rect 3791 30534 3797 30547
rect 3975 30534 3981 30547
rect 3791 30482 3792 30534
rect 3980 30482 3981 30534
rect 3791 30469 3797 30482
rect 3975 30469 3981 30482
rect 3791 30417 3792 30469
rect 3980 30417 3981 30469
rect 3791 30404 3797 30417
rect 3975 30404 3981 30417
rect 3791 30352 3792 30404
rect 3980 30352 3981 30404
rect 3791 30339 3797 30352
rect 3975 30339 3981 30352
rect 3791 30287 3792 30339
rect 3980 30287 3981 30339
rect 3791 30274 3797 30287
rect 3975 30274 3981 30287
rect 3791 30222 3792 30274
rect 3980 30222 3981 30274
rect 3791 30209 3797 30222
rect 3975 30209 3981 30222
rect 3791 30157 3792 30209
rect 3980 30157 3981 30209
rect 3791 30144 3797 30157
rect 3975 30144 3981 30157
rect 3791 30092 3792 30144
rect 3980 30092 3981 30144
rect 3791 30079 3797 30092
rect 3975 30079 3981 30092
rect 3791 30027 3792 30079
rect 3980 30027 3981 30079
rect 3791 30014 3797 30027
rect 3975 30014 3981 30027
rect 3791 29962 3792 30014
rect 3980 29962 3981 30014
rect 3791 28560 3797 29962
rect 3975 28560 3981 29962
rect 3791 28521 3981 28560
rect 3791 28487 3797 28521
rect 3831 28487 3869 28521
rect 3903 28487 3941 28521
rect 3975 28487 3981 28521
rect 3791 28448 3981 28487
rect 3791 28414 3797 28448
rect 3831 28414 3869 28448
rect 3903 28414 3941 28448
rect 3975 28414 3981 28448
rect 3791 28375 3981 28414
rect 3791 28341 3797 28375
rect 3831 28341 3869 28375
rect 3903 28341 3941 28375
rect 3975 28341 3981 28375
rect 3791 28302 3981 28341
rect 3791 28268 3797 28302
rect 3831 28268 3869 28302
rect 3903 28268 3941 28302
rect 3975 28268 3981 28302
rect 3791 28229 3981 28268
rect 3791 28195 3797 28229
rect 3831 28195 3869 28229
rect 3903 28195 3941 28229
rect 3975 28195 3981 28229
rect 3791 28156 3981 28195
rect 3791 28122 3797 28156
rect 3831 28122 3869 28156
rect 3903 28122 3941 28156
rect 3975 28122 3981 28156
rect 3791 28083 3981 28122
rect 3791 28049 3797 28083
rect 3831 28049 3869 28083
rect 3903 28049 3941 28083
rect 3975 28049 3981 28083
rect 3791 28010 3981 28049
rect 3791 27976 3797 28010
rect 3831 27976 3869 28010
rect 3903 27976 3941 28010
rect 3975 27976 3981 28010
rect 3791 27937 3981 27976
rect 3791 27903 3797 27937
rect 3831 27903 3869 27937
rect 3903 27903 3941 27937
rect 3975 27903 3981 27937
rect 3791 27891 3981 27903
rect 4281 37997 4411 38003
rect 4333 37945 4359 37997
rect 4281 37929 4411 37945
rect 4333 37877 4359 37929
rect 4281 37861 4411 37877
rect 4333 37809 4359 37861
rect 4281 37793 4411 37809
rect 4333 37741 4359 37793
rect 4281 37725 4411 37741
rect 4333 37673 4359 37725
rect 4281 37657 4411 37673
rect 4333 37605 4359 37657
rect 4281 37589 4411 37605
rect 4333 37537 4359 37589
rect 4281 37521 4411 37537
rect 4333 37469 4359 37521
rect 4281 37453 4411 37469
rect 4333 37401 4359 37453
rect 4281 37385 4411 37401
rect 4333 37333 4359 37385
rect 4281 37318 4411 37333
rect 4333 37266 4359 37318
rect 4281 37251 4411 37266
rect 4333 37199 4359 37251
rect 4281 37184 4411 37199
rect 4333 37132 4359 37184
rect 4281 37117 4411 37132
rect 4333 37065 4359 37117
rect 4281 34225 4411 37065
rect 4333 34173 4359 34225
rect 4281 34161 4411 34173
rect 4333 34109 4359 34161
rect 4281 34097 4411 34109
rect 4333 34045 4359 34097
rect 4281 34033 4411 34045
rect 4333 33981 4359 34033
rect 4281 33969 4411 33981
rect 4333 33917 4359 33969
rect 4281 33905 4411 33917
rect 4333 33853 4359 33905
rect 4281 33841 4411 33853
rect 4333 33789 4359 33841
rect 4281 33777 4411 33789
rect 4333 33725 4359 33777
rect 4281 33713 4411 33725
rect 4333 33661 4359 33713
rect 4281 33649 4411 33661
rect 4333 33597 4359 33649
rect 4281 33585 4411 33597
rect 4333 33533 4359 33585
rect 4281 33521 4411 33533
rect 4333 33469 4359 33521
rect 4281 33457 4411 33469
rect 4333 33405 4359 33457
rect 4281 33393 4411 33405
rect 4333 33341 4359 33393
rect 4281 33329 4411 33341
rect 4333 33277 4359 33329
rect 4281 33264 4411 33277
rect 4333 33212 4359 33264
rect 4281 33199 4411 33212
rect 4333 33147 4359 33199
rect 4281 33134 4411 33147
rect 4333 33082 4359 33134
rect 4281 33069 4411 33082
rect 4333 33017 4359 33069
rect 4281 33004 4411 33017
rect 4333 32952 4359 33004
rect 4281 32939 4411 32952
rect 4333 32887 4359 32939
rect 4281 32874 4411 32887
rect 4333 32822 4359 32874
rect 4281 32809 4411 32822
rect 4333 32757 4359 32809
rect 4281 32744 4411 32757
rect 4333 32692 4359 32744
rect 4281 32679 4411 32692
rect 4333 32627 4359 32679
rect 4281 32614 4411 32627
rect 4333 32562 4359 32614
rect 4281 32549 4411 32562
rect 4333 32497 4359 32549
rect 4281 29625 4411 32497
rect 4333 29573 4359 29625
rect 4281 29561 4411 29573
rect 4333 29509 4359 29561
rect 4281 29497 4411 29509
rect 4333 29445 4359 29497
rect 4281 29433 4411 29445
rect 4333 29381 4359 29433
rect 4281 29369 4411 29381
rect 4333 29317 4359 29369
rect 4281 29305 4411 29317
rect 4333 29253 4359 29305
rect 4281 29241 4411 29253
rect 4333 29189 4359 29241
rect 4281 29177 4411 29189
rect 4333 29125 4359 29177
rect 4281 29113 4411 29125
rect 4333 29061 4359 29113
rect 4281 29049 4411 29061
rect 4333 28997 4359 29049
rect 4281 28985 4411 28997
rect 4333 28933 4359 28985
rect 4281 28921 4411 28933
rect 4333 28869 4359 28921
rect 4281 28857 4411 28869
rect 4333 28805 4359 28857
rect 4281 28793 4411 28805
rect 4333 28741 4359 28793
rect 4281 28729 4411 28741
rect 4333 28677 4359 28729
rect 4281 28664 4411 28677
rect 4333 28612 4359 28664
rect 4281 28599 4411 28612
rect 4333 28547 4359 28599
rect 4281 28534 4411 28547
rect 4333 28482 4359 28534
rect 4281 28469 4411 28482
rect 4333 28417 4359 28469
rect 4281 28404 4411 28417
rect 4333 28352 4359 28404
rect 4281 28339 4411 28352
rect 4333 28287 4359 28339
rect 4281 28274 4411 28287
rect 4333 28222 4359 28274
rect 4281 28209 4411 28222
rect 4333 28157 4359 28209
rect 4281 28144 4411 28157
rect 4333 28092 4359 28144
rect 4281 28079 4411 28092
rect 4333 28027 4359 28079
rect 4281 28014 4411 28027
rect 4333 27962 4359 28014
rect 4281 27949 4411 27962
rect 4333 27897 4359 27949
rect 4281 27891 4411 27897
rect 4711 37962 4901 38003
rect 4711 37928 4717 37962
rect 4751 37928 4789 37962
rect 4823 37928 4861 37962
rect 4895 37928 4901 37962
rect 4711 37887 4901 37928
rect 4711 37853 4717 37887
rect 4751 37853 4789 37887
rect 4823 37853 4861 37887
rect 4895 37853 4901 37887
rect 4711 37812 4901 37853
rect 4711 37778 4717 37812
rect 4751 37778 4789 37812
rect 4823 37778 4861 37812
rect 4895 37778 4901 37812
rect 4711 37737 4901 37778
rect 4711 37703 4717 37737
rect 4751 37703 4789 37737
rect 4823 37703 4861 37737
rect 4895 37703 4901 37737
rect 4711 37662 4901 37703
rect 4711 37628 4717 37662
rect 4751 37628 4789 37662
rect 4823 37628 4861 37662
rect 4895 37628 4901 37662
rect 4711 37587 4901 37628
rect 4711 37553 4717 37587
rect 4751 37553 4789 37587
rect 4823 37553 4861 37587
rect 4895 37553 4901 37587
rect 4711 37512 4901 37553
rect 4711 37478 4717 37512
rect 4751 37478 4789 37512
rect 4823 37478 4861 37512
rect 4895 37478 4901 37512
rect 4711 37437 4901 37478
rect 4711 37403 4717 37437
rect 4751 37403 4789 37437
rect 4823 37403 4861 37437
rect 4895 37403 4901 37437
rect 4711 37362 4901 37403
rect 4711 37328 4717 37362
rect 4751 37328 4789 37362
rect 4823 37328 4861 37362
rect 4895 37328 4901 37362
rect 4711 37287 4901 37328
rect 4711 37253 4717 37287
rect 4751 37253 4789 37287
rect 4823 37253 4861 37287
rect 4895 37253 4901 37287
rect 4711 37212 4901 37253
rect 4711 37178 4717 37212
rect 4751 37178 4789 37212
rect 4823 37178 4861 37212
rect 4895 37178 4901 37212
rect 4711 37137 4901 37178
rect 4711 37103 4717 37137
rect 4751 37103 4789 37137
rect 4823 37103 4861 37137
rect 4895 37103 4901 37137
rect 4711 36353 4901 37103
rect 4711 36290 4717 36353
rect 4895 36290 4901 36353
rect 4711 36238 4712 36290
rect 4900 36238 4901 36290
rect 4711 36226 4717 36238
rect 4895 36226 4901 36238
rect 4711 36174 4712 36226
rect 4900 36174 4901 36226
rect 4711 36162 4717 36174
rect 4895 36162 4901 36174
rect 4711 36110 4712 36162
rect 4900 36110 4901 36162
rect 4711 36098 4717 36110
rect 4895 36098 4901 36110
rect 4711 36046 4712 36098
rect 4900 36046 4901 36098
rect 4711 36034 4717 36046
rect 4895 36034 4901 36046
rect 4711 35982 4712 36034
rect 4900 35982 4901 36034
rect 4711 35970 4717 35982
rect 4895 35970 4901 35982
rect 4711 35918 4712 35970
rect 4900 35918 4901 35970
rect 4711 35906 4717 35918
rect 4895 35906 4901 35918
rect 4711 35854 4712 35906
rect 4900 35854 4901 35906
rect 4711 35842 4717 35854
rect 4895 35842 4901 35854
rect 4711 35790 4712 35842
rect 4900 35790 4901 35842
rect 4711 35778 4717 35790
rect 4895 35778 4901 35790
rect 4711 35726 4712 35778
rect 4900 35726 4901 35778
rect 4711 35714 4717 35726
rect 4895 35714 4901 35726
rect 4711 35662 4712 35714
rect 4900 35662 4901 35714
rect 4711 35650 4717 35662
rect 4895 35650 4901 35662
rect 4711 35598 4712 35650
rect 4900 35598 4901 35650
rect 4711 35586 4717 35598
rect 4895 35586 4901 35598
rect 4711 35534 4712 35586
rect 4900 35534 4901 35586
rect 4711 35522 4717 35534
rect 4895 35522 4901 35534
rect 4711 35470 4712 35522
rect 4900 35470 4901 35522
rect 4711 35458 4717 35470
rect 4895 35458 4901 35470
rect 4711 35406 4712 35458
rect 4900 35406 4901 35458
rect 4711 35394 4717 35406
rect 4895 35394 4901 35406
rect 4711 35342 4712 35394
rect 4900 35342 4901 35394
rect 4711 35329 4717 35342
rect 4895 35329 4901 35342
rect 4711 35277 4712 35329
rect 4900 35277 4901 35329
rect 4711 35264 4717 35277
rect 4895 35264 4901 35277
rect 4711 35212 4712 35264
rect 4900 35212 4901 35264
rect 4711 35199 4717 35212
rect 4895 35199 4901 35212
rect 4711 35147 4712 35199
rect 4900 35147 4901 35199
rect 4711 35134 4717 35147
rect 4895 35134 4901 35147
rect 4711 35082 4712 35134
rect 4900 35082 4901 35134
rect 4711 35069 4717 35082
rect 4895 35069 4901 35082
rect 4711 35017 4712 35069
rect 4900 35017 4901 35069
rect 4711 35004 4717 35017
rect 4895 35004 4901 35017
rect 4711 34952 4712 35004
rect 4900 34952 4901 35004
rect 4711 34939 4717 34952
rect 4895 34939 4901 34952
rect 4711 34887 4712 34939
rect 4900 34887 4901 34939
rect 4711 34874 4717 34887
rect 4895 34874 4901 34887
rect 4711 34822 4712 34874
rect 4900 34822 4901 34874
rect 4711 34809 4717 34822
rect 4895 34809 4901 34822
rect 4711 34757 4712 34809
rect 4900 34757 4901 34809
rect 4711 34744 4717 34757
rect 4895 34744 4901 34757
rect 4711 34692 4712 34744
rect 4900 34692 4901 34744
rect 4711 34679 4717 34692
rect 4895 34679 4901 34692
rect 4711 34627 4712 34679
rect 4900 34627 4901 34679
rect 4711 34614 4717 34627
rect 4895 34614 4901 34627
rect 4711 34562 4712 34614
rect 4900 34562 4901 34614
rect 4711 32503 4717 34562
rect 4895 32503 4901 34562
rect 4711 31753 4901 32503
rect 4711 31690 4717 31753
rect 4895 31690 4901 31753
rect 4711 31638 4712 31690
rect 4900 31638 4901 31690
rect 4711 31626 4717 31638
rect 4895 31626 4901 31638
rect 4711 31574 4712 31626
rect 4900 31574 4901 31626
rect 4711 31562 4717 31574
rect 4895 31562 4901 31574
rect 4711 31510 4712 31562
rect 4900 31510 4901 31562
rect 4711 31498 4717 31510
rect 4895 31498 4901 31510
rect 4711 31446 4712 31498
rect 4900 31446 4901 31498
rect 4711 31434 4717 31446
rect 4895 31434 4901 31446
rect 4711 31382 4712 31434
rect 4900 31382 4901 31434
rect 4711 31370 4717 31382
rect 4895 31370 4901 31382
rect 4711 31318 4712 31370
rect 4900 31318 4901 31370
rect 4711 31306 4717 31318
rect 4895 31306 4901 31318
rect 4711 31254 4712 31306
rect 4900 31254 4901 31306
rect 4711 31242 4717 31254
rect 4895 31242 4901 31254
rect 4711 31190 4712 31242
rect 4900 31190 4901 31242
rect 4711 31178 4717 31190
rect 4895 31178 4901 31190
rect 4711 31126 4712 31178
rect 4900 31126 4901 31178
rect 4711 31114 4717 31126
rect 4895 31114 4901 31126
rect 4711 31062 4712 31114
rect 4900 31062 4901 31114
rect 4711 31050 4717 31062
rect 4895 31050 4901 31062
rect 4711 30998 4712 31050
rect 4900 30998 4901 31050
rect 4711 30986 4717 30998
rect 4895 30986 4901 30998
rect 4711 30934 4712 30986
rect 4900 30934 4901 30986
rect 4711 30922 4717 30934
rect 4895 30922 4901 30934
rect 4711 30870 4712 30922
rect 4900 30870 4901 30922
rect 4711 30858 4717 30870
rect 4895 30858 4901 30870
rect 4711 30806 4712 30858
rect 4900 30806 4901 30858
rect 4711 30794 4717 30806
rect 4895 30794 4901 30806
rect 4711 30742 4712 30794
rect 4900 30742 4901 30794
rect 4711 30729 4717 30742
rect 4895 30729 4901 30742
rect 4711 30677 4712 30729
rect 4900 30677 4901 30729
rect 4711 30664 4717 30677
rect 4895 30664 4901 30677
rect 4711 30612 4712 30664
rect 4900 30612 4901 30664
rect 4711 30599 4717 30612
rect 4895 30599 4901 30612
rect 4711 30547 4712 30599
rect 4900 30547 4901 30599
rect 4711 30534 4717 30547
rect 4895 30534 4901 30547
rect 4711 30482 4712 30534
rect 4900 30482 4901 30534
rect 4711 30469 4717 30482
rect 4895 30469 4901 30482
rect 4711 30417 4712 30469
rect 4900 30417 4901 30469
rect 4711 30404 4717 30417
rect 4895 30404 4901 30417
rect 4711 30352 4712 30404
rect 4900 30352 4901 30404
rect 4711 30339 4717 30352
rect 4895 30339 4901 30352
rect 4711 30287 4712 30339
rect 4900 30287 4901 30339
rect 4711 30274 4717 30287
rect 4895 30274 4901 30287
rect 4711 30222 4712 30274
rect 4900 30222 4901 30274
rect 4711 30209 4717 30222
rect 4895 30209 4901 30222
rect 4711 30157 4712 30209
rect 4900 30157 4901 30209
rect 4711 30144 4717 30157
rect 4895 30144 4901 30157
rect 4711 30092 4712 30144
rect 4900 30092 4901 30144
rect 4711 30079 4717 30092
rect 4895 30079 4901 30092
rect 4711 30027 4712 30079
rect 4900 30027 4901 30079
rect 4711 30014 4717 30027
rect 4895 30014 4901 30027
rect 4711 29962 4712 30014
rect 4900 29962 4901 30014
rect 4711 27903 4717 29962
rect 4895 27903 4901 29962
rect 2308 27826 2314 27860
rect 2348 27826 2386 27860
rect 2420 27826 2426 27860
rect 2308 27787 2426 27826
rect 2308 27753 2314 27787
rect 2348 27753 2386 27787
rect 2420 27753 2426 27787
rect 2308 27714 2426 27753
rect 2308 27680 2314 27714
rect 2348 27680 2386 27714
rect 2420 27680 2426 27714
rect 2308 27641 2426 27680
rect 2308 27607 2314 27641
rect 2348 27607 2386 27641
rect 2420 27607 2426 27641
rect 2308 27568 2426 27607
rect 2308 27534 2314 27568
rect 2348 27534 2386 27568
rect 2420 27534 2426 27568
rect 2308 27495 2426 27534
rect 2308 27461 2314 27495
rect 2348 27461 2386 27495
rect 2420 27461 2426 27495
rect 2308 27422 2426 27461
rect 2308 27388 2314 27422
rect 2348 27388 2386 27422
rect 2420 27388 2426 27422
rect 2308 27349 2426 27388
rect 2308 27315 2314 27349
rect 2348 27315 2386 27349
rect 2420 27315 2426 27349
rect 2308 27276 2426 27315
rect 3158 27574 3366 27580
rect 3158 27540 3170 27574
rect 3204 27540 3245 27574
rect 3279 27540 3320 27574
rect 3354 27540 3366 27574
rect 3158 27534 3366 27540
rect 3158 27502 3241 27534
tri 3241 27502 3273 27534 nw
rect 2308 27242 2314 27276
rect 2348 27242 2386 27276
rect 2420 27252 2426 27276
tri 2426 27252 2457 27283 sw
rect 2420 27242 2457 27252
rect 2308 27231 2457 27242
tri 2457 27231 2478 27252 sw
rect 2308 27209 2478 27231
tri 2478 27209 2500 27231 sw
rect 2308 27203 2833 27209
rect 2308 27169 2314 27203
rect 2348 27169 2386 27203
rect 2420 27169 2471 27203
rect 2505 27169 2550 27203
rect 2584 27169 2629 27203
rect 2663 27169 2708 27203
rect 2742 27169 2787 27203
rect 2821 27169 2833 27203
rect 2308 27131 2833 27169
rect 2308 27097 2392 27131
rect 2426 27097 2471 27131
rect 2505 27097 2550 27131
rect 2584 27097 2629 27131
rect 2663 27097 2708 27131
rect 2742 27097 2787 27131
rect 2821 27097 2833 27131
rect 2308 27091 2833 27097
rect 1834 27073 1986 27078
rect 1834 27039 1946 27073
rect 1980 27039 1986 27073
rect 1834 27005 1840 27039
rect 1874 27005 1986 27039
rect 1834 27000 1986 27005
rect 1834 26966 1946 27000
rect 1980 26966 1986 27000
rect 1834 26932 1840 26966
rect 1874 26932 1986 26966
rect 1834 26927 1986 26932
rect 1834 26893 1946 26927
rect 1980 26893 1986 26927
rect 1834 26859 1840 26893
rect 1874 26859 1986 26893
rect 1834 26854 1986 26859
rect 1834 26820 1946 26854
rect 1980 26820 1986 26854
rect 1834 26786 1840 26820
rect 1874 26787 1986 26820
tri 1986 26787 2060 26861 sw
rect 1874 26786 2850 26787
rect 1834 26781 2850 26786
rect 1834 26747 1946 26781
rect 1980 26747 2024 26781
rect 2058 26747 2102 26781
rect 2136 26747 2180 26781
rect 2214 26747 2258 26781
rect 2292 26747 2336 26781
rect 2370 26747 2414 26781
rect 2448 26747 2492 26781
rect 2526 26747 2570 26781
rect 2604 26747 2648 26781
rect 2682 26747 2726 26781
rect 2760 26747 2804 26781
rect 2838 26747 2850 26781
rect 1834 26713 1840 26747
rect 1874 26713 2850 26747
rect 1834 26675 2850 26713
rect 1834 26641 1914 26675
rect 1948 26641 1988 26675
rect 2022 26641 2062 26675
rect 2096 26641 2136 26675
rect 2170 26641 2210 26675
rect 2244 26641 2284 26675
rect 2318 26641 2358 26675
rect 2392 26641 2432 26675
rect 2466 26641 2506 26675
rect 2540 26641 2580 26675
rect 2614 26641 2654 26675
rect 2688 26641 2729 26675
rect 2763 26641 2804 26675
rect 2838 26641 2850 26675
rect 1834 26635 2850 26641
tri 1498 26341 1499 26342 sw
tri 3157 26341 3158 26342 se
rect 3158 26341 3239 27502
tri 3239 27500 3241 27502 nw
rect 4711 27367 4901 27903
tri 4711 27358 4720 27367 ne
rect 4720 27358 4901 27367
tri 4720 27324 4754 27358 ne
rect 4754 27324 4901 27358
tri 4754 27301 4777 27324 ne
rect 3572 27231 4477 27237
rect 3572 27197 3584 27231
rect 3618 27197 3662 27231
rect 3696 27197 3740 27231
rect 3774 27197 3818 27231
rect 3852 27197 3896 27231
rect 3930 27197 3974 27231
rect 4008 27197 4052 27231
rect 4086 27197 4130 27231
rect 4164 27197 4208 27231
rect 4242 27197 4286 27231
rect 4320 27197 4363 27231
rect 4397 27197 4477 27231
rect 3572 27123 4477 27197
rect 3572 27089 3584 27123
rect 3618 27089 3662 27123
rect 3696 27089 3740 27123
rect 3774 27089 3818 27123
rect 3852 27089 3896 27123
rect 3930 27089 3974 27123
rect 4008 27089 4052 27123
rect 4086 27089 4130 27123
rect 4164 27089 4208 27123
rect 4242 27089 4286 27123
rect 4320 27089 4363 27123
rect 4397 27089 4477 27123
rect 3572 27083 4477 27089
tri 4261 27059 4285 27083 ne
rect 4285 27059 4477 27083
tri 4285 27055 4289 27059 ne
rect 4289 27055 4477 27059
tri 4289 27047 4297 27055 ne
rect 4297 27047 4477 27055
tri 4297 26985 4359 27047 ne
rect 3555 26769 4059 26775
rect 3555 26735 3567 26769
rect 3601 26735 3643 26769
rect 3677 26735 3719 26769
rect 3753 26735 3795 26769
rect 3829 26735 3871 26769
rect 3905 26735 3947 26769
rect 3981 26735 4059 26769
rect 3555 26697 4059 26735
rect 3555 26663 4019 26697
rect 4053 26663 4059 26697
rect 3555 26629 3567 26663
rect 3601 26629 3653 26663
rect 3687 26629 3739 26663
rect 3773 26629 3826 26663
rect 3860 26629 3913 26663
rect 3947 26629 4059 26663
rect 3555 26625 4059 26629
rect 3555 26623 4019 26625
tri 3873 26591 3905 26623 ne
rect 3905 26591 4019 26623
rect 4053 26591 4059 26625
tri 3905 26589 3907 26591 ne
rect 3907 26557 3913 26591
rect 3947 26557 4059 26591
rect 3907 26553 4059 26557
rect 3907 26519 4019 26553
rect 4053 26519 4059 26553
rect 3907 26485 3913 26519
rect 3947 26485 4059 26519
rect 3907 26481 4059 26485
rect 3907 26447 4019 26481
rect 4053 26447 4059 26481
rect 3907 26413 3913 26447
rect 3947 26413 4059 26447
rect 3907 26409 4059 26413
rect 3907 26375 4019 26409
rect 4053 26375 4059 26409
tri 3239 26341 3240 26342 sw
rect 3907 26341 3913 26375
rect 3947 26341 4059 26375
rect 1418 26337 1499 26341
tri 1499 26337 1503 26341 sw
tri 3153 26337 3157 26341 se
rect 3157 26337 3240 26341
tri 3240 26337 3244 26341 sw
rect 3907 26337 4059 26341
rect 1418 26308 1503 26337
tri 1503 26308 1532 26337 sw
tri 3124 26308 3153 26337 se
rect 3153 26308 3244 26337
tri 3244 26308 3273 26337 sw
rect 1418 26228 3521 26308
tri 3407 26197 3438 26228 ne
rect 3438 26197 3521 26228
tri 3438 26194 3441 26197 ne
rect 3441 23432 3521 26197
rect 3441 23380 3456 23432
rect 3508 23380 3521 23432
rect 3441 23357 3521 23380
rect 3441 23305 3456 23357
rect 3508 23305 3521 23357
rect 3441 23282 3521 23305
rect 3441 23230 3456 23282
rect 3508 23230 3521 23282
rect 222 14870 1999 14877
rect 222 14836 1881 14870
rect 1915 14836 1953 14870
rect 1987 14836 1999 14870
rect 222 14829 1999 14836
rect 222 14822 320 14829
tri 320 14822 327 14829 nw
rect 222 14796 294 14822
tri 294 14796 320 14822 nw
rect 222 14785 283 14796
tri 283 14785 294 14796 nw
rect 222 14784 282 14785
tri 282 14784 283 14785 nw
rect 222 14783 281 14784
tri 281 14783 282 14784 nw
rect 222 8762 270 14783
tri 270 14772 281 14783 nw
tri 3426 14749 3441 14764 se
rect 3441 14749 3521 23230
rect 3907 26303 4019 26337
rect 4053 26303 4059 26337
rect 3907 26269 3913 26303
rect 3947 26269 4059 26303
rect 3907 26265 4059 26269
rect 3907 26231 4019 26265
rect 4053 26231 4059 26265
rect 3907 26197 3913 26231
rect 3947 26197 4059 26231
rect 3907 26193 4059 26197
rect 3907 26159 4019 26193
rect 4053 26159 4059 26193
rect 3907 26125 3913 26159
rect 3947 26125 4059 26159
rect 3907 26121 4059 26125
rect 3907 26087 4019 26121
rect 4053 26087 4059 26121
rect 3907 26053 3913 26087
rect 3947 26053 4059 26087
rect 3907 26049 4059 26053
rect 3907 26015 4019 26049
rect 4053 26015 4059 26049
rect 3907 25981 3913 26015
rect 3947 25981 4059 26015
rect 3907 25977 4059 25981
rect 3907 25943 4019 25977
rect 4053 25943 4059 25977
rect 3907 25909 3913 25943
rect 3947 25909 4059 25943
rect 3907 25905 4059 25909
rect 3907 25871 4019 25905
rect 4053 25871 4059 25905
rect 3907 25837 3913 25871
rect 3947 25837 4059 25871
rect 3907 25833 4059 25837
rect 3907 25799 4019 25833
rect 4053 25799 4059 25833
rect 3907 25765 3913 25799
rect 3947 25765 4059 25799
rect 3907 25761 4059 25765
rect 3907 25727 4019 25761
rect 4053 25727 4059 25761
rect 3907 25693 3913 25727
rect 3947 25693 4059 25727
rect 3907 25689 4059 25693
rect 3907 25655 4019 25689
rect 4053 25655 4059 25689
rect 3907 25621 3913 25655
rect 3947 25621 4059 25655
rect 3907 25617 4059 25621
rect 3907 25583 4019 25617
rect 4053 25583 4059 25617
rect 3907 25549 3913 25583
rect 3947 25549 4059 25583
rect 3907 25545 4059 25549
rect 3907 25511 4019 25545
rect 4053 25511 4059 25545
rect 3907 25477 3913 25511
rect 3947 25477 4059 25511
rect 3907 25473 4059 25477
rect 3907 25439 4019 25473
rect 4053 25439 4059 25473
rect 3907 25405 3913 25439
rect 3947 25405 4059 25439
rect 3907 25401 4059 25405
rect 3907 25367 4019 25401
rect 4053 25367 4059 25401
rect 3907 25333 3913 25367
rect 3947 25333 4059 25367
rect 3907 25329 4059 25333
rect 3907 25295 4019 25329
rect 4053 25295 4059 25329
rect 3907 25261 3913 25295
rect 3947 25261 4059 25295
rect 3907 25257 4059 25261
rect 3907 25223 4019 25257
rect 4053 25223 4059 25257
rect 3907 25189 3913 25223
rect 3947 25189 4059 25223
rect 3907 25185 4059 25189
rect 3907 25151 4019 25185
rect 4053 25151 4059 25185
rect 3907 25117 3913 25151
rect 3947 25117 4059 25151
rect 3907 25113 4059 25117
rect 3907 25079 4019 25113
rect 4053 25079 4059 25113
rect 3907 25045 3913 25079
rect 3947 25045 4059 25079
rect 3907 25041 4059 25045
rect 3907 25007 4019 25041
rect 4053 25007 4059 25041
rect 3907 24973 3913 25007
rect 3947 24973 4059 25007
rect 3907 24969 4059 24973
rect 3907 24935 4019 24969
rect 4053 24935 4059 24969
rect 3907 24901 3913 24935
rect 3947 24901 4059 24935
rect 3907 24897 4059 24901
rect 3907 24863 4019 24897
rect 4053 24863 4059 24897
rect 3907 24829 3913 24863
rect 3947 24829 4059 24863
rect 3907 24825 4059 24829
rect 3907 24791 4019 24825
rect 4053 24791 4059 24825
rect 3907 24757 3913 24791
rect 3947 24757 4059 24791
rect 3907 24753 4059 24757
rect 3907 24719 4019 24753
rect 4053 24719 4059 24753
rect 3907 24685 3913 24719
rect 3947 24685 4059 24719
rect 3907 24681 4059 24685
rect 3907 24647 4019 24681
rect 4053 24647 4059 24681
rect 3907 24613 3913 24647
rect 3947 24613 4059 24647
rect 3907 24609 4059 24613
rect 3907 24575 4019 24609
rect 4053 24575 4059 24609
rect 3907 24541 3913 24575
rect 3947 24541 4059 24575
rect 3907 24537 4059 24541
rect 3907 24503 4019 24537
rect 4053 24503 4059 24537
rect 3907 24469 3913 24503
rect 3947 24469 4059 24503
rect 3907 24465 4059 24469
rect 3907 24431 4019 24465
rect 4053 24431 4059 24465
rect 3907 24397 3913 24431
rect 3947 24397 4059 24431
rect 3907 24393 4059 24397
rect 3907 24359 4019 24393
rect 4053 24359 4059 24393
rect 3907 24325 3913 24359
rect 3947 24325 4059 24359
rect 3907 24321 4059 24325
rect 3907 24287 4019 24321
rect 4053 24287 4059 24321
rect 3907 24253 3913 24287
rect 3947 24253 4059 24287
rect 3907 24249 4059 24253
rect 3907 24215 4019 24249
rect 4053 24215 4059 24249
rect 3907 24181 3913 24215
rect 3947 24181 4059 24215
rect 3907 24177 4059 24181
rect 3907 24143 4019 24177
rect 4053 24143 4059 24177
rect 3907 24109 3913 24143
rect 3947 24109 4059 24143
rect 3907 24105 4059 24109
rect 3907 24071 4019 24105
rect 4053 24071 4059 24105
rect 3907 24037 3913 24071
rect 3947 24037 4059 24071
rect 3907 24033 4059 24037
rect 3907 23999 4019 24033
rect 4053 23999 4059 24033
rect 3907 23965 3913 23999
rect 3947 23965 4059 23999
rect 3907 23961 4059 23965
rect 3907 23927 4019 23961
rect 4053 23927 4059 23961
rect 3907 23893 3913 23927
rect 3947 23893 4059 23927
rect 3907 23889 4059 23893
rect 3907 23855 4019 23889
rect 4053 23855 4059 23889
rect 3907 23821 3913 23855
rect 3947 23821 4059 23855
rect 3907 23817 4059 23821
rect 3907 23783 4019 23817
rect 4053 23783 4059 23817
rect 3907 23749 3913 23783
rect 3947 23749 4059 23783
rect 3907 23745 4059 23749
rect 3907 23711 4019 23745
rect 4053 23711 4059 23745
rect 3907 23677 3913 23711
rect 3947 23677 4059 23711
rect 3907 23673 4059 23677
rect 3907 23639 4019 23673
rect 4053 23639 4059 23673
rect 3907 23605 3913 23639
rect 3947 23605 4059 23639
rect 3907 23601 4059 23605
rect 3907 23567 4019 23601
rect 4053 23567 4059 23601
rect 3907 23533 3913 23567
rect 3947 23533 4059 23567
rect 3907 23529 4059 23533
rect 3907 23495 4019 23529
rect 4053 23495 4059 23529
rect 3907 23461 3913 23495
rect 3947 23461 4059 23495
rect 3907 23457 4059 23461
rect 3907 23423 4019 23457
rect 4053 23423 4059 23457
rect 3907 23389 3913 23423
rect 3947 23389 4059 23423
rect 3907 23385 4059 23389
rect 3907 23351 4019 23385
rect 4053 23351 4059 23385
rect 3907 23317 3913 23351
rect 3947 23317 4059 23351
rect 3907 23313 4059 23317
rect 3907 23279 4019 23313
rect 4053 23279 4059 23313
rect 3907 23245 3913 23279
rect 3947 23245 4059 23279
rect 3907 23241 4059 23245
rect 3907 23207 4019 23241
rect 4053 23207 4059 23241
rect 3907 23173 3913 23207
rect 3947 23173 4059 23207
rect 3907 23169 4059 23173
rect 3907 23135 4019 23169
rect 4053 23135 4059 23169
rect 3907 23101 3913 23135
rect 3947 23101 4059 23135
rect 3907 23097 4059 23101
rect 3907 23063 4019 23097
rect 4053 23063 4059 23097
rect 3907 23029 3913 23063
rect 3947 23029 4059 23063
rect 3907 23025 4059 23029
rect 3907 22991 4019 23025
rect 4053 22991 4059 23025
rect 3907 22957 3913 22991
rect 3947 22957 4059 22991
rect 3907 22953 4059 22957
rect 3907 22919 4019 22953
rect 4053 22919 4059 22953
rect 3907 22885 3913 22919
rect 3947 22885 4059 22919
rect 3907 22881 4059 22885
rect 3907 22847 4019 22881
rect 4053 22847 4059 22881
rect 3907 22813 3913 22847
rect 3947 22813 4059 22847
rect 3907 22809 4059 22813
rect 3907 22775 4019 22809
rect 4053 22775 4059 22809
rect 3907 22741 3913 22775
rect 3947 22741 4059 22775
rect 3907 22737 4059 22741
rect 3907 22703 4019 22737
rect 4053 22703 4059 22737
rect 3907 22669 3913 22703
rect 3947 22669 4059 22703
rect 3907 22665 4059 22669
rect 3907 22631 4019 22665
rect 4053 22631 4059 22665
rect 3907 22597 3913 22631
rect 3947 22597 4059 22631
rect 3907 22593 4059 22597
rect 3907 22559 4019 22593
rect 4053 22559 4059 22593
rect 3907 22525 3913 22559
rect 3947 22525 4059 22559
rect 3907 22521 4059 22525
rect 3907 22487 4019 22521
rect 4053 22487 4059 22521
rect 3907 22453 3913 22487
rect 3947 22453 4059 22487
rect 3907 22449 4059 22453
rect 3907 22415 4019 22449
rect 4053 22415 4059 22449
rect 3907 22381 3913 22415
rect 3947 22381 4059 22415
rect 3907 22377 4059 22381
rect 3907 22343 4019 22377
rect 4053 22343 4059 22377
rect 3907 22309 3913 22343
rect 3947 22309 4059 22343
rect 3907 22305 4059 22309
rect 3907 22271 4019 22305
rect 4053 22271 4059 22305
rect 3907 22237 3913 22271
rect 3947 22237 4059 22271
rect 3907 22233 4059 22237
rect 3907 22199 4019 22233
rect 4053 22199 4059 22233
rect 3907 22165 3913 22199
rect 3947 22165 4059 22199
rect 3907 22161 4059 22165
rect 3907 22127 4019 22161
rect 4053 22127 4059 22161
rect 3907 22093 3913 22127
rect 3947 22093 4059 22127
rect 3907 22089 4059 22093
rect 3907 22055 4019 22089
rect 4053 22055 4059 22089
rect 3907 22021 3913 22055
rect 3947 22021 4059 22055
rect 3907 22016 4059 22021
rect 3907 21983 4019 22016
rect 3907 21949 3913 21983
rect 3947 21982 4019 21983
rect 4053 21982 4059 22016
rect 3947 21949 4059 21982
rect 3907 21943 4059 21949
rect 3907 21911 4019 21943
rect 3907 21877 3913 21911
rect 3947 21909 4019 21911
rect 4053 21909 4059 21943
rect 3947 21877 4059 21909
rect 3907 21870 4059 21877
rect 3907 21839 4019 21870
rect 3907 21805 3913 21839
rect 3947 21836 4019 21839
rect 4053 21836 4059 21870
rect 3947 21805 4059 21836
rect 3907 21797 4059 21805
rect 3907 21767 4019 21797
rect 3907 21733 3913 21767
rect 3947 21763 4019 21767
rect 4053 21763 4059 21797
rect 3947 21733 4059 21763
rect 3907 21724 4059 21733
rect 3907 21695 4019 21724
rect 3907 21661 3913 21695
rect 3947 21690 4019 21695
rect 4053 21690 4059 21724
rect 3947 21661 4059 21690
rect 3907 21651 4059 21661
rect 3907 21623 4019 21651
rect 3907 21589 3913 21623
rect 3947 21617 4019 21623
rect 4053 21617 4059 21651
rect 3947 21589 4059 21617
rect 3907 21578 4059 21589
rect 3907 21551 4019 21578
rect 3907 21517 3913 21551
rect 3947 21544 4019 21551
rect 4053 21544 4059 21578
rect 3947 21517 4059 21544
rect 3907 21505 4059 21517
rect 3907 21479 4019 21505
rect 3907 21445 3913 21479
rect 3947 21471 4019 21479
rect 4053 21471 4059 21505
rect 3947 21445 4059 21471
rect 3907 21432 4059 21445
rect 3907 21407 4019 21432
rect 3907 21373 3913 21407
rect 3947 21398 4019 21407
rect 4053 21398 4059 21432
rect 3947 21373 4059 21398
rect 3907 21359 4059 21373
rect 3907 21335 4019 21359
rect 3907 21301 3913 21335
rect 3947 21325 4019 21335
rect 4053 21325 4059 21359
rect 3947 21301 4059 21325
rect 3907 21286 4059 21301
rect 3907 21263 4019 21286
rect 3907 21229 3913 21263
rect 3947 21252 4019 21263
rect 4053 21252 4059 21286
rect 3947 21229 4059 21252
rect 3907 21213 4059 21229
rect 3907 21191 4019 21213
rect 3907 21157 3913 21191
rect 3947 21179 4019 21191
rect 4053 21179 4059 21213
rect 3947 21157 4059 21179
rect 3907 21140 4059 21157
rect 3907 21119 4019 21140
rect 3907 21085 3913 21119
rect 3947 21106 4019 21119
rect 4053 21106 4059 21140
rect 3947 21085 4059 21106
rect 3907 21067 4059 21085
rect 3907 21047 4019 21067
rect 3907 21013 3913 21047
rect 3947 21033 4019 21047
rect 4053 21033 4059 21067
rect 3947 21013 4059 21033
rect 3907 20994 4059 21013
rect 3907 20975 4019 20994
rect 3907 20941 3913 20975
rect 3947 20960 4019 20975
rect 4053 20960 4059 20994
rect 3947 20941 4059 20960
rect 3907 20921 4059 20941
rect 3907 20903 4019 20921
rect 3907 20869 3913 20903
rect 3947 20887 4019 20903
rect 4053 20887 4059 20921
rect 3947 20869 4059 20887
rect 3907 20848 4059 20869
rect 3907 20831 4019 20848
rect 3907 20797 3913 20831
rect 3947 20814 4019 20831
rect 4053 20814 4059 20848
rect 3947 20797 4059 20814
rect 3907 20775 4059 20797
rect 3907 20759 4019 20775
rect 3907 20725 3913 20759
rect 3947 20741 4019 20759
rect 4053 20741 4059 20775
rect 3947 20725 4059 20741
rect 3907 20702 4059 20725
rect 3907 20687 4019 20702
rect 3907 20653 3913 20687
rect 3947 20668 4019 20687
rect 4053 20668 4059 20702
rect 3947 20653 4059 20668
rect 3907 20629 4059 20653
rect 3907 20615 4019 20629
rect 3907 20581 3913 20615
rect 3947 20595 4019 20615
rect 4053 20595 4059 20629
rect 3947 20581 4059 20595
rect 3907 20556 4059 20581
rect 3907 20543 4019 20556
rect 3907 20509 3913 20543
rect 3947 20522 4019 20543
rect 4053 20522 4059 20556
rect 3947 20509 4059 20522
rect 3907 20483 4059 20509
rect 3907 20471 4019 20483
rect 3907 20437 3913 20471
rect 3947 20449 4019 20471
rect 4053 20449 4059 20483
rect 3947 20437 4059 20449
rect 3907 20410 4059 20437
rect 3907 20399 4019 20410
rect 3907 20365 3913 20399
rect 3947 20376 4019 20399
rect 4053 20376 4059 20410
rect 3947 20365 4059 20376
rect 3907 20337 4059 20365
rect 3907 20327 4019 20337
rect 3907 20293 3913 20327
rect 3947 20303 4019 20327
rect 4053 20303 4059 20337
rect 3947 20293 4059 20303
rect 3907 20264 4059 20293
rect 3907 20255 4019 20264
rect 3907 20221 3913 20255
rect 3947 20230 4019 20255
rect 4053 20230 4059 20264
rect 3947 20221 4059 20230
rect 3907 20191 4059 20221
rect 3907 20183 4019 20191
rect 3907 20149 3913 20183
rect 3947 20157 4019 20183
rect 4053 20157 4059 20191
rect 3947 20149 4059 20157
rect 3907 20118 4059 20149
rect 3907 20111 4019 20118
rect 3907 20077 3913 20111
rect 3947 20084 4019 20111
rect 4053 20084 4059 20118
rect 3947 20077 4059 20084
rect 3907 20045 4059 20077
rect 3907 20039 4019 20045
rect 3907 20005 3913 20039
rect 3947 20011 4019 20039
rect 4053 20011 4059 20045
rect 3947 20005 4059 20011
rect 3907 19972 4059 20005
rect 3907 19967 4019 19972
rect 3907 19933 3913 19967
rect 3947 19938 4019 19967
rect 4053 19938 4059 19972
rect 3947 19933 4059 19938
rect 3907 19899 4059 19933
rect 3907 19895 4019 19899
rect 3907 19861 3913 19895
rect 3947 19865 4019 19895
rect 4053 19865 4059 19899
rect 3947 19861 4059 19865
rect 3907 19826 4059 19861
rect 3907 19823 4019 19826
rect 3907 19789 3913 19823
rect 3947 19792 4019 19823
rect 4053 19792 4059 19826
rect 3947 19789 4059 19792
rect 3907 19753 4059 19789
rect 3907 19751 4019 19753
rect 3907 19717 3913 19751
rect 3947 19719 4019 19751
rect 4053 19719 4059 19753
rect 3947 19717 4059 19719
rect 3907 19680 4059 19717
rect 3907 19679 4019 19680
rect 3907 19645 3913 19679
rect 3947 19646 4019 19679
rect 4053 19646 4059 19680
rect 3947 19645 4059 19646
rect 3907 19607 4059 19645
rect 3907 19573 3913 19607
rect 3947 19573 4019 19607
rect 4053 19573 4059 19607
rect 3907 19534 4059 19573
rect 3907 19500 3913 19534
rect 3947 19500 4019 19534
rect 4053 19500 4059 19534
rect 4359 23557 4365 27047
rect 4471 23557 4477 27047
rect 4359 23518 4477 23557
rect 4359 23484 4365 23518
rect 4399 23484 4437 23518
rect 4471 23484 4477 23518
rect 4359 23445 4477 23484
rect 4359 23411 4365 23445
rect 4399 23411 4437 23445
rect 4471 23411 4477 23445
rect 4359 23372 4477 23411
rect 4359 23338 4365 23372
rect 4399 23338 4437 23372
rect 4471 23338 4477 23372
rect 4359 23299 4477 23338
rect 4777 27162 4901 27324
rect 4777 27128 4783 27162
rect 4817 27128 4861 27162
rect 4895 27128 4901 27162
rect 4777 27090 4901 27128
rect 4777 27038 4780 27090
rect 4832 27038 4848 27090
rect 4900 27038 4901 27090
rect 4777 27026 4901 27038
rect 4777 26974 4780 27026
rect 4832 26974 4848 27026
rect 4900 26974 4901 27026
rect 4777 26962 4901 26974
rect 4777 26910 4780 26962
rect 4832 26910 4848 26962
rect 4900 26910 4901 26962
rect 4777 26909 4783 26910
rect 4817 26909 4861 26910
rect 4895 26909 4901 26910
rect 4777 26898 4901 26909
rect 4777 26846 4780 26898
rect 4832 26846 4848 26898
rect 4900 26846 4901 26898
rect 4777 26836 4783 26846
rect 4817 26836 4861 26846
rect 4895 26836 4901 26846
rect 4777 26834 4901 26836
rect 4777 26782 4780 26834
rect 4832 26782 4848 26834
rect 4900 26782 4901 26834
rect 4777 26770 4783 26782
rect 4817 26770 4861 26782
rect 4895 26770 4901 26782
rect 4777 26718 4780 26770
rect 4832 26718 4848 26770
rect 4900 26718 4901 26770
rect 4777 26706 4783 26718
rect 4817 26706 4861 26718
rect 4895 26706 4901 26718
rect 4777 26654 4780 26706
rect 4832 26654 4848 26706
rect 4900 26654 4901 26706
rect 4777 26651 4901 26654
rect 4777 26642 4783 26651
rect 4817 26642 4861 26651
rect 4895 26642 4901 26651
rect 4777 26590 4780 26642
rect 4832 26590 4848 26642
rect 4900 26590 4901 26642
rect 4777 26578 4901 26590
rect 4777 26526 4780 26578
rect 4832 26526 4848 26578
rect 4900 26526 4901 26578
rect 4777 26514 4901 26526
rect 4777 26462 4780 26514
rect 4832 26462 4848 26514
rect 4900 26462 4901 26514
rect 4777 26450 4901 26462
rect 4777 26398 4780 26450
rect 4832 26398 4848 26450
rect 4900 26398 4901 26450
rect 4777 26386 4901 26398
rect 4777 26334 4780 26386
rect 4832 26334 4848 26386
rect 4900 26334 4901 26386
rect 4777 26325 4783 26334
rect 4817 26325 4861 26334
rect 4895 26325 4901 26334
rect 4777 26322 4901 26325
rect 4777 26270 4780 26322
rect 4832 26270 4848 26322
rect 4900 26270 4901 26322
rect 4777 26258 4783 26270
rect 4817 26258 4861 26270
rect 4895 26258 4901 26270
rect 4777 26206 4780 26258
rect 4832 26206 4848 26258
rect 4900 26206 4901 26258
rect 4777 26194 4783 26206
rect 4817 26194 4861 26206
rect 4895 26194 4901 26206
rect 4777 26142 4780 26194
rect 4832 26142 4848 26194
rect 4900 26142 4901 26194
rect 4777 26140 4901 26142
rect 4777 26129 4783 26140
rect 4817 26129 4861 26140
rect 4895 26129 4901 26140
rect 4777 26077 4780 26129
rect 4832 26077 4848 26129
rect 4900 26077 4901 26129
rect 4777 26067 4901 26077
rect 4777 26064 4783 26067
rect 4817 26064 4861 26067
rect 4895 26064 4901 26067
rect 4777 26012 4780 26064
rect 4832 26012 4848 26064
rect 4900 26012 4901 26064
rect 4777 25999 4901 26012
rect 4777 25947 4780 25999
rect 4832 25947 4848 25999
rect 4900 25947 4901 25999
rect 4777 25934 4901 25947
rect 4777 25882 4780 25934
rect 4832 25882 4848 25934
rect 4900 25882 4901 25934
rect 4777 25869 4901 25882
rect 4777 25817 4780 25869
rect 4832 25817 4848 25869
rect 4900 25817 4901 25869
rect 4777 25814 4783 25817
rect 4817 25814 4861 25817
rect 4895 25814 4901 25817
rect 4777 25804 4901 25814
rect 4777 25752 4780 25804
rect 4832 25752 4848 25804
rect 4900 25752 4901 25804
rect 4777 25741 4783 25752
rect 4817 25741 4861 25752
rect 4895 25741 4901 25752
rect 4777 25739 4901 25741
rect 4777 25687 4780 25739
rect 4832 25687 4848 25739
rect 4900 25687 4901 25739
rect 4777 25674 4783 25687
rect 4817 25674 4861 25687
rect 4895 25674 4901 25687
rect 4777 25622 4780 25674
rect 4832 25622 4848 25674
rect 4900 25622 4901 25674
rect 4777 25609 4783 25622
rect 4817 25609 4861 25622
rect 4895 25609 4901 25622
rect 4777 25557 4780 25609
rect 4832 25557 4848 25609
rect 4900 25557 4901 25609
rect 4777 25556 4901 25557
rect 4777 25544 4783 25556
rect 4817 25544 4861 25556
rect 4895 25544 4901 25556
rect 4777 25492 4780 25544
rect 4832 25492 4848 25544
rect 4900 25492 4901 25544
rect 4777 25483 4901 25492
rect 4777 25479 4783 25483
rect 4817 25479 4861 25483
rect 4895 25479 4901 25483
rect 4777 25427 4780 25479
rect 4832 25427 4848 25479
rect 4900 25427 4901 25479
rect 4777 25414 4901 25427
rect 4777 25362 4780 25414
rect 4832 25362 4848 25414
rect 4900 25362 4901 25414
rect 4777 25337 4901 25362
rect 4777 25303 4783 25337
rect 4817 25303 4861 25337
rect 4895 25303 4901 25337
rect 4777 25264 4901 25303
rect 4777 25230 4783 25264
rect 4817 25230 4861 25264
rect 4895 25230 4901 25264
rect 4777 25191 4901 25230
rect 4777 25157 4783 25191
rect 4817 25157 4861 25191
rect 4895 25157 4901 25191
rect 4777 25118 4901 25157
rect 4777 25084 4783 25118
rect 4817 25084 4861 25118
rect 4895 25084 4901 25118
rect 4777 25045 4901 25084
rect 4777 25011 4783 25045
rect 4817 25011 4861 25045
rect 4895 25011 4901 25045
rect 4777 24972 4901 25011
rect 4777 24938 4783 24972
rect 4817 24938 4861 24972
rect 4895 24938 4901 24972
rect 4777 24899 4901 24938
rect 4777 24865 4783 24899
rect 4817 24865 4861 24899
rect 4895 24865 4901 24899
rect 4777 24826 4901 24865
rect 4777 24792 4783 24826
rect 4817 24792 4861 24826
rect 4895 24792 4901 24826
rect 4777 24753 4901 24792
rect 4777 24719 4783 24753
rect 4817 24719 4861 24753
rect 4895 24719 4901 24753
rect 4777 24680 4901 24719
rect 4777 24646 4783 24680
rect 4817 24646 4861 24680
rect 4895 24646 4901 24680
rect 4777 24606 4901 24646
rect 4777 24572 4783 24606
rect 4817 24572 4861 24606
rect 4895 24572 4901 24606
rect 4777 24532 4901 24572
rect 4777 24498 4783 24532
rect 4817 24498 4861 24532
rect 4895 24498 4901 24532
rect 4777 24458 4901 24498
rect 4777 24424 4783 24458
rect 4817 24424 4861 24458
rect 4895 24424 4901 24458
rect 4777 24384 4901 24424
rect 4777 24350 4783 24384
rect 4817 24350 4861 24384
rect 4895 24350 4901 24384
rect 4777 24310 4901 24350
rect 4777 24276 4783 24310
rect 4817 24276 4861 24310
rect 4895 24276 4901 24310
rect 4777 24236 4901 24276
rect 4777 24202 4783 24236
rect 4817 24202 4861 24236
rect 4895 24202 4901 24236
rect 4777 24162 4901 24202
rect 4777 24128 4783 24162
rect 4817 24128 4861 24162
rect 4895 24128 4901 24162
rect 4777 24088 4901 24128
rect 4777 24054 4783 24088
rect 4817 24054 4861 24088
rect 4895 24054 4901 24088
rect 4777 24014 4901 24054
rect 4777 23980 4783 24014
rect 4817 23980 4861 24014
rect 4895 23980 4901 24014
rect 4777 23940 4901 23980
rect 4777 23906 4783 23940
rect 4817 23906 4861 23940
rect 4895 23906 4901 23940
rect 4777 23866 4901 23906
rect 4777 23832 4783 23866
rect 4817 23832 4861 23866
rect 4895 23832 4901 23866
rect 4777 23792 4901 23832
rect 4777 23758 4783 23792
rect 4817 23758 4861 23792
rect 4895 23758 4901 23792
rect 4777 23718 4901 23758
rect 4777 23684 4783 23718
rect 4817 23684 4861 23718
rect 4895 23684 4901 23718
rect 4777 23644 4901 23684
rect 4777 23610 4783 23644
rect 4817 23610 4861 23644
rect 4895 23610 4901 23644
rect 4777 23570 4901 23610
rect 4777 23536 4783 23570
rect 4817 23536 4861 23570
rect 4895 23536 4901 23570
rect 4777 23496 4901 23536
rect 4777 23462 4783 23496
rect 4817 23462 4861 23496
rect 4895 23462 4901 23496
rect 4777 23422 4901 23462
rect 4777 23388 4783 23422
rect 4817 23388 4861 23422
rect 4895 23388 4901 23422
rect 4777 23348 4901 23388
rect 4777 23314 4783 23348
rect 4817 23314 4861 23348
rect 4895 23314 4901 23348
rect 4777 23302 4901 23314
rect 5201 37997 5331 38003
rect 5253 37945 5279 37997
rect 5201 37929 5331 37945
rect 5253 37877 5279 37929
rect 5201 37861 5331 37877
rect 5253 37809 5279 37861
rect 5201 37793 5331 37809
rect 5253 37741 5279 37793
rect 5201 37725 5331 37741
rect 5253 37673 5279 37725
rect 5201 37657 5331 37673
rect 5253 37605 5279 37657
rect 5201 37589 5331 37605
rect 5253 37537 5279 37589
rect 5201 37521 5331 37537
rect 5253 37469 5279 37521
rect 5201 37453 5331 37469
rect 5253 37401 5279 37453
rect 5201 37385 5331 37401
rect 5253 37333 5279 37385
rect 5201 37318 5331 37333
rect 5253 37266 5279 37318
rect 5201 37251 5331 37266
rect 5253 37199 5279 37251
rect 5201 37184 5331 37199
rect 5253 37132 5279 37184
rect 5201 37117 5331 37132
rect 5253 37065 5279 37117
rect 5201 34225 5331 37065
rect 5253 34173 5279 34225
rect 5201 34161 5331 34173
rect 5253 34109 5279 34161
rect 5201 34097 5331 34109
rect 5253 34045 5279 34097
rect 5201 34033 5331 34045
rect 5253 33981 5279 34033
rect 5201 33969 5331 33981
rect 5253 33917 5279 33969
rect 5201 33905 5331 33917
rect 5253 33853 5279 33905
rect 5201 33841 5331 33853
rect 5253 33789 5279 33841
rect 5201 33777 5331 33789
rect 5253 33725 5279 33777
rect 5201 33713 5331 33725
rect 5253 33661 5279 33713
rect 5201 33649 5331 33661
rect 5253 33597 5279 33649
rect 5201 33585 5331 33597
rect 5253 33533 5279 33585
rect 5201 33521 5331 33533
rect 5253 33469 5279 33521
rect 5201 33457 5331 33469
rect 5253 33405 5279 33457
rect 5201 33393 5331 33405
rect 5253 33341 5279 33393
rect 5201 33329 5331 33341
rect 5253 33277 5279 33329
rect 5201 33264 5331 33277
rect 5253 33212 5279 33264
rect 5201 33199 5331 33212
rect 5253 33147 5279 33199
rect 5201 33134 5331 33147
rect 5253 33082 5279 33134
rect 5201 33069 5331 33082
rect 5253 33017 5279 33069
rect 5201 33004 5331 33017
rect 5253 32952 5279 33004
rect 5201 32939 5331 32952
rect 5253 32887 5279 32939
rect 5201 32874 5331 32887
rect 5253 32822 5279 32874
rect 5201 32809 5331 32822
rect 5253 32757 5279 32809
rect 5201 32744 5331 32757
rect 5253 32692 5279 32744
rect 5201 32679 5331 32692
rect 5253 32627 5279 32679
rect 5201 32614 5331 32627
rect 5253 32562 5279 32614
rect 5201 32549 5331 32562
rect 5253 32497 5279 32549
rect 5201 29625 5331 32497
rect 5253 29573 5279 29625
rect 5201 29561 5331 29573
rect 5253 29509 5279 29561
rect 5201 29497 5331 29509
rect 5253 29445 5279 29497
rect 5201 29433 5331 29445
rect 5253 29381 5279 29433
rect 5201 29369 5331 29381
rect 5253 29317 5279 29369
rect 5201 29305 5331 29317
rect 5253 29253 5279 29305
rect 5201 29241 5331 29253
rect 5253 29189 5279 29241
rect 5201 29177 5331 29189
rect 5253 29125 5279 29177
rect 5201 29113 5331 29125
rect 5253 29061 5279 29113
rect 5201 29049 5331 29061
rect 5253 28997 5279 29049
rect 5201 28985 5331 28997
rect 5253 28933 5279 28985
rect 5201 28921 5331 28933
rect 5253 28869 5279 28921
rect 5201 28857 5331 28869
rect 5253 28805 5279 28857
rect 5201 28793 5331 28805
rect 5253 28741 5279 28793
rect 5201 28729 5331 28741
rect 5253 28677 5279 28729
rect 5201 28664 5331 28677
rect 5253 28612 5279 28664
rect 5201 28599 5331 28612
rect 5253 28547 5279 28599
rect 5201 28534 5331 28547
rect 5253 28482 5279 28534
rect 5201 28469 5331 28482
rect 5253 28417 5279 28469
rect 5201 28404 5331 28417
rect 5253 28352 5279 28404
rect 5201 28339 5331 28352
rect 5253 28287 5279 28339
rect 5201 28274 5331 28287
rect 5253 28222 5279 28274
rect 5201 28209 5331 28222
rect 5253 28157 5279 28209
rect 5201 28144 5331 28157
rect 5253 28092 5279 28144
rect 5201 28079 5331 28092
rect 5253 28027 5279 28079
rect 5201 28014 5331 28027
rect 5253 27962 5279 28014
rect 5201 27949 5331 27962
rect 5253 27897 5279 27949
rect 5201 25025 5331 27897
rect 5253 24973 5279 25025
rect 5201 24961 5331 24973
rect 5253 24909 5279 24961
rect 5201 24897 5331 24909
rect 5253 24845 5279 24897
rect 5201 24833 5331 24845
rect 5253 24781 5279 24833
rect 5201 24769 5331 24781
rect 5253 24717 5279 24769
rect 5201 24705 5331 24717
rect 5253 24653 5279 24705
rect 5201 24641 5331 24653
rect 5253 24589 5279 24641
rect 5201 24577 5331 24589
rect 5253 24525 5279 24577
rect 5201 24513 5331 24525
rect 5253 24461 5279 24513
rect 5201 24449 5331 24461
rect 5253 24397 5279 24449
rect 5201 24385 5331 24397
rect 5253 24333 5279 24385
rect 5201 24321 5331 24333
rect 5253 24269 5279 24321
rect 5201 24257 5331 24269
rect 5253 24205 5279 24257
rect 5201 24193 5331 24205
rect 5253 24141 5279 24193
rect 5201 24129 5331 24141
rect 5253 24077 5279 24129
rect 5201 24064 5331 24077
rect 5253 24012 5279 24064
rect 5201 23999 5331 24012
rect 5253 23947 5279 23999
rect 5201 23934 5331 23947
rect 5253 23882 5279 23934
rect 5201 23869 5331 23882
rect 5253 23817 5279 23869
rect 5201 23804 5331 23817
rect 5253 23752 5279 23804
rect 5201 23739 5331 23752
rect 5253 23687 5279 23739
rect 5201 23674 5331 23687
rect 5253 23622 5279 23674
rect 5201 23609 5331 23622
rect 5253 23557 5279 23609
rect 5201 23544 5331 23557
rect 5253 23492 5279 23544
rect 5201 23479 5331 23492
rect 5253 23427 5279 23479
rect 5201 23414 5331 23427
rect 5253 23362 5279 23414
rect 5201 23349 5331 23362
rect 4359 23265 4365 23299
rect 4399 23265 4437 23299
rect 4471 23265 4477 23299
rect 4359 23226 4477 23265
rect 4359 23192 4365 23226
rect 4399 23192 4437 23226
rect 4471 23192 4477 23226
rect 4359 23153 4477 23192
rect 4359 23119 4365 23153
rect 4399 23119 4437 23153
rect 4471 23119 4477 23153
rect 4359 23080 4477 23119
rect 4359 23046 4365 23080
rect 4399 23046 4437 23080
rect 4471 23046 4477 23080
rect 4359 23007 4477 23046
rect 4359 22973 4365 23007
rect 4399 22973 4437 23007
rect 4471 22973 4477 23007
rect 5253 23297 5279 23349
rect 4359 22934 4477 22973
rect 4359 22900 4365 22934
rect 4399 22900 4437 22934
rect 4471 22900 4477 22934
rect 4359 22861 4477 22900
rect 4777 22995 4841 22999
rect 4777 22943 4783 22995
rect 4835 22943 4841 22995
rect 4777 22931 4841 22943
rect 4777 22879 4783 22931
rect 4835 22879 4841 22931
rect 4359 22827 4365 22861
rect 4399 22827 4437 22861
rect 4471 22827 4477 22861
rect 4359 22788 4477 22827
rect 4359 22754 4365 22788
rect 4399 22754 4437 22788
rect 4471 22754 4477 22788
rect 4359 22715 4477 22754
rect 4359 22681 4365 22715
rect 4399 22681 4437 22715
rect 4471 22681 4477 22715
rect 4359 22642 4477 22681
rect 4359 22608 4365 22642
rect 4399 22608 4437 22642
rect 4471 22608 4477 22642
rect 4359 22569 4477 22608
rect 4359 22535 4365 22569
rect 4399 22535 4437 22569
rect 4471 22535 4477 22569
rect 4359 22496 4477 22535
rect 4359 22462 4365 22496
rect 4399 22462 4437 22496
rect 4471 22462 4477 22496
rect 4359 22423 4477 22462
rect 4359 22389 4365 22423
rect 4399 22389 4437 22423
rect 4471 22389 4477 22423
rect 4359 22350 4477 22389
rect 4359 22316 4365 22350
rect 4399 22316 4437 22350
rect 4471 22316 4477 22350
rect 4359 22277 4477 22316
rect 4359 22243 4365 22277
rect 4399 22243 4437 22277
rect 4471 22243 4477 22277
rect 4359 22204 4477 22243
rect 4359 22170 4365 22204
rect 4399 22170 4437 22204
rect 4471 22170 4477 22204
rect 4359 22131 4477 22170
rect 4359 22097 4365 22131
rect 4399 22097 4437 22131
rect 4471 22097 4477 22131
rect 4359 22058 4477 22097
rect 4359 22024 4365 22058
rect 4399 22024 4437 22058
rect 4471 22024 4477 22058
rect 4359 21985 4477 22024
rect 4359 21951 4365 21985
rect 4399 21951 4437 21985
rect 4471 21951 4477 21985
rect 4359 21912 4477 21951
rect 4359 21878 4365 21912
rect 4399 21878 4437 21912
rect 4471 21878 4477 21912
rect 4359 21839 4477 21878
rect 4359 21805 4365 21839
rect 4399 21805 4437 21839
rect 4471 21805 4477 21839
rect 4359 21766 4477 21805
rect 4359 21732 4365 21766
rect 4399 21732 4437 21766
rect 4471 21732 4477 21766
rect 4359 21693 4477 21732
rect 4359 21659 4365 21693
rect 4399 21659 4437 21693
rect 4471 21659 4477 21693
rect 4359 21620 4477 21659
rect 4359 21586 4365 21620
rect 4399 21586 4437 21620
rect 4471 21586 4477 21620
rect 4359 21547 4477 21586
rect 4359 21513 4365 21547
rect 4399 21513 4437 21547
rect 4471 21513 4477 21547
rect 4359 21474 4477 21513
rect 4359 21440 4365 21474
rect 4399 21440 4437 21474
rect 4471 21440 4477 21474
rect 4359 21401 4477 21440
rect 4359 21367 4365 21401
rect 4399 21367 4437 21401
rect 4471 21367 4477 21401
rect 4359 21328 4477 21367
rect 4359 21294 4365 21328
rect 4399 21294 4437 21328
rect 4471 21294 4477 21328
rect 4359 21255 4477 21294
rect 4359 21221 4365 21255
rect 4399 21221 4437 21255
rect 4471 21221 4477 21255
rect 4359 21182 4477 21221
rect 4359 21148 4365 21182
rect 4399 21148 4437 21182
rect 4471 21148 4477 21182
rect 4359 21109 4477 21148
rect 4359 21075 4365 21109
rect 4399 21075 4437 21109
rect 4471 21075 4477 21109
rect 4359 21036 4477 21075
rect 4359 21002 4365 21036
rect 4399 21002 4437 21036
rect 4471 21002 4477 21036
rect 4359 20963 4477 21002
rect 4359 20929 4365 20963
rect 4399 20929 4437 20963
rect 4471 20929 4477 20963
rect 4359 20890 4477 20929
rect 4359 20856 4365 20890
rect 4399 20856 4437 20890
rect 4471 20856 4477 20890
rect 4359 20817 4477 20856
rect 4359 20783 4365 20817
rect 4399 20783 4437 20817
rect 4471 20783 4477 20817
rect 4359 20744 4477 20783
rect 4359 20710 4365 20744
rect 4399 20710 4437 20744
rect 4471 20710 4477 20744
rect 4359 20671 4477 20710
rect 4359 20637 4365 20671
rect 4399 20637 4437 20671
rect 4471 20637 4477 20671
rect 4359 20598 4477 20637
rect 4359 20564 4365 20598
rect 4399 20564 4437 20598
rect 4471 20564 4477 20598
rect 4359 20525 4477 20564
rect 4359 20491 4365 20525
rect 4399 20491 4437 20525
rect 4471 20491 4477 20525
rect 4359 20452 4477 20491
rect 4359 20418 4365 20452
rect 4399 20418 4437 20452
rect 4471 20418 4477 20452
rect 4359 20379 4477 20418
rect 4359 20345 4365 20379
rect 4399 20345 4437 20379
rect 4471 20345 4477 20379
rect 4359 20306 4477 20345
rect 4359 20272 4365 20306
rect 4399 20272 4437 20306
rect 4471 20272 4477 20306
rect 4359 20233 4477 20272
rect 4359 20199 4365 20233
rect 4399 20199 4437 20233
rect 4471 20199 4477 20233
rect 4359 20160 4477 20199
rect 4359 20126 4365 20160
rect 4399 20126 4437 20160
rect 4471 20126 4477 20160
rect 4359 20087 4477 20126
rect 4359 20053 4365 20087
rect 4399 20053 4437 20087
rect 4471 20053 4477 20087
rect 4359 20014 4477 20053
rect 4359 19980 4365 20014
rect 4399 19980 4437 20014
rect 4471 19980 4477 20014
rect 4359 19941 4477 19980
rect 4359 19907 4365 19941
rect 4399 19907 4437 19941
rect 4471 19907 4477 19941
rect 4359 19868 4477 19907
rect 4359 19834 4365 19868
rect 4399 19834 4437 19868
rect 4471 19834 4477 19868
rect 4359 19795 4477 19834
rect 4359 19761 4365 19795
rect 4399 19761 4437 19795
rect 4471 19761 4477 19795
rect 4359 19722 4477 19761
rect 4359 19688 4365 19722
rect 4399 19688 4437 19722
rect 4471 19688 4477 19722
rect 4359 19649 4477 19688
rect 4359 19615 4365 19649
rect 4399 19615 4437 19649
rect 4471 19615 4477 19649
rect 4359 19576 4477 19615
rect 4359 19542 4365 19576
rect 4399 19542 4437 19576
rect 4471 19542 4477 19576
rect 3907 19391 4059 19500
tri 4352 19523 4359 19530 se
rect 4359 19529 4477 19542
rect 4777 22490 4901 22496
rect 4829 22484 4849 22490
rect 4777 22426 4784 22438
rect 4890 22426 4901 22438
rect 4777 22362 4784 22374
rect 4890 22362 4901 22374
rect 4777 22298 4784 22310
rect 4890 22298 4901 22310
rect 4777 22234 4784 22246
rect 4890 22234 4901 22246
rect 4777 22170 4784 22182
rect 4890 22170 4901 22182
rect 4777 22106 4784 22118
rect 4890 22106 4901 22118
rect 4777 22042 4784 22054
rect 4890 22042 4901 22054
rect 4777 21978 4784 21990
rect 4890 21978 4901 21990
rect 4777 21914 4784 21926
rect 4890 21914 4901 21926
rect 4777 21850 4784 21862
rect 4890 21850 4901 21862
rect 4777 21786 4784 21798
rect 4890 21786 4901 21798
rect 4777 21722 4784 21734
rect 4890 21722 4901 21734
rect 4777 21658 4784 21670
rect 4890 21658 4901 21670
rect 4777 21594 4784 21606
rect 4890 21594 4901 21606
rect 4777 21529 4784 21542
rect 4890 21529 4901 21542
rect 4777 21464 4784 21477
rect 4890 21464 4901 21477
rect 4777 21399 4784 21412
rect 4890 21399 4901 21412
rect 4777 21334 4784 21347
rect 4890 21334 4901 21347
rect 4777 21269 4784 21282
rect 4890 21269 4901 21282
rect 4777 21204 4784 21217
rect 4890 21204 4901 21217
rect 4777 21139 4784 21152
rect 4890 21139 4901 21152
rect 4777 21074 4784 21087
rect 4890 21074 4901 21087
rect 4777 21009 4784 21022
rect 4890 21009 4901 21022
rect 4777 20944 4784 20957
rect 4890 20944 4901 20957
rect 4777 20879 4784 20892
rect 4890 20879 4901 20892
rect 4777 20814 4784 20827
rect 4890 20814 4901 20827
tri 4477 19529 4478 19530 sw
rect 4359 19523 4478 19529
rect 4352 19502 4478 19523
tri 4478 19502 4505 19529 sw
tri 4750 19502 4777 19529 se
rect 4777 19502 4784 20762
rect 4352 19490 4542 19502
tri 4059 19391 4152 19484 sw
rect 3907 19382 4223 19391
tri 3907 19379 3910 19382 ne
rect 3910 19379 4223 19382
tri 3910 19328 3961 19379 ne
rect 3961 19129 3967 19379
rect 3961 19090 4039 19129
rect 3961 19056 3967 19090
rect 4001 19057 4039 19090
rect 4001 19056 4111 19057
rect 3961 19018 4111 19056
rect 3961 19017 4039 19018
rect 3961 18983 3967 19017
rect 4001 18984 4039 19017
rect 4073 18985 4111 19018
rect 4217 18985 4223 19379
rect 4073 18984 4223 18985
rect 4001 18983 4223 18984
rect 3961 18946 4223 18983
rect 3961 18945 4111 18946
rect 3961 18944 4039 18945
rect 3961 18910 3967 18944
rect 4001 18911 4039 18944
rect 4073 18912 4111 18945
rect 4145 18912 4183 18946
rect 4217 18912 4223 18946
rect 4073 18911 4223 18912
rect 4001 18910 4223 18911
rect 3961 18873 4223 18910
rect 3961 18872 4111 18873
rect 3961 18871 4039 18872
rect 3961 18837 3967 18871
rect 4001 18838 4039 18871
rect 4073 18839 4111 18872
rect 4145 18839 4183 18873
rect 4217 18839 4223 18873
rect 4073 18838 4223 18839
rect 4001 18837 4223 18838
rect 3961 18800 4223 18837
rect 3961 18799 4111 18800
rect 3961 18798 4039 18799
rect 3961 18764 3967 18798
rect 4001 18765 4039 18798
rect 4073 18766 4111 18799
rect 4145 18766 4183 18800
rect 4217 18766 4223 18800
rect 4073 18765 4223 18766
rect 4001 18764 4223 18765
rect 3961 18727 4223 18764
rect 3961 18726 4111 18727
rect 3961 18725 4039 18726
rect 3961 18691 3967 18725
rect 4001 18692 4039 18725
rect 4073 18693 4111 18726
rect 4145 18693 4183 18727
rect 4217 18693 4223 18727
rect 4073 18692 4223 18693
rect 4001 18691 4223 18692
rect 3961 18654 4223 18691
rect 3961 18653 4111 18654
rect 3961 18652 4039 18653
rect 3961 18618 3967 18652
rect 4001 18619 4039 18652
rect 4073 18620 4111 18653
rect 4145 18620 4183 18654
rect 4217 18620 4223 18654
rect 4073 18619 4223 18620
rect 4001 18618 4223 18619
rect 3961 18581 4223 18618
rect 3961 18580 4111 18581
rect 3961 18579 4039 18580
rect 3961 18545 3967 18579
rect 4001 18546 4039 18579
rect 4073 18547 4111 18580
rect 4145 18547 4183 18581
rect 4217 18547 4223 18581
rect 4073 18546 4223 18547
rect 4001 18545 4223 18546
rect 3961 18508 4223 18545
rect 3961 18507 4111 18508
rect 3961 18506 4039 18507
rect 3961 18472 3967 18506
rect 4001 18473 4039 18506
rect 4073 18474 4111 18507
rect 4145 18474 4183 18508
rect 4217 18474 4223 18508
rect 4073 18473 4223 18474
rect 4001 18472 4223 18473
rect 3961 18435 4223 18472
rect 3961 18434 4111 18435
rect 3961 18433 4039 18434
rect 3961 18399 3967 18433
rect 4001 18400 4039 18433
rect 4073 18401 4111 18434
rect 4145 18401 4183 18435
rect 4217 18401 4223 18435
rect 4073 18400 4223 18401
rect 4001 18399 4223 18400
rect 3961 18362 4223 18399
rect 3961 18361 4111 18362
rect 3961 18360 4039 18361
rect 3961 18326 3967 18360
rect 4001 18327 4039 18360
rect 4073 18328 4111 18361
rect 4145 18328 4183 18362
rect 4217 18328 4223 18362
rect 4073 18327 4223 18328
rect 4001 18326 4223 18327
rect 3961 18289 4223 18326
rect 3961 18288 4111 18289
rect 3961 18287 4039 18288
rect 3961 18253 3967 18287
rect 4001 18254 4039 18287
rect 4073 18255 4111 18288
rect 4145 18255 4183 18289
rect 4217 18255 4223 18289
rect 4073 18254 4223 18255
rect 4001 18253 4223 18254
rect 3961 18216 4223 18253
rect 3961 18215 4111 18216
rect 3961 18214 4039 18215
rect 3961 18180 3967 18214
rect 4001 18181 4039 18214
rect 4073 18182 4111 18215
rect 4145 18182 4183 18216
rect 4217 18182 4223 18216
rect 4073 18181 4223 18182
rect 4001 18180 4223 18181
rect 3961 18143 4223 18180
rect 3961 18142 4111 18143
rect 3961 18141 4039 18142
rect 3961 18107 3967 18141
rect 4001 18108 4039 18141
rect 4073 18109 4111 18142
rect 4145 18109 4183 18143
rect 4217 18109 4223 18143
rect 4073 18108 4223 18109
rect 4001 18107 4223 18108
rect 3961 18070 4223 18107
rect 3961 18069 4111 18070
rect 3961 18068 4039 18069
rect 3961 18034 3967 18068
rect 4001 18035 4039 18068
rect 4073 18036 4111 18069
rect 4145 18036 4183 18070
rect 4217 18036 4223 18070
rect 4073 18035 4223 18036
rect 4001 18034 4223 18035
rect 3961 17997 4223 18034
rect 3961 17996 4111 17997
rect 3961 17995 4039 17996
rect 3961 17961 3967 17995
rect 4001 17962 4039 17995
rect 4073 17963 4111 17996
rect 4145 17963 4183 17997
rect 4217 17963 4223 17997
rect 4073 17962 4223 17963
rect 4001 17961 4223 17962
rect 3961 17924 4223 17961
rect 3961 17923 4111 17924
rect 3961 17922 4039 17923
rect 3961 17888 3967 17922
rect 4001 17889 4039 17922
rect 4073 17890 4111 17923
rect 4145 17890 4183 17924
rect 4217 17890 4223 17924
rect 4073 17889 4223 17890
rect 4001 17888 4223 17889
rect 3961 17851 4223 17888
rect 3961 17850 4111 17851
rect 3961 17849 4039 17850
rect 3961 17815 3967 17849
rect 4001 17816 4039 17849
rect 4073 17817 4111 17850
rect 4145 17817 4183 17851
rect 4217 17817 4223 17851
rect 4073 17816 4223 17817
rect 4001 17815 4223 17816
rect 3961 17778 4223 17815
rect 3961 17777 4111 17778
rect 3961 17776 4039 17777
rect 3961 17742 3967 17776
rect 4001 17743 4039 17776
rect 4073 17744 4111 17777
rect 4145 17744 4183 17778
rect 4217 17744 4223 17778
rect 4073 17743 4223 17744
rect 4001 17742 4223 17743
rect 3961 17705 4223 17742
rect 3961 17704 4111 17705
rect 3961 17703 4039 17704
rect 3961 17669 3967 17703
rect 4001 17670 4039 17703
rect 4073 17671 4111 17704
rect 4145 17671 4183 17705
rect 4217 17671 4223 17705
rect 4073 17670 4223 17671
rect 4001 17669 4223 17670
rect 3961 17632 4223 17669
rect 3961 17631 4111 17632
rect 3961 17630 4039 17631
rect 3961 17596 3967 17630
rect 4001 17597 4039 17630
rect 4073 17598 4111 17631
rect 4145 17598 4183 17632
rect 4217 17598 4223 17632
rect 4073 17597 4223 17598
rect 4001 17596 4223 17597
rect 3961 17559 4223 17596
rect 3961 17558 4111 17559
rect 3961 17557 4039 17558
rect 3961 17523 3967 17557
rect 4001 17524 4039 17557
rect 4073 17525 4111 17558
rect 4145 17525 4183 17559
rect 4217 17525 4223 17559
rect 4073 17524 4223 17525
rect 4001 17523 4223 17524
rect 3961 17486 4223 17523
rect 3961 17485 4111 17486
rect 3961 17484 4039 17485
rect 3961 17450 3967 17484
rect 4001 17451 4039 17484
rect 4073 17452 4111 17485
rect 4145 17452 4183 17486
rect 4217 17452 4223 17486
rect 4073 17451 4223 17452
rect 4001 17450 4223 17451
rect 3961 17413 4223 17450
rect 3961 17412 4111 17413
rect 3961 17411 4039 17412
rect 3961 17377 3967 17411
rect 4001 17378 4039 17411
rect 4073 17379 4111 17412
rect 4145 17379 4183 17413
rect 4217 17379 4223 17413
rect 4073 17378 4223 17379
rect 4001 17377 4223 17378
rect 3961 17340 4223 17377
rect 3961 17339 4111 17340
rect 3961 17338 4039 17339
rect 3961 17304 3967 17338
rect 4001 17305 4039 17338
rect 4073 17306 4111 17339
rect 4145 17306 4183 17340
rect 4217 17306 4223 17340
rect 4073 17305 4223 17306
rect 4001 17304 4223 17305
rect 3961 17267 4223 17304
rect 3961 17266 4111 17267
rect 3961 17265 4039 17266
rect 3961 17231 3967 17265
rect 4001 17232 4039 17265
rect 4073 17233 4111 17266
rect 4145 17233 4183 17267
rect 4217 17233 4223 17267
rect 4073 17232 4223 17233
rect 4001 17231 4223 17232
rect 3961 17194 4223 17231
rect 3961 17193 4111 17194
rect 3961 17192 4039 17193
rect 3961 17158 3967 17192
rect 4001 17159 4039 17192
rect 4073 17160 4111 17193
rect 4145 17160 4183 17194
rect 4217 17160 4223 17194
rect 4073 17159 4223 17160
rect 4001 17158 4223 17159
rect 3961 17121 4223 17158
rect 3961 17120 4111 17121
rect 3961 17119 4039 17120
rect 3961 17085 3967 17119
rect 4001 17086 4039 17119
rect 4073 17087 4111 17120
rect 4145 17087 4183 17121
rect 4217 17087 4223 17121
rect 4073 17086 4223 17087
rect 4001 17085 4223 17086
rect 3961 17048 4223 17085
rect 3961 17047 4111 17048
rect 3961 17046 4039 17047
rect 3961 17012 3967 17046
rect 4001 17013 4039 17046
rect 4073 17014 4111 17047
rect 4145 17014 4183 17048
rect 4217 17014 4223 17048
rect 4073 17013 4223 17014
rect 4001 17012 4223 17013
rect 3961 16975 4223 17012
rect 3961 16974 4111 16975
rect 3961 16973 4039 16974
rect 3961 16939 3967 16973
rect 4001 16940 4039 16973
rect 4073 16941 4111 16974
rect 4145 16941 4183 16975
rect 4217 16941 4223 16975
rect 4073 16940 4223 16941
rect 4001 16939 4223 16940
rect 3961 16902 4223 16939
rect 3961 16901 4111 16902
rect 3961 16900 4039 16901
rect 3961 16866 3967 16900
rect 4001 16867 4039 16900
rect 4073 16868 4111 16901
rect 4145 16868 4183 16902
rect 4217 16868 4223 16902
rect 4073 16867 4223 16868
rect 4001 16866 4223 16867
rect 3961 16829 4223 16866
rect 3961 16828 4111 16829
rect 3961 16827 4039 16828
rect 3961 16793 3967 16827
rect 4001 16794 4039 16827
rect 4073 16795 4111 16828
rect 4145 16795 4183 16829
rect 4217 16795 4223 16829
rect 4073 16794 4223 16795
rect 4001 16793 4223 16794
rect 3961 16756 4223 16793
rect 3961 16755 4111 16756
rect 3961 16754 4039 16755
rect 3961 16720 3967 16754
rect 4001 16721 4039 16754
rect 4073 16722 4111 16755
rect 4145 16722 4183 16756
rect 4217 16722 4223 16756
rect 4073 16721 4223 16722
rect 4001 16720 4223 16721
rect 3961 16683 4223 16720
rect 3961 16682 4111 16683
rect 3961 16681 4039 16682
rect 3961 16647 3967 16681
rect 4001 16648 4039 16681
rect 4073 16649 4111 16682
rect 4145 16649 4183 16683
rect 4217 16649 4223 16683
rect 4073 16648 4223 16649
rect 4001 16647 4223 16648
rect 3961 16610 4223 16647
rect 3961 16609 4111 16610
rect 3961 16608 4039 16609
rect 3961 16574 3967 16608
rect 4001 16575 4039 16608
rect 4073 16576 4111 16609
rect 4145 16576 4183 16610
rect 4217 16576 4223 16610
rect 4073 16575 4223 16576
rect 4001 16574 4223 16575
rect 3961 16537 4223 16574
rect 3961 16536 4111 16537
rect 3961 16535 4039 16536
rect 3961 16501 3967 16535
rect 4001 16502 4039 16535
rect 4073 16503 4111 16536
rect 4145 16503 4183 16537
rect 4217 16503 4223 16537
rect 4073 16502 4223 16503
rect 4001 16501 4223 16502
rect 3961 16464 4223 16501
rect 3961 16463 4111 16464
rect 3961 16462 4039 16463
rect 3961 16428 3967 16462
rect 4001 16429 4039 16462
rect 4073 16430 4111 16463
rect 4145 16430 4183 16464
rect 4217 16430 4223 16464
rect 4073 16429 4223 16430
rect 4001 16428 4223 16429
rect 3961 16391 4223 16428
rect 3961 16390 4111 16391
rect 3961 16389 4039 16390
rect 3961 16355 3967 16389
rect 4001 16356 4039 16389
rect 4073 16357 4111 16390
rect 4145 16357 4183 16391
rect 4217 16357 4223 16391
rect 4073 16356 4223 16357
rect 4001 16355 4223 16356
rect 3961 16318 4223 16355
rect 3961 16317 4111 16318
rect 3961 16316 4039 16317
rect 3961 16282 3967 16316
rect 4001 16283 4039 16316
rect 4073 16284 4111 16317
rect 4145 16284 4183 16318
rect 4217 16284 4223 16318
rect 4073 16283 4223 16284
rect 4001 16282 4223 16283
rect 3961 16245 4223 16282
rect 3961 16244 4111 16245
rect 3961 16243 4039 16244
rect 3961 16209 3967 16243
rect 4001 16210 4039 16243
rect 4073 16211 4111 16244
rect 4145 16211 4183 16245
rect 4217 16211 4223 16245
rect 4073 16210 4223 16211
rect 4001 16209 4223 16210
rect 3961 16172 4223 16209
rect 3961 16171 4111 16172
rect 3961 16170 4039 16171
rect 3961 16136 3967 16170
rect 4001 16137 4039 16170
rect 4073 16138 4111 16171
rect 4145 16138 4183 16172
rect 4217 16138 4223 16172
rect 4073 16137 4223 16138
rect 4001 16136 4223 16137
rect 3961 16099 4223 16136
rect 3961 16098 4111 16099
rect 3961 16097 4039 16098
rect 3961 16063 3967 16097
rect 4001 16064 4039 16097
rect 4073 16065 4111 16098
rect 4145 16065 4183 16099
rect 4217 16065 4223 16099
rect 4073 16064 4223 16065
rect 4001 16063 4223 16064
rect 3961 16026 4223 16063
rect 3961 16025 4111 16026
rect 3961 16024 4039 16025
rect 3961 15990 3967 16024
rect 4001 15991 4039 16024
rect 4073 15992 4111 16025
rect 4145 15992 4183 16026
rect 4217 15992 4223 16026
rect 4073 15991 4223 15992
rect 4001 15990 4223 15991
rect 3961 15953 4223 15990
rect 3961 15952 4111 15953
rect 3961 15951 4039 15952
rect 3961 15917 3967 15951
rect 4001 15918 4039 15951
rect 4073 15919 4111 15952
rect 4145 15919 4183 15953
rect 4217 15919 4223 15953
rect 4073 15918 4223 15919
rect 4001 15917 4223 15918
rect 3961 15880 4223 15917
rect 3961 15879 4111 15880
rect 3961 15878 4039 15879
rect 3961 15844 3967 15878
rect 4001 15845 4039 15878
rect 4073 15846 4111 15879
rect 4145 15846 4183 15880
rect 4217 15846 4223 15880
rect 4073 15845 4223 15846
rect 4001 15844 4223 15845
rect 3961 15807 4223 15844
rect 3961 15806 4111 15807
rect 3961 15805 4039 15806
rect 3961 15771 3967 15805
rect 4001 15772 4039 15805
rect 4073 15773 4111 15806
rect 4145 15773 4183 15807
rect 4217 15773 4223 15807
rect 4073 15772 4223 15773
rect 4001 15771 4223 15772
rect 3961 15734 4223 15771
rect 3961 15733 4111 15734
rect 3961 15732 4039 15733
rect 3961 15698 3967 15732
rect 4001 15699 4039 15732
rect 4073 15700 4111 15733
rect 4145 15700 4183 15734
rect 4217 15700 4223 15734
rect 4073 15699 4223 15700
rect 4001 15698 4223 15699
rect 3961 15661 4223 15698
rect 3961 15660 4111 15661
rect 3961 15659 4039 15660
rect 3961 15625 3967 15659
rect 4001 15626 4039 15659
rect 4073 15627 4111 15660
rect 4145 15627 4183 15661
rect 4217 15627 4223 15661
rect 4073 15626 4223 15627
rect 4001 15625 4223 15626
rect 3961 15588 4223 15625
rect 3961 15587 4111 15588
rect 3961 15586 4039 15587
rect 3961 15552 3967 15586
rect 4001 15553 4039 15586
rect 4073 15554 4111 15587
rect 4145 15554 4183 15588
rect 4217 15554 4223 15588
rect 4073 15553 4223 15554
rect 4001 15552 4223 15553
rect 3961 15515 4223 15552
rect 3961 15514 4111 15515
rect 3961 15513 4039 15514
rect 3961 15479 3967 15513
rect 4001 15480 4039 15513
rect 4073 15481 4111 15514
rect 4145 15481 4183 15515
rect 4217 15481 4223 15515
rect 4073 15480 4223 15481
rect 4001 15479 4223 15480
rect 3961 15442 4223 15479
rect 3961 15441 4111 15442
rect 3961 15440 4039 15441
rect 3961 15406 3967 15440
rect 4001 15407 4039 15440
rect 4073 15408 4111 15441
rect 4145 15408 4183 15442
rect 4217 15408 4223 15442
rect 4073 15407 4223 15408
rect 4001 15406 4223 15407
rect 3961 15369 4223 15406
rect 3961 15368 4111 15369
rect 3961 15367 4039 15368
rect 3961 15333 3967 15367
rect 4001 15334 4039 15367
rect 4073 15335 4111 15368
rect 4145 15335 4183 15369
rect 4217 15335 4223 15369
rect 4073 15334 4223 15335
rect 4001 15333 4223 15334
rect 3961 15296 4223 15333
rect 3961 15295 4111 15296
rect 3961 15294 4039 15295
rect 3961 15260 3967 15294
rect 4001 15261 4039 15294
rect 4073 15262 4111 15295
rect 4145 15262 4183 15296
rect 4217 15262 4223 15296
rect 4073 15261 4223 15262
rect 4001 15260 4223 15261
rect 3961 15223 4223 15260
rect 3961 15222 4111 15223
rect 3961 15221 4039 15222
rect 3961 15187 3967 15221
rect 4001 15188 4039 15221
rect 4073 15189 4111 15222
rect 4145 15189 4183 15223
rect 4217 15189 4223 15223
rect 4073 15188 4223 15189
rect 4001 15187 4223 15188
rect 3961 15150 4223 15187
rect 3961 15149 4111 15150
rect 3961 15148 4039 15149
rect 3961 15114 3967 15148
rect 4001 15115 4039 15148
rect 4073 15116 4111 15149
rect 4145 15116 4183 15150
rect 4217 15116 4223 15150
rect 4073 15115 4223 15116
rect 4001 15114 4223 15115
rect 3961 15077 4223 15114
rect 3961 15076 4111 15077
rect 3961 15075 4039 15076
rect 3961 15041 3967 15075
rect 4001 15042 4039 15075
rect 4073 15043 4111 15076
rect 4145 15043 4183 15077
rect 4217 15043 4223 15077
rect 4073 15042 4223 15043
rect 4001 15041 4223 15042
rect 3961 15004 4223 15041
rect 3961 15003 4111 15004
rect 3961 15002 4039 15003
rect 3961 14968 3967 15002
rect 4001 14969 4039 15002
rect 4073 14970 4111 15003
rect 4145 14970 4183 15004
rect 4217 14970 4223 15004
rect 4073 14969 4223 14970
rect 4001 14968 4223 14969
rect 3961 14931 4223 14968
rect 3961 14930 4111 14931
rect 3961 14929 4039 14930
rect 3961 14895 3967 14929
rect 4001 14896 4039 14929
rect 4073 14897 4111 14930
rect 4145 14897 4183 14931
rect 4217 14897 4223 14931
rect 4073 14896 4223 14897
rect 4001 14895 4223 14896
rect 3682 14831 3688 14883
rect 3740 14831 3754 14883
rect 3806 14831 3812 14883
rect 3961 14858 4223 14895
rect 3961 14857 4111 14858
rect 3961 14856 4039 14857
tri 3407 14730 3426 14749 se
rect 3426 14730 3521 14749
rect 1635 14702 3521 14730
rect 3961 14822 3967 14856
rect 4001 14823 4039 14856
rect 4073 14824 4111 14857
rect 4145 14824 4183 14858
rect 4217 14824 4223 14858
rect 4073 14823 4223 14824
rect 4001 14822 4223 14823
rect 3961 14785 4223 14822
rect 3961 14784 4111 14785
rect 3961 14783 4039 14784
rect 3961 14749 3967 14783
rect 4001 14750 4039 14783
rect 4073 14751 4111 14784
rect 4145 14751 4183 14785
rect 4217 14751 4223 14785
rect 4073 14750 4223 14751
rect 4001 14749 4223 14750
rect 3961 14712 4223 14749
tri 3960 14711 3961 14712 se
rect 3961 14711 4111 14712
tri 3959 14710 3960 14711 se
rect 3960 14710 4039 14711
rect 1635 14650 3359 14702
rect 3411 14650 3448 14702
rect 3500 14650 3521 14702
tri 3925 14676 3959 14710 se
rect 3959 14676 3967 14710
rect 4001 14677 4039 14710
rect 4073 14678 4111 14711
rect 4145 14678 4183 14712
rect 4217 14678 4223 14712
rect 4073 14677 4223 14678
rect 4001 14676 4223 14677
tri 3899 14650 3925 14676 se
rect 3925 14650 4223 14676
rect 1635 14648 1747 14650
tri 1747 14648 1749 14650 nw
tri 3897 14648 3899 14650 se
rect 3899 14648 4223 14650
rect 1635 14639 1738 14648
tri 1738 14639 1747 14648 nw
tri 3888 14639 3897 14648 se
rect 3897 14639 4223 14648
rect 1635 14638 1737 14639
tri 1737 14638 1738 14639 nw
tri 3887 14638 3888 14639 se
rect 3888 14638 4111 14639
rect 1635 14637 1736 14638
tri 1736 14637 1737 14638 nw
tri 3886 14637 3887 14638 se
rect 3887 14637 4039 14638
tri 1608 8880 1635 8907 se
rect 1635 8880 1715 14637
tri 1715 14616 1736 14637 nw
tri 3865 14616 3886 14637 se
rect 3886 14616 3967 14637
tri 3852 14603 3865 14616 se
rect 3865 14603 3967 14616
rect 4001 14604 4039 14637
rect 4073 14605 4111 14638
rect 4145 14605 4183 14639
rect 4217 14605 4223 14639
rect 4073 14604 4223 14605
rect 4001 14603 4223 14604
tri 3826 14577 3852 14603 se
rect 3852 14577 4223 14603
tri 3824 14575 3826 14577 se
rect 3826 14575 4223 14577
tri 3819 14570 3824 14575 se
rect 3824 14570 4223 14575
tri 1587 8859 1608 8880 se
rect 1608 8859 1715 8880
rect 222 8728 229 8762
rect 263 8728 270 8762
rect 222 8690 270 8728
rect 222 8656 229 8690
rect 263 8656 270 8690
rect 222 8644 270 8656
rect 357 8779 1715 8859
rect 1821 14566 4223 14570
rect 1821 14565 4111 14566
rect 1821 14564 4039 14565
rect 1821 14530 1899 14564
rect 1933 14530 1973 14564
rect 2007 14530 2047 14564
rect 2081 14530 2121 14564
rect 2155 14530 2195 14564
rect 2229 14530 2269 14564
rect 2303 14530 2343 14564
rect 2377 14530 2417 14564
rect 2451 14530 2491 14564
rect 2525 14530 2565 14564
rect 2599 14530 2639 14564
rect 2673 14530 2713 14564
rect 2747 14530 2787 14564
rect 2821 14530 2861 14564
rect 2895 14530 2935 14564
rect 2969 14530 3009 14564
rect 3043 14530 3083 14564
rect 3117 14530 3157 14564
rect 3191 14530 3231 14564
rect 3265 14530 3305 14564
rect 3339 14530 3379 14564
rect 3413 14530 3453 14564
rect 3487 14530 3527 14564
rect 3561 14530 3601 14564
rect 3635 14530 3675 14564
rect 3709 14530 3748 14564
rect 3782 14530 3821 14564
rect 3855 14530 3894 14564
rect 3928 14530 3967 14564
rect 4001 14531 4039 14564
rect 4073 14532 4111 14565
rect 4145 14532 4183 14566
rect 4217 14532 4223 14566
rect 4073 14531 4223 14532
rect 4001 14530 4223 14531
rect 1821 14493 4223 14530
rect 1821 14492 4111 14493
rect 1821 13882 1827 14492
rect 1933 14458 1973 14492
rect 2007 14458 2047 14492
rect 2081 14458 2121 14492
rect 2155 14458 2195 14492
rect 2229 14458 2269 14492
rect 2303 14458 2343 14492
rect 2377 14458 2417 14492
rect 2451 14458 2491 14492
rect 2525 14458 2565 14492
rect 2599 14458 2639 14492
rect 2673 14458 2713 14492
rect 2747 14458 2787 14492
rect 2821 14458 2861 14492
rect 2895 14458 2935 14492
rect 2969 14458 3009 14492
rect 3043 14458 3083 14492
rect 3117 14458 3157 14492
rect 3191 14458 3231 14492
rect 3265 14458 3305 14492
rect 3339 14458 3379 14492
rect 3413 14458 3453 14492
rect 3487 14458 3527 14492
rect 3561 14458 3601 14492
rect 3635 14458 3674 14492
rect 3708 14458 3747 14492
rect 3781 14458 3820 14492
rect 3854 14458 3893 14492
rect 3927 14458 3966 14492
rect 4000 14458 4039 14492
rect 4073 14459 4111 14492
rect 4145 14459 4183 14493
rect 4217 14459 4223 14493
rect 4073 14458 4223 14459
rect 1933 14420 4223 14458
rect 2005 14386 2045 14420
rect 2079 14386 2119 14420
rect 2153 14386 2193 14420
rect 2227 14386 2267 14420
rect 2301 14386 2341 14420
rect 2375 14386 2415 14420
rect 2449 14386 2489 14420
rect 2523 14386 2563 14420
rect 2597 14386 2637 14420
rect 2671 14386 2711 14420
rect 2745 14386 2785 14420
rect 2819 14386 2859 14420
rect 2893 14386 2933 14420
rect 2967 14386 3007 14420
rect 3041 14386 3081 14420
rect 3115 14386 3155 14420
rect 3189 14386 3229 14420
rect 3263 14386 3303 14420
rect 3337 14386 3377 14420
rect 3411 14386 3451 14420
rect 3485 14386 3525 14420
rect 3559 14386 3599 14420
rect 3633 14386 3672 14420
rect 3706 14386 3745 14420
rect 3779 14386 3818 14420
rect 3852 14386 3891 14420
rect 3925 14386 3964 14420
rect 3998 14386 4037 14420
rect 4071 14386 4111 14420
rect 4145 14386 4183 14420
rect 4217 14386 4223 14420
rect 2005 14348 4223 14386
rect 2077 14314 2117 14348
rect 2151 14314 2191 14348
rect 2225 14314 2265 14348
rect 2299 14314 2339 14348
rect 2373 14314 2413 14348
rect 2447 14314 2487 14348
rect 2521 14314 2561 14348
rect 2595 14314 2635 14348
rect 2669 14314 2709 14348
rect 2743 14314 2783 14348
rect 2817 14314 2857 14348
rect 2891 14314 2931 14348
rect 2965 14314 3005 14348
rect 3039 14314 3079 14348
rect 3113 14314 3153 14348
rect 3187 14314 3227 14348
rect 3261 14314 3301 14348
rect 3335 14314 3375 14348
rect 3409 14314 3449 14348
rect 3483 14314 3523 14348
rect 3557 14314 3597 14348
rect 3631 14314 3671 14348
rect 3705 14314 3745 14348
rect 3779 14314 3818 14348
rect 3852 14314 3891 14348
rect 3925 14314 3964 14348
rect 3998 14314 4037 14348
rect 4071 14314 4110 14348
rect 4144 14314 4223 14348
rect 2077 14308 4223 14314
rect 4352 18592 4358 19490
rect 4352 18553 4430 18592
rect 4352 18519 4358 18553
rect 4392 18520 4430 18553
rect 4536 18520 4542 19490
tri 4714 19466 4750 19502 se
rect 4750 19466 4784 19502
rect 4711 18922 4784 19466
rect 4890 18922 4901 20762
rect 4711 18883 4901 18922
rect 4711 18849 4784 18883
rect 4818 18849 4856 18883
rect 4890 18849 4901 18883
rect 4711 18810 4901 18849
rect 4711 18776 4784 18810
rect 4818 18776 4856 18810
rect 4890 18776 4901 18810
rect 4711 18737 4901 18776
rect 4711 18703 4784 18737
rect 4818 18703 4856 18737
rect 4890 18703 4901 18737
rect 4392 18519 4542 18520
rect 4352 18481 4542 18519
rect 4352 18480 4430 18481
rect 4352 18446 4358 18480
rect 4392 18447 4430 18480
rect 4464 18447 4502 18481
rect 4536 18447 4542 18481
rect 4392 18446 4542 18447
rect 4352 18408 4542 18446
rect 4352 18407 4430 18408
rect 4352 18373 4358 18407
rect 4392 18374 4430 18407
rect 4464 18374 4502 18408
rect 4536 18374 4542 18408
rect 4392 18373 4542 18374
rect 4352 18335 4542 18373
rect 4352 18334 4430 18335
rect 4352 18300 4358 18334
rect 4392 18301 4430 18334
rect 4464 18301 4502 18335
rect 4536 18301 4542 18335
rect 4392 18300 4542 18301
rect 4352 18262 4542 18300
rect 4352 18261 4430 18262
rect 4352 18227 4358 18261
rect 4392 18228 4430 18261
rect 4464 18228 4502 18262
rect 4536 18228 4542 18262
rect 4392 18227 4542 18228
rect 4352 18189 4542 18227
rect 4352 18188 4430 18189
rect 4352 18154 4358 18188
rect 4392 18155 4430 18188
rect 4464 18155 4502 18189
rect 4536 18155 4542 18189
rect 4392 18154 4542 18155
rect 4352 18116 4542 18154
rect 4352 18115 4430 18116
rect 4352 18081 4358 18115
rect 4392 18082 4430 18115
rect 4464 18082 4502 18116
rect 4536 18082 4542 18116
rect 4392 18081 4542 18082
rect 4352 18043 4542 18081
rect 4352 18042 4430 18043
rect 4352 18008 4358 18042
rect 4392 18009 4430 18042
rect 4464 18009 4502 18043
rect 4536 18009 4542 18043
rect 4392 18008 4542 18009
rect 4352 17970 4542 18008
rect 4352 17969 4430 17970
rect 4352 17935 4358 17969
rect 4392 17936 4430 17969
rect 4464 17936 4502 17970
rect 4536 17936 4542 17970
rect 4392 17935 4542 17936
rect 4352 17897 4542 17935
rect 4352 17896 4430 17897
rect 4352 17862 4358 17896
rect 4392 17863 4430 17896
rect 4464 17863 4502 17897
rect 4536 17863 4542 17897
rect 4392 17862 4542 17863
rect 4352 17824 4542 17862
rect 4352 17823 4430 17824
rect 4352 17789 4358 17823
rect 4392 17790 4430 17823
rect 4464 17790 4502 17824
rect 4536 17790 4542 17824
rect 4392 17789 4542 17790
rect 4352 17751 4542 17789
rect 4352 17750 4430 17751
rect 4352 17716 4358 17750
rect 4392 17717 4430 17750
rect 4464 17717 4502 17751
rect 4536 17717 4542 17751
rect 4392 17716 4542 17717
rect 4352 17678 4542 17716
rect 4352 17677 4430 17678
rect 4352 17643 4358 17677
rect 4392 17644 4430 17677
rect 4464 17644 4502 17678
rect 4536 17644 4542 17678
rect 4392 17643 4542 17644
rect 4352 17605 4542 17643
rect 4352 17604 4430 17605
rect 4352 17570 4358 17604
rect 4392 17571 4430 17604
rect 4464 17571 4502 17605
rect 4536 17571 4542 17605
rect 4392 17570 4542 17571
rect 4352 17532 4542 17570
rect 4352 17531 4430 17532
rect 4352 17497 4358 17531
rect 4392 17498 4430 17531
rect 4464 17498 4502 17532
rect 4536 17498 4542 17532
rect 4392 17497 4542 17498
rect 4352 17459 4542 17497
rect 4352 17458 4430 17459
rect 4352 17424 4358 17458
rect 4392 17425 4430 17458
rect 4464 17425 4502 17459
rect 4536 17425 4542 17459
rect 4392 17424 4542 17425
rect 4352 17386 4542 17424
rect 4352 17385 4430 17386
rect 4352 17351 4358 17385
rect 4392 17352 4430 17385
rect 4464 17352 4502 17386
rect 4536 17352 4542 17386
rect 4392 17351 4542 17352
rect 4352 17313 4542 17351
rect 4352 17312 4430 17313
rect 4352 17278 4358 17312
rect 4392 17279 4430 17312
rect 4464 17279 4502 17313
rect 4536 17279 4542 17313
rect 4392 17278 4542 17279
rect 4352 17240 4542 17278
rect 4352 17239 4430 17240
rect 4352 17205 4358 17239
rect 4392 17206 4430 17239
rect 4464 17206 4502 17240
rect 4536 17206 4542 17240
rect 4392 17205 4542 17206
rect 4352 17167 4542 17205
rect 4352 17166 4430 17167
rect 4352 17132 4358 17166
rect 4392 17133 4430 17166
rect 4464 17133 4502 17167
rect 4536 17133 4542 17167
rect 4392 17132 4542 17133
rect 4352 17094 4542 17132
rect 4352 17093 4430 17094
rect 4352 17059 4358 17093
rect 4392 17060 4430 17093
rect 4464 17060 4502 17094
rect 4536 17060 4542 17094
rect 4392 17059 4542 17060
rect 4352 17021 4542 17059
rect 4352 17020 4430 17021
rect 4352 16986 4358 17020
rect 4392 16987 4430 17020
rect 4464 16987 4502 17021
rect 4536 16987 4542 17021
rect 4392 16986 4542 16987
rect 4352 16948 4542 16986
rect 4352 16947 4430 16948
rect 4352 16913 4358 16947
rect 4392 16914 4430 16947
rect 4464 16914 4502 16948
rect 4536 16914 4542 16948
rect 4392 16913 4542 16914
rect 4352 16875 4542 16913
rect 4352 16874 4430 16875
rect 4352 16840 4358 16874
rect 4392 16841 4430 16874
rect 4464 16841 4502 16875
rect 4536 16841 4542 16875
rect 4392 16840 4542 16841
rect 4352 16802 4542 16840
rect 4352 16801 4430 16802
rect 4352 16767 4358 16801
rect 4392 16768 4430 16801
rect 4464 16768 4502 16802
rect 4536 16768 4542 16802
rect 4392 16767 4542 16768
rect 4352 16729 4542 16767
rect 4352 16728 4430 16729
rect 4352 16694 4358 16728
rect 4392 16695 4430 16728
rect 4464 16695 4502 16729
rect 4536 16695 4542 16729
rect 4392 16694 4542 16695
rect 4352 16656 4542 16694
rect 4352 16655 4430 16656
rect 4352 16621 4358 16655
rect 4392 16622 4430 16655
rect 4464 16622 4502 16656
rect 4536 16622 4542 16656
rect 4392 16621 4542 16622
rect 4352 16583 4542 16621
rect 4352 16582 4430 16583
rect 4352 16548 4358 16582
rect 4392 16549 4430 16582
rect 4464 16549 4502 16583
rect 4536 16549 4542 16583
rect 4392 16548 4542 16549
rect 4352 16510 4542 16548
rect 4352 16509 4430 16510
rect 4352 16475 4358 16509
rect 4392 16476 4430 16509
rect 4464 16476 4502 16510
rect 4536 16476 4542 16510
rect 4392 16475 4542 16476
rect 4352 16437 4542 16475
rect 4352 16436 4430 16437
rect 4352 16402 4358 16436
rect 4392 16403 4430 16436
rect 4464 16403 4502 16437
rect 4536 16403 4542 16437
rect 4392 16402 4542 16403
rect 4352 16364 4542 16402
rect 4352 16363 4430 16364
rect 4352 16329 4358 16363
rect 4392 16330 4430 16363
rect 4464 16330 4502 16364
rect 4536 16330 4542 16364
rect 4392 16329 4542 16330
rect 4352 16291 4542 16329
rect 4352 16290 4430 16291
rect 4352 16256 4358 16290
rect 4392 16257 4430 16290
rect 4464 16257 4502 16291
rect 4536 16257 4542 16291
rect 4392 16256 4542 16257
rect 4352 16218 4542 16256
rect 4352 16217 4430 16218
rect 4352 16183 4358 16217
rect 4392 16184 4430 16217
rect 4464 16184 4502 16218
rect 4536 16184 4542 16218
rect 4392 16183 4542 16184
rect 4352 16145 4542 16183
rect 4352 16144 4430 16145
rect 4352 16110 4358 16144
rect 4392 16111 4430 16144
rect 4464 16111 4502 16145
rect 4536 16111 4542 16145
rect 4392 16110 4542 16111
rect 4352 16072 4542 16110
rect 4352 16071 4430 16072
rect 4352 16037 4358 16071
rect 4392 16038 4430 16071
rect 4464 16038 4502 16072
rect 4536 16038 4542 16072
rect 4392 16037 4542 16038
rect 4352 15999 4542 16037
rect 4352 15998 4430 15999
rect 4352 15964 4358 15998
rect 4392 15965 4430 15998
rect 4464 15965 4502 15999
rect 4536 15965 4542 15999
rect 4392 15964 4542 15965
rect 4352 15926 4542 15964
rect 4352 15925 4430 15926
rect 4352 15891 4358 15925
rect 4392 15892 4430 15925
rect 4464 15892 4502 15926
rect 4536 15892 4542 15926
rect 4392 15891 4542 15892
rect 4352 15853 4542 15891
rect 4352 15852 4430 15853
rect 4352 15818 4358 15852
rect 4392 15819 4430 15852
rect 4464 15819 4502 15853
rect 4536 15819 4542 15853
rect 4392 15818 4542 15819
rect 4352 15780 4542 15818
rect 4352 15779 4430 15780
rect 4352 15745 4358 15779
rect 4392 15746 4430 15779
rect 4464 15746 4502 15780
rect 4536 15746 4542 15780
rect 4392 15745 4542 15746
rect 4352 15707 4542 15745
rect 4352 15706 4430 15707
rect 4352 15672 4358 15706
rect 4392 15673 4430 15706
rect 4464 15673 4502 15707
rect 4536 15673 4542 15707
rect 4392 15672 4542 15673
rect 4352 15634 4542 15672
rect 4352 15633 4430 15634
rect 4352 15599 4358 15633
rect 4392 15600 4430 15633
rect 4464 15600 4502 15634
rect 4536 15600 4542 15634
rect 4392 15599 4542 15600
rect 4352 15561 4542 15599
rect 4352 15560 4430 15561
rect 4352 15526 4358 15560
rect 4392 15527 4430 15560
rect 4464 15527 4502 15561
rect 4536 15527 4542 15561
rect 4392 15526 4542 15527
rect 4352 15488 4542 15526
rect 4352 15487 4430 15488
rect 4352 15453 4358 15487
rect 4392 15454 4430 15487
rect 4464 15454 4502 15488
rect 4536 15454 4542 15488
rect 4392 15453 4542 15454
rect 4352 15415 4542 15453
rect 4352 15414 4430 15415
rect 4352 15380 4358 15414
rect 4392 15381 4430 15414
rect 4464 15381 4502 15415
rect 4536 15381 4542 15415
rect 4392 15380 4542 15381
rect 4352 15342 4542 15380
rect 4352 15341 4430 15342
rect 4352 15307 4358 15341
rect 4392 15308 4430 15341
rect 4464 15308 4502 15342
rect 4536 15308 4542 15342
rect 4392 15307 4542 15308
rect 4352 15269 4542 15307
rect 4352 15268 4430 15269
rect 4352 15234 4358 15268
rect 4392 15235 4430 15268
rect 4464 15235 4502 15269
rect 4536 15235 4542 15269
rect 4392 15234 4542 15235
rect 4352 15196 4542 15234
rect 4352 15195 4430 15196
rect 4352 15161 4358 15195
rect 4392 15162 4430 15195
rect 4464 15162 4502 15196
rect 4536 15162 4542 15196
rect 4392 15161 4542 15162
rect 4352 15123 4542 15161
rect 4352 15122 4430 15123
rect 4352 15088 4358 15122
rect 4392 15089 4430 15122
rect 4464 15089 4502 15123
rect 4536 15089 4542 15123
rect 4392 15088 4542 15089
rect 4352 15050 4542 15088
rect 4352 15049 4430 15050
rect 4352 15015 4358 15049
rect 4392 15016 4430 15049
rect 4464 15016 4502 15050
rect 4536 15016 4542 15050
rect 4392 15015 4542 15016
rect 4352 14977 4542 15015
rect 4352 14976 4430 14977
rect 4352 14942 4358 14976
rect 4392 14943 4430 14976
rect 4464 14943 4502 14977
rect 4536 14943 4542 14977
rect 4392 14942 4542 14943
rect 4352 14904 4542 14942
rect 4352 14903 4430 14904
rect 4352 14869 4358 14903
rect 4392 14870 4430 14903
rect 4464 14870 4502 14904
rect 4536 14870 4542 14904
rect 4392 14869 4542 14870
rect 4352 14831 4542 14869
rect 4352 14830 4430 14831
rect 4352 14796 4358 14830
rect 4392 14797 4430 14830
rect 4464 14797 4502 14831
rect 4536 14797 4542 14831
rect 4392 14796 4542 14797
rect 4352 14758 4542 14796
rect 4352 14757 4430 14758
rect 4352 14723 4358 14757
rect 4392 14724 4430 14757
rect 4464 14724 4502 14758
rect 4536 14724 4542 14758
rect 4392 14723 4542 14724
rect 4352 14685 4542 14723
rect 4352 14684 4430 14685
rect 4352 14650 4358 14684
rect 4392 14651 4430 14684
rect 4464 14651 4502 14685
rect 4536 14651 4542 14685
rect 4392 14650 4542 14651
rect 4352 14612 4542 14650
rect 4352 14611 4430 14612
rect 4352 14577 4358 14611
rect 4392 14578 4430 14611
rect 4464 14578 4502 14612
rect 4536 14578 4542 14612
rect 4392 14577 4542 14578
rect 4352 14539 4542 14577
rect 4352 14538 4430 14539
rect 4352 14504 4358 14538
rect 4392 14505 4430 14538
rect 4464 14505 4502 14539
rect 4536 14505 4542 14539
rect 4392 14504 4542 14505
rect 4352 14466 4542 14504
rect 4352 14465 4430 14466
rect 4352 14431 4358 14465
rect 4392 14432 4430 14465
rect 4464 14432 4502 14466
rect 4536 14432 4542 14466
rect 4392 14431 4542 14432
rect 4352 14393 4542 14431
rect 4352 14392 4430 14393
rect 4352 14358 4358 14392
rect 4392 14359 4430 14392
rect 4464 14359 4502 14393
rect 4536 14359 4542 14393
rect 4392 14358 4542 14359
rect 4352 14320 4542 14358
rect 4352 14319 4430 14320
rect 2077 14285 2234 14308
tri 2234 14285 2257 14308 nw
rect 4352 14285 4358 14319
rect 4392 14286 4430 14319
rect 4464 14286 4502 14320
rect 4536 14286 4542 14320
rect 4392 14285 4542 14286
rect 2077 14283 2232 14285
tri 2232 14283 2234 14285 nw
rect 2077 14249 2198 14283
tri 2198 14249 2232 14283 nw
tri 4347 14249 4352 14254 se
rect 4352 14249 4542 14285
rect 2077 14247 2196 14249
tri 2196 14247 2198 14249 nw
tri 4345 14247 4347 14249 se
rect 4347 14247 4542 14249
rect 2077 14246 2195 14247
tri 2195 14246 2196 14247 nw
tri 4344 14246 4345 14247 se
rect 4345 14246 4430 14247
rect 2077 14212 2161 14246
tri 2161 14212 2195 14246 nw
tri 4310 14212 4344 14246 se
rect 4344 14212 4358 14246
rect 4392 14213 4430 14246
rect 4464 14213 4502 14247
rect 4536 14213 4542 14247
rect 4392 14212 4542 14213
rect 2077 14210 2159 14212
tri 2159 14210 2161 14212 nw
tri 4308 14210 4310 14212 se
rect 4310 14210 4542 14212
rect 2077 14179 2128 14210
tri 2128 14179 2159 14210 nw
tri 4277 14179 4308 14210 se
rect 4308 14179 4542 14210
rect 2077 14176 2125 14179
tri 2125 14176 2128 14179 nw
rect 2077 14174 2123 14176
tri 2123 14174 2125 14176 nw
rect 2215 14174 4542 14179
rect 2077 14173 2122 14174
tri 2122 14173 2123 14174 nw
rect 2215 14173 4430 14174
rect 2077 14139 2088 14173
tri 2088 14139 2122 14173 nw
rect 2215 14139 2293 14173
rect 2327 14139 2367 14173
rect 2401 14139 2441 14173
rect 2475 14139 2515 14173
rect 2549 14139 2589 14173
rect 2623 14139 2663 14173
rect 2697 14139 2737 14173
rect 2771 14139 2811 14173
rect 2845 14139 2885 14173
rect 2919 14139 2959 14173
rect 2993 14139 3033 14173
rect 3067 14139 3107 14173
rect 3141 14139 3181 14173
rect 3215 14139 3255 14173
rect 3289 14139 3329 14173
rect 3363 14139 3403 14173
rect 3437 14139 3477 14173
rect 3511 14139 3551 14173
rect 3585 14139 3625 14173
rect 3659 14139 3699 14173
rect 3733 14139 3773 14173
rect 3807 14139 3847 14173
rect 3881 14139 3920 14173
rect 3954 14139 3993 14173
rect 4027 14139 4066 14173
rect 4100 14139 4139 14173
rect 4173 14139 4212 14173
rect 4246 14139 4285 14173
rect 4319 14139 4358 14173
rect 4392 14140 4430 14173
rect 4464 14140 4502 14174
rect 4536 14140 4542 14174
rect 4392 14139 4542 14140
rect 2077 14137 2086 14139
tri 2086 14137 2088 14139 nw
rect 2077 13882 2083 14137
tri 2083 14134 2086 14137 nw
rect 1821 13843 2083 13882
rect 1821 13809 1827 13843
rect 1861 13809 1899 13843
rect 1933 13809 1971 13843
rect 2005 13809 2043 13843
rect 2077 13809 2083 13843
rect 1821 13770 2083 13809
rect 1821 13736 1827 13770
rect 1861 13736 1899 13770
rect 1933 13736 1971 13770
rect 2005 13736 2043 13770
rect 2077 13736 2083 13770
rect 1821 13697 2083 13736
rect 1821 13663 1827 13697
rect 1861 13663 1899 13697
rect 1933 13663 1971 13697
rect 2005 13663 2043 13697
rect 2077 13663 2083 13697
rect 1821 13624 2083 13663
rect 1821 13590 1827 13624
rect 1861 13590 1899 13624
rect 1933 13590 1971 13624
rect 2005 13590 2043 13624
rect 2077 13590 2083 13624
rect 1821 13543 2083 13590
rect 1821 12861 1827 13543
rect 2077 13005 2083 13543
rect 2005 12966 2083 13005
rect 2005 12933 2043 12966
rect 1933 12932 2043 12933
rect 2077 12932 2083 12966
rect 1933 12894 2083 12932
rect 1933 12861 1971 12894
rect 1821 12860 1971 12861
rect 2005 12893 2083 12894
rect 2005 12860 2043 12893
rect 1821 12859 2043 12860
rect 2077 12859 2083 12893
rect 1821 12822 2083 12859
rect 1821 12788 1827 12822
rect 1861 12788 1899 12822
rect 1933 12821 2083 12822
rect 1933 12788 1971 12821
rect 1821 12787 1971 12788
rect 2005 12820 2083 12821
rect 2005 12787 2043 12820
rect 1821 12786 2043 12787
rect 2077 12786 2083 12820
rect 1821 12749 2083 12786
rect 1821 12715 1827 12749
rect 1861 12715 1899 12749
rect 1933 12748 2083 12749
rect 1933 12715 1971 12748
rect 1821 12714 1971 12715
rect 2005 12747 2083 12748
rect 2005 12714 2043 12747
rect 1821 12713 2043 12714
rect 2077 12713 2083 12747
rect 1821 12676 2083 12713
rect 1821 12642 1827 12676
rect 1861 12642 1899 12676
rect 1933 12675 2083 12676
rect 1933 12642 1971 12675
rect 1821 12641 1971 12642
rect 2005 12674 2083 12675
rect 2005 12641 2043 12674
rect 1821 12640 2043 12641
rect 2077 12640 2083 12674
rect 1821 12603 2083 12640
rect 1821 12569 1827 12603
rect 1861 12569 1899 12603
rect 1933 12602 2083 12603
rect 1933 12569 1971 12602
rect 1821 12568 1971 12569
rect 2005 12601 2083 12602
rect 2005 12568 2043 12601
rect 1821 12567 2043 12568
rect 2077 12567 2083 12601
rect 1821 12530 2083 12567
rect 1821 12496 1827 12530
rect 1861 12496 1899 12530
rect 1933 12529 2083 12530
rect 1933 12496 1971 12529
rect 1821 12495 1971 12496
rect 2005 12528 2083 12529
rect 2005 12495 2043 12528
rect 1821 12494 2043 12495
rect 2077 12494 2083 12528
rect 1821 12457 2083 12494
rect 1821 12423 1827 12457
rect 1861 12423 1899 12457
rect 1933 12456 2083 12457
rect 1933 12423 1971 12456
rect 1821 12422 1971 12423
rect 2005 12455 2083 12456
rect 2005 12422 2043 12455
rect 1821 12421 2043 12422
rect 2077 12421 2083 12455
rect 1821 12384 2083 12421
rect 1821 12350 1827 12384
rect 1861 12350 1899 12384
rect 1933 12383 2083 12384
rect 1933 12350 1971 12383
rect 1821 12349 1971 12350
rect 2005 12382 2083 12383
rect 2005 12349 2043 12382
rect 1821 12348 2043 12349
rect 2077 12348 2083 12382
rect 1821 12311 2083 12348
rect 1821 12277 1827 12311
rect 1861 12277 1899 12311
rect 1933 12310 2083 12311
rect 1933 12277 1971 12310
rect 1821 12276 1971 12277
rect 2005 12309 2083 12310
rect 2005 12276 2043 12309
rect 1821 12275 2043 12276
rect 2077 12275 2083 12309
rect 1821 12238 2083 12275
rect 1821 12204 1827 12238
rect 1861 12204 1899 12238
rect 1933 12237 2083 12238
rect 1933 12204 1971 12237
rect 1821 12203 1971 12204
rect 2005 12236 2083 12237
rect 2005 12203 2043 12236
rect 1821 12202 2043 12203
rect 2077 12202 2083 12236
rect 1821 12165 2083 12202
rect 1821 12131 1827 12165
rect 1861 12131 1899 12165
rect 1933 12164 2083 12165
rect 1933 12131 1971 12164
rect 1821 12130 1971 12131
rect 2005 12163 2083 12164
rect 2005 12130 2043 12163
rect 1821 12129 2043 12130
rect 2077 12129 2083 12163
rect 1821 12092 2083 12129
rect 1821 12058 1827 12092
rect 1861 12058 1899 12092
rect 1933 12091 2083 12092
rect 1933 12058 1971 12091
rect 1821 12057 1971 12058
rect 2005 12090 2083 12091
rect 2005 12057 2043 12090
rect 1821 12056 2043 12057
rect 2077 12056 2083 12090
rect 1821 12019 2083 12056
rect 1821 11985 1827 12019
rect 1861 11985 1899 12019
rect 1933 12018 2083 12019
rect 1933 11985 1971 12018
rect 1821 11984 1971 11985
rect 2005 12017 2083 12018
rect 2005 11984 2043 12017
rect 1821 11983 2043 11984
rect 2077 11983 2083 12017
rect 1821 11946 2083 11983
rect 1821 11912 1827 11946
rect 1861 11912 1899 11946
rect 1933 11945 2083 11946
rect 1933 11912 1971 11945
rect 1821 11911 1971 11912
rect 2005 11944 2083 11945
rect 2005 11911 2043 11944
rect 1821 11910 2043 11911
rect 2077 11910 2083 11944
rect 1821 11873 2083 11910
rect 1821 11839 1827 11873
rect 1861 11839 1899 11873
rect 1933 11872 2083 11873
rect 1933 11839 1971 11872
rect 1821 11838 1971 11839
rect 2005 11871 2083 11872
rect 2005 11838 2043 11871
rect 1821 11837 2043 11838
rect 2077 11837 2083 11871
rect 1821 11800 2083 11837
rect 1821 11766 1827 11800
rect 1861 11766 1899 11800
rect 1933 11799 2083 11800
rect 1933 11766 1971 11799
rect 1821 11765 1971 11766
rect 2005 11798 2083 11799
rect 2005 11765 2043 11798
rect 1821 11764 2043 11765
rect 2077 11764 2083 11798
rect 1821 11727 2083 11764
rect 1821 11693 1827 11727
rect 1861 11693 1899 11727
rect 1933 11726 2083 11727
rect 1933 11693 1971 11726
rect 1821 11692 1971 11693
rect 2005 11725 2083 11726
rect 2005 11692 2043 11725
rect 1821 11691 2043 11692
rect 2077 11691 2083 11725
rect 1821 11654 2083 11691
rect 1821 11620 1827 11654
rect 1861 11620 1899 11654
rect 1933 11653 2083 11654
rect 1933 11620 1971 11653
rect 1821 11619 1971 11620
rect 2005 11652 2083 11653
rect 2005 11619 2043 11652
rect 1821 11618 2043 11619
rect 2077 11618 2083 11652
rect 1821 11581 2083 11618
rect 1821 11547 1827 11581
rect 1861 11547 1899 11581
rect 1933 11580 2083 11581
rect 1933 11547 1971 11580
rect 1821 11546 1971 11547
rect 2005 11579 2083 11580
rect 2005 11546 2043 11579
rect 1821 11545 2043 11546
rect 2077 11545 2083 11579
rect 1821 11508 2083 11545
rect 1821 11474 1827 11508
rect 1861 11474 1899 11508
rect 1933 11507 2083 11508
rect 1933 11474 1971 11507
rect 1821 11473 1971 11474
rect 2005 11506 2083 11507
rect 2005 11473 2043 11506
rect 1821 11472 2043 11473
rect 2077 11472 2083 11506
rect 1821 11435 2083 11472
rect 1821 11401 1827 11435
rect 1861 11401 1899 11435
rect 1933 11434 2083 11435
rect 1933 11401 1971 11434
rect 1821 11400 1971 11401
rect 2005 11433 2083 11434
rect 2005 11400 2043 11433
rect 1821 11399 2043 11400
rect 2077 11399 2083 11433
rect 1821 11362 2083 11399
rect 1821 11328 1827 11362
rect 1861 11328 1899 11362
rect 1933 11361 2083 11362
rect 1933 11328 1971 11361
rect 1821 11327 1971 11328
rect 2005 11360 2083 11361
rect 2005 11327 2043 11360
rect 1821 11326 2043 11327
rect 2077 11326 2083 11360
rect 1821 11289 2083 11326
rect 1821 11255 1827 11289
rect 1861 11255 1899 11289
rect 1933 11288 2083 11289
rect 1933 11255 1971 11288
rect 1821 11254 1971 11255
rect 2005 11287 2083 11288
rect 2005 11254 2043 11287
rect 1821 11253 2043 11254
rect 2077 11253 2083 11287
rect 1821 11216 2083 11253
rect 1821 11182 1827 11216
rect 1861 11182 1899 11216
rect 1933 11215 2083 11216
rect 1933 11182 1971 11215
rect 1821 11181 1971 11182
rect 2005 11214 2083 11215
rect 2005 11181 2043 11214
rect 1821 11180 2043 11181
rect 2077 11180 2083 11214
rect 1821 11143 2083 11180
rect 1821 11109 1827 11143
rect 1861 11109 1899 11143
rect 1933 11142 2083 11143
rect 1933 11109 1971 11142
rect 1821 11108 1971 11109
rect 2005 11141 2083 11142
rect 2005 11108 2043 11141
rect 1821 11107 2043 11108
rect 2077 11107 2083 11141
rect 1821 11070 2083 11107
rect 1821 11036 1827 11070
rect 1861 11036 1899 11070
rect 1933 11069 2083 11070
rect 1933 11036 1971 11069
rect 1821 11035 1971 11036
rect 2005 11068 2083 11069
rect 2005 11035 2043 11068
rect 1821 11034 2043 11035
rect 2077 11034 2083 11068
rect 1821 10997 2083 11034
rect 1821 10963 1827 10997
rect 1861 10963 1899 10997
rect 1933 10996 2083 10997
rect 1933 10963 1971 10996
rect 1821 10962 1971 10963
rect 2005 10995 2083 10996
rect 2005 10962 2043 10995
rect 1821 10961 2043 10962
rect 2077 10961 2083 10995
rect 1821 10924 2083 10961
rect 1821 10890 1827 10924
rect 1861 10890 1899 10924
rect 1933 10923 2083 10924
rect 1933 10890 1971 10923
rect 1821 10889 1971 10890
rect 2005 10922 2083 10923
rect 2005 10889 2043 10922
rect 1821 10888 2043 10889
rect 2077 10888 2083 10922
rect 1821 10851 2083 10888
rect 1821 10817 1827 10851
rect 1861 10817 1899 10851
rect 1933 10850 2083 10851
rect 1933 10817 1971 10850
rect 1821 10816 1971 10817
rect 2005 10849 2083 10850
rect 2005 10816 2043 10849
rect 1821 10815 2043 10816
rect 2077 10815 2083 10849
rect 1821 10778 2083 10815
rect 1821 10744 1827 10778
rect 1861 10744 1899 10778
rect 1933 10777 2083 10778
rect 1933 10744 1971 10777
rect 1821 10743 1971 10744
rect 2005 10776 2083 10777
rect 2005 10743 2043 10776
rect 1821 10742 2043 10743
rect 2077 10742 2083 10776
rect 1821 10705 2083 10742
rect 1821 10671 1827 10705
rect 1861 10671 1899 10705
rect 1933 10704 2083 10705
rect 1933 10671 1971 10704
rect 1821 10670 1971 10671
rect 2005 10703 2083 10704
rect 2005 10670 2043 10703
rect 1821 10669 2043 10670
rect 2077 10669 2083 10703
rect 1821 10632 2083 10669
rect 1821 10598 1827 10632
rect 1861 10598 1899 10632
rect 1933 10631 2083 10632
rect 1933 10598 1971 10631
rect 1821 10597 1971 10598
rect 2005 10630 2083 10631
rect 2005 10597 2043 10630
rect 1821 10596 2043 10597
rect 2077 10596 2083 10630
rect 1821 10559 2083 10596
rect 1821 10525 1827 10559
rect 1861 10525 1899 10559
rect 1933 10558 2083 10559
rect 1933 10525 1971 10558
rect 1821 10524 1971 10525
rect 2005 10557 2083 10558
rect 2005 10524 2043 10557
rect 1821 10523 2043 10524
rect 2077 10523 2083 10557
rect 1821 10486 2083 10523
rect 1821 10452 1827 10486
rect 1861 10452 1899 10486
rect 1933 10485 2083 10486
rect 1933 10452 1971 10485
rect 1821 10451 1971 10452
rect 2005 10484 2083 10485
rect 2005 10451 2043 10484
rect 1821 10450 2043 10451
rect 2077 10450 2083 10484
rect 1821 10413 2083 10450
rect 1821 10379 1827 10413
rect 1861 10379 1899 10413
rect 1933 10412 2083 10413
rect 1933 10379 1971 10412
rect 1821 10378 1971 10379
rect 2005 10411 2083 10412
rect 2005 10378 2043 10411
rect 1821 10377 2043 10378
rect 2077 10377 2083 10411
rect 1821 10340 2083 10377
rect 1821 10306 1827 10340
rect 1861 10306 1899 10340
rect 1933 10339 2083 10340
rect 1933 10306 1971 10339
rect 1821 10305 1971 10306
rect 2005 10338 2083 10339
rect 2005 10305 2043 10338
rect 1821 10304 2043 10305
rect 2077 10304 2083 10338
rect 1821 10267 2083 10304
rect 1821 10233 1827 10267
rect 1861 10233 1899 10267
rect 1933 10266 2083 10267
rect 1933 10233 1971 10266
rect 1821 10232 1971 10233
rect 2005 10265 2083 10266
rect 2005 10232 2043 10265
rect 1821 10231 2043 10232
rect 2077 10231 2083 10265
rect 1821 10194 2083 10231
rect 1821 10160 1827 10194
rect 1861 10160 1899 10194
rect 1933 10193 2083 10194
rect 1933 10160 1971 10193
rect 1821 10159 1971 10160
rect 2005 10192 2083 10193
rect 2005 10159 2043 10192
rect 1821 10158 2043 10159
rect 2077 10158 2083 10192
rect 1821 10121 2083 10158
rect 1821 10087 1827 10121
rect 1861 10087 1899 10121
rect 1933 10120 2083 10121
rect 1933 10087 1971 10120
rect 1821 10086 1971 10087
rect 2005 10119 2083 10120
rect 2005 10086 2043 10119
rect 1821 10085 2043 10086
rect 2077 10085 2083 10119
rect 1821 10048 2083 10085
rect 1821 10014 1827 10048
rect 1861 10014 1899 10048
rect 1933 10047 2083 10048
rect 1933 10014 1971 10047
rect 1821 10013 1971 10014
rect 2005 10046 2083 10047
rect 2005 10013 2043 10046
rect 1821 10012 2043 10013
rect 2077 10012 2083 10046
rect 1821 9975 2083 10012
rect 1821 9941 1827 9975
rect 1861 9941 1899 9975
rect 1933 9974 2083 9975
rect 1933 9941 1971 9974
rect 1821 9940 1971 9941
rect 2005 9973 2083 9974
rect 2005 9940 2043 9973
rect 1821 9939 2043 9940
rect 2077 9939 2083 9973
rect 1821 9902 2083 9939
rect 1821 9868 1827 9902
rect 1861 9868 1899 9902
rect 1933 9901 2083 9902
rect 1933 9868 1971 9901
rect 1821 9867 1971 9868
rect 2005 9900 2083 9901
rect 2005 9867 2043 9900
rect 1821 9866 2043 9867
rect 2077 9866 2083 9900
rect 1821 9829 2083 9866
rect 1821 9795 1827 9829
rect 1861 9795 1899 9829
rect 1933 9828 2083 9829
rect 1933 9795 1971 9828
rect 1821 9794 1971 9795
rect 2005 9827 2083 9828
rect 2005 9794 2043 9827
rect 1821 9793 2043 9794
rect 2077 9793 2083 9827
rect 1821 9756 2083 9793
rect 1821 9722 1827 9756
rect 1861 9722 1899 9756
rect 1933 9755 2083 9756
rect 1933 9722 1971 9755
rect 1821 9721 1971 9722
rect 2005 9754 2083 9755
rect 2005 9721 2043 9754
rect 1821 9720 2043 9721
rect 2077 9720 2083 9754
rect 1821 9683 2083 9720
rect 1821 9649 1827 9683
rect 1861 9649 1899 9683
rect 1933 9682 2083 9683
rect 1933 9649 1971 9682
rect 1821 9648 1971 9649
rect 2005 9681 2083 9682
rect 2005 9648 2043 9681
rect 1821 9647 2043 9648
rect 2077 9647 2083 9681
rect 1821 9610 2083 9647
rect 1821 9576 1827 9610
rect 1861 9576 1899 9610
rect 1933 9609 2083 9610
rect 1933 9576 1971 9609
rect 1821 9575 1971 9576
rect 2005 9608 2083 9609
rect 2005 9575 2043 9608
rect 1821 9574 2043 9575
rect 2077 9574 2083 9608
rect 1821 9537 2083 9574
rect 1821 9503 1827 9537
rect 1861 9503 1899 9537
rect 1933 9536 2083 9537
rect 1933 9503 1971 9536
rect 1821 9502 1971 9503
rect 2005 9535 2083 9536
rect 2005 9502 2043 9535
rect 1821 9501 2043 9502
rect 2077 9501 2083 9535
rect 1821 9464 2083 9501
rect 1821 9430 1827 9464
rect 1861 9430 1899 9464
rect 1933 9463 2083 9464
rect 1933 9430 1971 9463
rect 1821 9429 1971 9430
rect 2005 9462 2083 9463
rect 2005 9429 2043 9462
rect 1821 9428 2043 9429
rect 2077 9428 2083 9462
rect 1821 9391 2083 9428
rect 1821 9357 1827 9391
rect 1861 9357 1899 9391
rect 1933 9390 2083 9391
rect 1933 9357 1971 9390
rect 1821 9356 1971 9357
rect 2005 9389 2083 9390
rect 2005 9356 2043 9389
rect 1821 9355 2043 9356
rect 2077 9355 2083 9389
rect 1821 9318 2083 9355
rect 1821 9284 1827 9318
rect 1861 9284 1899 9318
rect 1933 9317 2083 9318
rect 1933 9284 1971 9317
rect 1821 9283 1971 9284
rect 2005 9316 2083 9317
rect 2005 9283 2043 9316
rect 1821 9282 2043 9283
rect 2077 9282 2083 9316
rect 1821 9245 2083 9282
rect 1821 9211 1827 9245
rect 1861 9211 1899 9245
rect 1933 9244 2083 9245
rect 1933 9211 1971 9244
rect 1821 9210 1971 9211
rect 2005 9243 2083 9244
rect 2005 9210 2043 9243
rect 1821 9209 2043 9210
rect 2077 9209 2083 9243
rect 1821 9172 2083 9209
rect 1821 9138 1827 9172
rect 1861 9138 1899 9172
rect 1933 9171 2083 9172
rect 1933 9138 1971 9171
rect 1821 9137 1971 9138
rect 2005 9170 2083 9171
rect 2005 9137 2043 9170
rect 1821 9136 2043 9137
rect 2077 9136 2083 9170
rect 1821 9099 2083 9136
rect 2215 14101 4542 14139
rect 2215 14095 2293 14101
rect 2215 14061 2221 14095
rect 2255 14067 2293 14095
rect 2327 14067 2367 14101
rect 2401 14067 2441 14101
rect 2475 14067 2515 14101
rect 2549 14067 2589 14101
rect 2623 14067 2663 14101
rect 2697 14067 2737 14101
rect 2771 14067 2811 14101
rect 2845 14067 2885 14101
rect 2919 14067 2959 14101
rect 2993 14067 3033 14101
rect 3067 14067 3107 14101
rect 3141 14067 3181 14101
rect 3215 14067 3255 14101
rect 3289 14067 3329 14101
rect 3363 14067 3403 14101
rect 3437 14067 3477 14101
rect 3511 14067 3551 14101
rect 3585 14067 3625 14101
rect 3659 14067 3699 14101
rect 3733 14067 3772 14101
rect 3806 14067 3845 14101
rect 3879 14067 3918 14101
rect 3952 14067 3991 14101
rect 4025 14067 4064 14101
rect 4098 14067 4137 14101
rect 4171 14067 4210 14101
rect 4244 14067 4283 14101
rect 4317 14067 4356 14101
rect 4390 14067 4430 14101
rect 4464 14067 4502 14101
rect 4536 14067 4542 14101
rect 2255 14061 4542 14067
rect 2215 14029 4542 14061
rect 2215 14017 2365 14029
rect 2215 13983 2221 14017
rect 2255 13983 2293 14017
rect 2327 13995 2365 14017
rect 2399 13995 2439 14029
rect 2473 13995 2513 14029
rect 2547 13995 2587 14029
rect 2621 13995 2661 14029
rect 2695 13995 2735 14029
rect 2769 13995 2809 14029
rect 2843 13995 2883 14029
rect 2917 13995 2957 14029
rect 2991 13995 3031 14029
rect 3065 13995 3105 14029
rect 3139 13995 3179 14029
rect 3213 13995 3253 14029
rect 3287 13995 3327 14029
rect 3361 13995 3401 14029
rect 3435 13995 3475 14029
rect 3509 13995 3549 14029
rect 3583 13995 3623 14029
rect 3657 13995 3697 14029
rect 3731 13995 3771 14029
rect 3805 13995 3845 14029
rect 3879 13995 3918 14029
rect 3952 13995 3991 14029
rect 4025 13995 4064 14029
rect 4098 13995 4137 14029
rect 4171 13995 4210 14029
rect 4244 13995 4283 14029
rect 4317 13995 4356 14029
rect 4390 13995 4429 14029
rect 4463 13995 4542 14029
rect 2327 13989 4542 13995
rect 4605 18586 4651 18598
rect 4605 18552 4611 18586
rect 4645 18552 4651 18586
rect 4605 18513 4651 18552
rect 4605 18479 4611 18513
rect 4645 18479 4651 18513
rect 4605 18440 4651 18479
rect 4605 18406 4611 18440
rect 4645 18406 4651 18440
rect 4605 18367 4651 18406
rect 4605 18333 4611 18367
rect 4645 18333 4651 18367
rect 4605 18293 4651 18333
rect 4605 18259 4611 18293
rect 4645 18259 4651 18293
rect 4605 18219 4651 18259
rect 4605 18185 4611 18219
rect 4645 18185 4651 18219
rect 4605 18145 4651 18185
rect 4605 18111 4611 18145
rect 4645 18111 4651 18145
rect 2327 13983 2405 13989
rect 2215 13949 2405 13983
rect 2215 13939 2365 13949
rect 2215 13905 2221 13939
rect 2255 13905 2293 13939
rect 2327 13915 2365 13939
rect 2399 13915 2405 13949
rect 2327 13905 2405 13915
rect 2215 13869 2405 13905
rect 2215 13861 2365 13869
rect 2215 13827 2221 13861
rect 2255 13827 2293 13861
rect 2327 13835 2365 13861
rect 2399 13835 2405 13869
tri 2405 13859 2535 13989 nw
rect 2327 13827 2405 13835
rect 2215 13789 2405 13827
rect 2215 13783 2365 13789
rect 2215 13749 2221 13783
rect 2255 13749 2293 13783
rect 2327 13755 2365 13783
rect 2399 13755 2405 13789
rect 2327 13749 2405 13755
rect 2215 13708 2405 13749
rect 2215 13705 2365 13708
rect 2215 13671 2221 13705
rect 2255 13671 2293 13705
rect 2327 13674 2365 13705
rect 2399 13674 2405 13708
rect 2327 13671 2405 13674
rect 2215 13627 2405 13671
tri 4583 13660 4605 13682 se
rect 4605 13660 4651 18111
rect 2215 13593 2221 13627
rect 2255 13593 2293 13627
rect 2327 13593 2365 13627
rect 2399 13593 2405 13627
rect 2215 13550 2405 13593
rect 2569 13651 3514 13660
rect 2569 13642 3367 13651
rect 3419 13642 3456 13651
rect 3508 13648 3514 13651
tri 3514 13648 3526 13660 sw
tri 4571 13648 4583 13660 se
rect 4583 13648 4651 13660
rect 3508 13642 4651 13648
rect 2569 13608 3157 13642
rect 3191 13608 3230 13642
rect 3264 13608 3303 13642
rect 3337 13608 3367 13642
rect 3419 13608 3449 13642
rect 3508 13608 3522 13642
rect 3556 13608 3595 13642
rect 3629 13608 3668 13642
rect 3702 13608 3741 13642
rect 3775 13608 3813 13642
rect 3847 13608 3885 13642
rect 3919 13608 3957 13642
rect 3991 13608 4029 13642
rect 4063 13608 4101 13642
rect 4135 13608 4173 13642
rect 4207 13608 4245 13642
rect 4279 13608 4317 13642
rect 4351 13608 4389 13642
rect 4423 13608 4461 13642
rect 4495 13608 4533 13642
rect 4567 13608 4605 13642
rect 4639 13608 4651 13642
rect 2569 13599 3367 13608
rect 3419 13599 3456 13608
rect 3508 13602 4651 13608
rect 4711 17962 4901 18703
rect 4711 17890 4717 17962
rect 4895 17890 4901 17962
rect 4711 17838 4712 17890
rect 4900 17838 4901 17890
rect 4711 17826 4717 17838
rect 4895 17826 4901 17838
rect 4711 17774 4712 17826
rect 4900 17774 4901 17826
rect 4711 17762 4717 17774
rect 4895 17762 4901 17774
rect 4711 17710 4712 17762
rect 4900 17710 4901 17762
rect 4711 17698 4717 17710
rect 4895 17698 4901 17710
rect 4711 17646 4712 17698
rect 4900 17646 4901 17698
rect 4711 17634 4717 17646
rect 4895 17634 4901 17646
rect 4711 17582 4712 17634
rect 4900 17582 4901 17634
rect 4711 17570 4717 17582
rect 4895 17570 4901 17582
rect 4711 17518 4712 17570
rect 4900 17518 4901 17570
rect 4711 17506 4717 17518
rect 4895 17506 4901 17518
rect 4711 17454 4712 17506
rect 4900 17454 4901 17506
rect 4711 17442 4717 17454
rect 4895 17442 4901 17454
rect 4711 17390 4712 17442
rect 4900 17390 4901 17442
rect 4711 17378 4717 17390
rect 4895 17378 4901 17390
rect 4711 17326 4712 17378
rect 4900 17326 4901 17378
rect 4711 17314 4717 17326
rect 4895 17314 4901 17326
rect 4711 17262 4712 17314
rect 4900 17262 4901 17314
rect 4711 17250 4717 17262
rect 4895 17250 4901 17262
rect 4711 17198 4712 17250
rect 4900 17198 4901 17250
rect 4711 17186 4717 17198
rect 4895 17186 4901 17198
rect 4711 17134 4712 17186
rect 4900 17134 4901 17186
rect 4711 17122 4717 17134
rect 4895 17122 4901 17134
rect 4711 17070 4712 17122
rect 4900 17070 4901 17122
rect 4711 17058 4717 17070
rect 4895 17058 4901 17070
rect 4711 17006 4712 17058
rect 4900 17006 4901 17058
rect 4711 16994 4717 17006
rect 4895 16994 4901 17006
rect 4711 16942 4712 16994
rect 4900 16942 4901 16994
rect 4711 16929 4717 16942
rect 4895 16929 4901 16942
rect 4711 16877 4712 16929
rect 4900 16877 4901 16929
rect 4711 16864 4717 16877
rect 4895 16864 4901 16877
rect 4711 16812 4712 16864
rect 4900 16812 4901 16864
rect 4711 16799 4717 16812
rect 4895 16799 4901 16812
rect 4711 16747 4712 16799
rect 4900 16747 4901 16799
rect 4711 16734 4717 16747
rect 4895 16734 4901 16747
rect 4711 16682 4712 16734
rect 4900 16682 4901 16734
rect 4711 16669 4717 16682
rect 4895 16669 4901 16682
rect 4711 16617 4712 16669
rect 4900 16617 4901 16669
rect 4711 16604 4717 16617
rect 4895 16604 4901 16617
rect 4711 16552 4712 16604
rect 4900 16552 4901 16604
rect 4711 16539 4717 16552
rect 4895 16539 4901 16552
rect 4711 16487 4712 16539
rect 4900 16487 4901 16539
rect 4711 16474 4717 16487
rect 4895 16474 4901 16487
rect 4711 16422 4712 16474
rect 4900 16422 4901 16474
rect 4711 16409 4717 16422
rect 4895 16409 4901 16422
rect 4711 16357 4712 16409
rect 4900 16357 4901 16409
rect 4711 16344 4717 16357
rect 4895 16344 4901 16357
rect 4711 16292 4712 16344
rect 4900 16292 4901 16344
rect 4711 16279 4717 16292
rect 4895 16279 4901 16292
rect 4711 16227 4712 16279
rect 4900 16227 4901 16279
rect 4711 16214 4717 16227
rect 4895 16214 4901 16227
rect 4711 16162 4712 16214
rect 4900 16162 4901 16214
rect 4711 14760 4717 16162
rect 4895 14760 4901 16162
rect 4711 14721 4901 14760
rect 4711 14687 4717 14721
rect 4751 14687 4789 14721
rect 4823 14687 4861 14721
rect 4895 14687 4901 14721
rect 4711 14648 4901 14687
rect 4711 14614 4717 14648
rect 4751 14614 4789 14648
rect 4823 14614 4861 14648
rect 4895 14614 4901 14648
rect 4711 14575 4901 14614
rect 4711 14541 4717 14575
rect 4751 14541 4789 14575
rect 4823 14541 4861 14575
rect 4895 14541 4901 14575
rect 4711 14502 4901 14541
rect 4711 14468 4717 14502
rect 4751 14468 4789 14502
rect 4823 14468 4861 14502
rect 4895 14468 4901 14502
rect 4711 14429 4901 14468
rect 4711 14395 4717 14429
rect 4751 14395 4789 14429
rect 4823 14395 4861 14429
rect 4895 14395 4901 14429
rect 4711 14356 4901 14395
rect 4711 14322 4717 14356
rect 4751 14322 4789 14356
rect 4823 14322 4861 14356
rect 4895 14322 4901 14356
rect 4711 14283 4901 14322
rect 4711 14249 4717 14283
rect 4751 14249 4789 14283
rect 4823 14249 4861 14283
rect 4895 14249 4901 14283
rect 4711 14210 4901 14249
rect 4711 14176 4717 14210
rect 4751 14176 4789 14210
rect 4823 14176 4861 14210
rect 4895 14176 4901 14210
rect 4711 14137 4901 14176
rect 4711 14103 4717 14137
rect 4751 14103 4789 14137
rect 4823 14103 4861 14137
rect 4895 14103 4901 14137
rect 3508 13599 3514 13602
rect 2569 13593 3514 13599
rect 2569 13590 2617 13593
tri 2569 13581 2578 13590 ne
rect 2578 13581 2617 13590
tri 2578 13578 2581 13581 ne
rect 2581 13578 2617 13581
tri 2581 13559 2600 13578 ne
rect 2600 13559 2617 13578
rect 2651 13590 3514 13593
tri 3514 13590 3526 13602 nw
rect 2651 13559 2657 13590
tri 2600 13556 2603 13559 ne
rect 2603 13556 2657 13559
rect 2215 13544 2233 13550
rect 2285 13544 2335 13550
rect 2387 13544 2405 13550
tri 2603 13548 2611 13556 ne
rect 2215 11062 2221 13544
rect 2399 11134 2405 13544
rect 2327 11120 2335 11134
rect 2387 11120 2405 11134
rect 2327 11107 2405 11120
rect 2327 11062 2335 11107
rect 2387 11095 2405 11107
rect 2215 11055 2233 11062
rect 2285 11055 2335 11062
rect 2399 11061 2405 11095
rect 2387 11055 2405 11061
rect 2215 11042 2405 11055
rect 2215 11023 2233 11042
rect 2285 11023 2335 11042
rect 2215 10989 2221 11023
rect 2285 10990 2293 11023
rect 2255 10989 2293 10990
rect 2327 10990 2335 11023
rect 2387 11022 2405 11042
rect 2327 10989 2365 10990
rect 2215 10988 2365 10989
rect 2399 10988 2405 11022
rect 2215 10977 2405 10988
rect 2215 10950 2233 10977
rect 2285 10950 2335 10977
rect 2215 10916 2221 10950
rect 2285 10925 2293 10950
rect 2255 10916 2293 10925
rect 2327 10925 2335 10950
rect 2387 10949 2405 10977
rect 2327 10916 2365 10925
rect 2215 10915 2365 10916
rect 2399 10915 2405 10949
rect 2215 10912 2405 10915
rect 2215 10877 2233 10912
rect 2285 10877 2335 10912
rect 2215 10843 2221 10877
rect 2285 10860 2293 10877
rect 2255 10847 2293 10860
rect 2285 10843 2293 10847
rect 2327 10860 2335 10877
rect 2387 10876 2405 10912
rect 2327 10847 2365 10860
rect 2327 10843 2335 10847
rect 2215 10804 2233 10843
rect 2285 10804 2335 10843
rect 2399 10842 2405 10876
rect 2215 10770 2221 10804
rect 2285 10795 2293 10804
rect 2255 10782 2293 10795
rect 2285 10770 2293 10782
rect 2327 10795 2335 10804
rect 2387 10803 2405 10842
rect 2327 10782 2365 10795
rect 2327 10770 2335 10782
rect 2215 10731 2233 10770
rect 2285 10731 2335 10770
rect 2399 10769 2405 10803
rect 2215 10697 2221 10731
rect 2285 10730 2293 10731
rect 2255 10717 2293 10730
rect 2285 10697 2293 10717
rect 2327 10730 2335 10731
rect 2387 10730 2405 10769
rect 2327 10717 2365 10730
rect 2327 10697 2335 10717
rect 2215 10665 2233 10697
rect 2285 10665 2335 10697
rect 2399 10696 2405 10730
rect 2387 10665 2405 10696
rect 2215 10658 2405 10665
rect 2215 10624 2221 10658
rect 2255 10652 2293 10658
rect 2285 10624 2293 10652
rect 2327 10657 2405 10658
rect 2327 10652 2365 10657
rect 2327 10624 2335 10652
rect 2215 10600 2233 10624
rect 2285 10600 2335 10624
rect 2399 10623 2405 10657
rect 2387 10600 2405 10623
rect 2215 10587 2405 10600
rect 2215 10585 2233 10587
rect 2285 10585 2335 10587
rect 2215 10551 2221 10585
rect 2285 10551 2293 10585
rect 2327 10551 2335 10585
rect 2387 10584 2405 10587
rect 2215 10535 2233 10551
rect 2285 10535 2335 10551
rect 2399 10550 2405 10584
rect 2387 10535 2405 10550
rect 2215 10522 2405 10535
rect 2215 10512 2233 10522
rect 2285 10512 2335 10522
rect 2215 10478 2221 10512
rect 2285 10478 2293 10512
rect 2327 10478 2335 10512
rect 2387 10511 2405 10522
rect 2215 10470 2233 10478
rect 2285 10470 2335 10478
rect 2399 10477 2405 10511
rect 2387 10470 2405 10477
rect 2215 10457 2405 10470
rect 2215 10439 2233 10457
rect 2285 10439 2335 10457
rect 2215 10405 2221 10439
rect 2285 10405 2293 10439
rect 2327 10405 2335 10439
rect 2387 10438 2405 10457
rect 2215 10404 2365 10405
rect 2399 10404 2405 10438
rect 2215 10392 2405 10404
rect 2215 10366 2233 10392
rect 2285 10366 2335 10392
rect 2215 10332 2221 10366
rect 2285 10340 2293 10366
rect 2255 10332 2293 10340
rect 2327 10340 2335 10366
rect 2387 10365 2405 10392
rect 2327 10332 2365 10340
rect 2215 10331 2365 10332
rect 2399 10331 2405 10365
rect 2215 10327 2405 10331
rect 2215 10293 2233 10327
rect 2285 10293 2335 10327
rect 2215 10259 2221 10293
rect 2285 10275 2293 10293
rect 2255 10262 2293 10275
rect 2285 10259 2293 10262
rect 2327 10275 2335 10293
rect 2387 10292 2405 10327
rect 2327 10262 2365 10275
rect 2327 10259 2335 10262
rect 2215 10220 2233 10259
rect 2285 10220 2335 10259
rect 2399 10258 2405 10292
rect 2215 10186 2221 10220
rect 2285 10210 2293 10220
rect 2255 10197 2293 10210
rect 2285 10186 2293 10197
rect 2327 10210 2335 10220
rect 2387 10219 2405 10258
rect 2327 10197 2365 10210
rect 2327 10186 2335 10197
rect 2215 10147 2233 10186
rect 2285 10147 2335 10186
rect 2399 10185 2405 10219
rect 2215 10113 2221 10147
rect 2285 10145 2293 10147
rect 2255 10132 2293 10145
rect 2285 10113 2293 10132
rect 2327 10145 2335 10147
rect 2387 10146 2405 10185
rect 2327 10132 2365 10145
rect 2327 10113 2335 10132
rect 2215 10080 2233 10113
rect 2285 10080 2335 10113
rect 2399 10112 2405 10146
rect 2387 10080 2405 10112
rect 2215 10074 2405 10080
rect 2215 10040 2221 10074
rect 2255 10067 2293 10074
rect 2285 10040 2293 10067
rect 2327 10073 2405 10074
rect 2327 10067 2365 10073
rect 2327 10040 2335 10067
rect 2215 10015 2233 10040
rect 2285 10015 2335 10040
rect 2399 10039 2405 10073
rect 2387 10015 2405 10039
rect 2215 10002 2405 10015
rect 2215 10001 2233 10002
rect 2285 10001 2335 10002
rect 2215 9967 2221 10001
rect 2285 9967 2293 10001
rect 2327 9967 2335 10001
rect 2387 10000 2405 10002
rect 2215 9950 2233 9967
rect 2285 9950 2335 9967
rect 2399 9966 2405 10000
rect 2387 9950 2405 9966
rect 2215 9937 2405 9950
rect 2215 9928 2233 9937
rect 2285 9928 2335 9937
rect 2215 9894 2221 9928
rect 2285 9894 2293 9928
rect 2327 9894 2335 9928
rect 2387 9927 2405 9937
rect 2215 9885 2233 9894
rect 2285 9885 2335 9894
rect 2399 9893 2405 9927
rect 2387 9885 2405 9893
rect 2215 9872 2405 9885
rect 2215 9855 2233 9872
rect 2285 9855 2335 9872
rect 2215 9821 2221 9855
rect 2285 9821 2293 9855
rect 2327 9821 2335 9855
rect 2387 9854 2405 9872
rect 2215 9820 2233 9821
rect 2285 9820 2335 9821
rect 2399 9820 2405 9854
rect 2215 9807 2405 9820
rect 2215 9782 2233 9807
rect 2285 9782 2335 9807
rect 2215 9748 2221 9782
rect 2285 9755 2293 9782
rect 2255 9748 2293 9755
rect 2327 9755 2335 9782
rect 2387 9781 2405 9807
rect 2327 9748 2365 9755
rect 2215 9747 2365 9748
rect 2399 9747 2405 9781
rect 2215 9742 2405 9747
rect 2215 9709 2233 9742
rect 2285 9709 2335 9742
rect 2215 9675 2221 9709
rect 2285 9690 2293 9709
rect 2255 9677 2293 9690
rect 2285 9675 2293 9677
rect 2327 9690 2335 9709
rect 2387 9708 2405 9742
rect 2327 9677 2365 9690
rect 2327 9675 2335 9677
rect 2215 9636 2233 9675
rect 2285 9636 2335 9675
rect 2399 9674 2405 9708
rect 2215 9602 2221 9636
rect 2285 9625 2293 9636
rect 2255 9612 2293 9625
rect 2285 9602 2293 9612
rect 2327 9625 2335 9636
rect 2387 9635 2405 9674
rect 2327 9612 2365 9625
rect 2327 9602 2335 9612
rect 2215 9563 2233 9602
rect 2285 9563 2335 9602
rect 2399 9601 2405 9635
rect 2215 9529 2221 9563
rect 2285 9560 2293 9563
rect 2255 9547 2293 9560
rect 2285 9529 2293 9547
rect 2327 9560 2335 9563
rect 2387 9562 2405 9601
rect 2327 9547 2365 9560
rect 2327 9529 2335 9547
rect 2215 9495 2233 9529
rect 2285 9495 2335 9529
rect 2399 9528 2405 9562
rect 2387 9495 2405 9528
rect 2215 9490 2405 9495
rect 2215 9456 2221 9490
rect 2255 9482 2293 9490
rect 2285 9456 2293 9482
rect 2327 9489 2405 9490
rect 2327 9482 2365 9489
rect 2327 9456 2335 9482
rect 2215 9430 2233 9456
rect 2285 9430 2335 9456
rect 2399 9455 2405 9489
rect 2387 9430 2405 9455
rect 2215 9417 2405 9430
rect 2215 9383 2221 9417
rect 2285 9383 2293 9417
rect 2327 9383 2335 9417
rect 2387 9416 2405 9417
rect 2215 9365 2233 9383
rect 2285 9365 2335 9383
rect 2399 9382 2405 9416
rect 2387 9365 2405 9382
rect 2215 9352 2405 9365
rect 2611 13521 2657 13556
tri 2657 13548 2699 13590 nw
rect 2611 13487 2617 13521
rect 2651 13487 2657 13521
rect 2611 13449 2657 13487
rect 2611 13415 2617 13449
rect 2651 13415 2657 13449
rect 2611 13377 2657 13415
rect 2611 13343 2617 13377
rect 2651 13343 2657 13377
rect 2611 13305 2657 13343
rect 2611 13271 2617 13305
rect 2651 13271 2657 13305
rect 2611 13233 2657 13271
rect 2611 13199 2617 13233
rect 2651 13199 2657 13233
rect 2611 13161 2657 13199
rect 2611 13127 2617 13161
rect 2651 13127 2657 13161
rect 2611 13089 2657 13127
rect 2611 13055 2617 13089
rect 2651 13055 2657 13089
rect 2611 13017 2657 13055
rect 2611 12983 2617 13017
rect 2651 12983 2657 13017
rect 2611 12945 2657 12983
rect 2611 12911 2617 12945
rect 2651 12911 2657 12945
rect 2611 12873 2657 12911
rect 2611 12839 2617 12873
rect 2651 12839 2657 12873
rect 2611 12801 2657 12839
rect 2611 12767 2617 12801
rect 2651 12767 2657 12801
rect 2611 12729 2657 12767
rect 2611 12695 2617 12729
rect 2651 12695 2657 12729
rect 2611 12657 2657 12695
rect 2611 12623 2617 12657
rect 2651 12623 2657 12657
rect 2611 12585 2657 12623
rect 2611 12551 2617 12585
rect 2651 12551 2657 12585
rect 2611 12513 2657 12551
rect 2611 12479 2617 12513
rect 2651 12479 2657 12513
rect 2611 12441 2657 12479
rect 2611 12407 2617 12441
rect 2651 12407 2657 12441
rect 2611 12369 2657 12407
rect 2611 12335 2617 12369
rect 2651 12335 2657 12369
rect 2611 12297 2657 12335
rect 2611 12263 2617 12297
rect 2651 12263 2657 12297
rect 2611 12225 2657 12263
rect 2611 12191 2617 12225
rect 2651 12191 2657 12225
rect 2611 12153 2657 12191
rect 2611 12119 2617 12153
rect 2651 12119 2657 12153
rect 2611 12081 2657 12119
rect 2611 12047 2617 12081
rect 2651 12047 2657 12081
rect 2611 12009 2657 12047
rect 2611 11975 2617 12009
rect 2651 11975 2657 12009
rect 2611 11937 2657 11975
rect 2611 11903 2617 11937
rect 2651 11903 2657 11937
rect 2611 11865 2657 11903
rect 2611 11831 2617 11865
rect 2651 11831 2657 11865
rect 2611 11793 2657 11831
rect 2611 11759 2617 11793
rect 2651 11759 2657 11793
rect 2611 11721 2657 11759
rect 2611 11687 2617 11721
rect 2651 11687 2657 11721
rect 2611 11649 2657 11687
rect 2611 11615 2617 11649
rect 2651 11615 2657 11649
rect 2611 11577 2657 11615
rect 2611 11543 2617 11577
rect 2651 11543 2657 11577
rect 2611 11505 2657 11543
rect 2611 11471 2617 11505
rect 2651 11471 2657 11505
rect 2611 11433 2657 11471
rect 2611 11399 2617 11433
rect 2651 11399 2657 11433
rect 2611 11361 2657 11399
rect 2611 11327 2617 11361
rect 2651 11327 2657 11361
rect 2611 11289 2657 11327
rect 2611 11255 2617 11289
rect 2651 11255 2657 11289
rect 2611 11217 2657 11255
rect 2611 11183 2617 11217
rect 2651 11183 2657 11217
rect 2611 11145 2657 11183
rect 2611 11111 2617 11145
rect 2651 11111 2657 11145
rect 2611 11073 2657 11111
rect 2611 11039 2617 11073
rect 2651 11039 2657 11073
rect 2611 11001 2657 11039
rect 2611 10967 2617 11001
rect 2651 10967 2657 11001
rect 2611 10929 2657 10967
rect 2611 10895 2617 10929
rect 2651 10895 2657 10929
rect 2611 10857 2657 10895
rect 2611 10823 2617 10857
rect 2651 10823 2657 10857
rect 2611 10784 2657 10823
rect 2611 10750 2617 10784
rect 2651 10750 2657 10784
rect 2611 10711 2657 10750
rect 2611 10677 2617 10711
rect 2651 10677 2657 10711
rect 2611 10638 2657 10677
rect 2611 10604 2617 10638
rect 2651 10604 2657 10638
rect 2611 10565 2657 10604
rect 2611 10531 2617 10565
rect 2651 10531 2657 10565
rect 2611 10492 2657 10531
rect 2611 10458 2617 10492
rect 2651 10458 2657 10492
rect 2611 10419 2657 10458
rect 2611 10385 2617 10419
rect 2651 10385 2657 10419
rect 2611 10346 2657 10385
rect 2611 10312 2617 10346
rect 2651 10312 2657 10346
rect 2611 10273 2657 10312
rect 2611 10239 2617 10273
rect 2651 10239 2657 10273
rect 2611 10200 2657 10239
rect 2611 10166 2617 10200
rect 2651 10166 2657 10200
rect 2611 10127 2657 10166
rect 2611 10093 2617 10127
rect 2651 10093 2657 10127
rect 2611 10054 2657 10093
rect 2611 10020 2617 10054
rect 2651 10020 2657 10054
rect 2611 9981 2657 10020
rect 2611 9947 2617 9981
rect 2651 9947 2657 9981
rect 2611 9908 2657 9947
rect 2611 9874 2617 9908
rect 2651 9874 2657 9908
rect 2611 9835 2657 9874
rect 2611 9801 2617 9835
rect 2651 9801 2657 9835
rect 2611 9762 2657 9801
rect 2611 9728 2617 9762
rect 2651 9728 2657 9762
rect 2611 9689 2657 9728
rect 2611 9655 2617 9689
rect 2651 9655 2657 9689
rect 2611 9616 2657 9655
rect 2611 9582 2617 9616
rect 2651 9582 2657 9616
rect 2611 9543 2657 9582
rect 2611 9509 2617 9543
rect 2651 9509 2657 9543
rect 2611 9470 2657 9509
rect 2871 13377 3061 13383
rect 2871 13325 2872 13377
rect 2924 13371 2940 13377
rect 2992 13371 3008 13377
rect 3060 13325 3061 13377
rect 2871 13312 2877 13325
rect 3055 13312 3061 13325
rect 2871 13260 2872 13312
rect 3060 13260 3061 13312
rect 2871 13247 2877 13260
rect 3055 13247 3061 13260
rect 2871 13195 2872 13247
rect 3060 13195 3061 13247
rect 2871 13182 2877 13195
rect 3055 13182 3061 13195
rect 2871 13130 2872 13182
rect 3060 13130 3061 13182
rect 2871 13117 2877 13130
rect 3055 13117 3061 13130
rect 2871 13065 2872 13117
rect 3060 13065 3061 13117
rect 2871 13052 2877 13065
rect 3055 13052 3061 13065
rect 2871 13000 2872 13052
rect 3060 13000 3061 13052
rect 2871 12987 2877 13000
rect 3055 12987 3061 13000
rect 2871 12935 2872 12987
rect 3060 12935 3061 12987
rect 2871 12922 2877 12935
rect 3055 12922 3061 12935
rect 2871 12870 2872 12922
rect 3060 12870 3061 12922
rect 2871 12857 2877 12870
rect 3055 12857 3061 12870
rect 2871 12805 2872 12857
rect 3060 12805 3061 12857
rect 2871 12792 2877 12805
rect 3055 12792 3061 12805
rect 2871 12740 2872 12792
rect 3060 12740 3061 12792
rect 2871 12727 2877 12740
rect 3055 12727 3061 12740
rect 2871 12675 2872 12727
rect 3060 12675 3061 12727
rect 2871 12662 2877 12675
rect 3055 12662 3061 12675
rect 2871 12610 2872 12662
rect 3060 12610 3061 12662
rect 2871 12597 2877 12610
rect 3055 12597 3061 12610
rect 2871 12545 2872 12597
rect 3060 12545 3061 12597
rect 2871 12532 2877 12545
rect 3055 12532 3061 12545
rect 2871 12480 2872 12532
rect 3060 12480 3061 12532
rect 2871 12467 2877 12480
rect 3055 12467 3061 12480
rect 2871 12415 2872 12467
rect 3060 12415 3061 12467
rect 2871 12402 2877 12415
rect 3055 12402 3061 12415
rect 2871 12350 2872 12402
rect 3060 12350 3061 12402
rect 2871 12337 2877 12350
rect 3055 12337 3061 12350
rect 2871 12285 2872 12337
rect 3060 12285 3061 12337
rect 2871 12272 2877 12285
rect 3055 12272 3061 12285
rect 2871 12220 2872 12272
rect 3060 12220 3061 12272
rect 2871 12207 2877 12220
rect 3055 12207 3061 12220
rect 2871 12155 2872 12207
rect 3060 12155 3061 12207
rect 2871 12142 2877 12155
rect 3055 12142 3061 12155
rect 2871 12090 2872 12142
rect 3060 12090 3061 12142
rect 2871 12076 2877 12090
rect 3055 12076 3061 12090
rect 2871 12024 2872 12076
rect 3060 12024 3061 12076
rect 2871 12010 2877 12024
rect 3055 12010 3061 12024
rect 2871 11958 2872 12010
rect 3060 11958 3061 12010
rect 2871 11944 2877 11958
rect 3055 11944 3061 11958
rect 2871 11892 2872 11944
rect 3060 11892 3061 11944
rect 2871 11878 2877 11892
rect 3055 11878 3061 11892
rect 2871 11826 2872 11878
rect 3060 11826 3061 11878
rect 2871 11812 2877 11826
rect 3055 11812 3061 11826
rect 2871 11760 2872 11812
rect 3060 11760 3061 11812
rect 2871 11746 2877 11760
rect 3055 11746 3061 11760
rect 2871 11694 2872 11746
rect 3060 11694 3061 11746
rect 2871 11680 2877 11694
rect 3055 11680 3061 11694
rect 2871 11628 2872 11680
rect 3060 11628 3061 11680
rect 2871 11614 2877 11628
rect 3055 11614 3061 11628
rect 2871 11562 2872 11614
rect 3060 11562 3061 11614
rect 2871 10817 2877 11562
rect 3055 10817 3061 11562
rect 3791 13371 3981 13383
rect 3791 13290 3797 13371
rect 3975 13290 3981 13371
rect 3791 13238 3792 13290
rect 3980 13238 3981 13290
rect 3791 13226 3797 13238
rect 3975 13226 3981 13238
rect 3791 13174 3792 13226
rect 3980 13174 3981 13226
rect 3791 13162 3797 13174
rect 3975 13162 3981 13174
rect 3791 13110 3792 13162
rect 3980 13110 3981 13162
rect 3791 13098 3797 13110
rect 3975 13098 3981 13110
rect 3791 13046 3792 13098
rect 3980 13046 3981 13098
rect 3791 13034 3797 13046
rect 3975 13034 3981 13046
rect 3791 12982 3792 13034
rect 3980 12982 3981 13034
rect 3791 12970 3797 12982
rect 3975 12970 3981 12982
rect 3791 12918 3792 12970
rect 3980 12918 3981 12970
rect 3791 12906 3797 12918
rect 3975 12906 3981 12918
rect 3791 12854 3792 12906
rect 3980 12854 3981 12906
rect 3791 12842 3797 12854
rect 3975 12842 3981 12854
rect 3791 12790 3792 12842
rect 3980 12790 3981 12842
rect 3791 12778 3797 12790
rect 3975 12778 3981 12790
rect 3791 12726 3792 12778
rect 3980 12726 3981 12778
rect 3791 12714 3797 12726
rect 3975 12714 3981 12726
rect 3791 12662 3792 12714
rect 3980 12662 3981 12714
rect 3791 12650 3797 12662
rect 3975 12650 3981 12662
rect 3791 12598 3792 12650
rect 3980 12598 3981 12650
rect 3791 12586 3797 12598
rect 3975 12586 3981 12598
rect 3791 12534 3792 12586
rect 3980 12534 3981 12586
rect 3791 12522 3797 12534
rect 3975 12522 3981 12534
rect 3791 12470 3792 12522
rect 3980 12470 3981 12522
rect 3791 12458 3797 12470
rect 3975 12458 3981 12470
rect 3791 12406 3792 12458
rect 3980 12406 3981 12458
rect 3791 12394 3797 12406
rect 3975 12394 3981 12406
rect 3791 12342 3792 12394
rect 3980 12342 3981 12394
rect 3791 12329 3797 12342
rect 3975 12329 3981 12342
rect 3791 12277 3792 12329
rect 3980 12277 3981 12329
rect 3791 12264 3797 12277
rect 3975 12264 3981 12277
rect 3791 12212 3792 12264
rect 3980 12212 3981 12264
rect 3791 12199 3797 12212
rect 3975 12199 3981 12212
rect 3791 12147 3792 12199
rect 3980 12147 3981 12199
rect 3791 12134 3797 12147
rect 3975 12134 3981 12147
rect 3791 12082 3792 12134
rect 3980 12082 3981 12134
rect 3791 12069 3797 12082
rect 3975 12069 3981 12082
rect 3791 12017 3792 12069
rect 3980 12017 3981 12069
rect 3791 12004 3797 12017
rect 3975 12004 3981 12017
rect 3791 11952 3792 12004
rect 3980 11952 3981 12004
rect 3791 11939 3797 11952
rect 3975 11939 3981 11952
rect 3791 11887 3792 11939
rect 3980 11887 3981 11939
rect 3791 11874 3797 11887
rect 3975 11874 3981 11887
rect 3791 11822 3792 11874
rect 3980 11822 3981 11874
rect 3791 11809 3797 11822
rect 3975 11809 3981 11822
rect 3791 11757 3792 11809
rect 3980 11757 3981 11809
rect 3791 11744 3797 11757
rect 3975 11744 3981 11757
rect 3791 11692 3792 11744
rect 3980 11692 3981 11744
rect 3791 11679 3797 11692
rect 3975 11679 3981 11692
rect 3791 11627 3792 11679
rect 3980 11627 3981 11679
rect 3791 11614 3797 11627
rect 3975 11614 3981 11627
rect 3791 11562 3792 11614
rect 3980 11562 3981 11614
rect 2871 10778 3061 10817
rect 2871 10744 2877 10778
rect 2911 10744 2949 10778
rect 2983 10744 3021 10778
rect 3055 10744 3061 10778
rect 2871 10705 3061 10744
rect 2871 10671 2877 10705
rect 2911 10671 2949 10705
rect 2983 10671 3021 10705
rect 3055 10671 3061 10705
rect 2871 10632 3061 10671
rect 2871 10598 2877 10632
rect 2911 10598 2949 10632
rect 2983 10598 3021 10632
rect 3055 10598 3061 10632
rect 2871 10559 3061 10598
rect 2871 10525 2877 10559
rect 2911 10525 2949 10559
rect 2983 10525 3021 10559
rect 3055 10525 3061 10559
rect 2871 10486 3061 10525
rect 2871 10452 2877 10486
rect 2911 10452 2949 10486
rect 2983 10452 3021 10486
rect 3055 10452 3061 10486
rect 2871 10413 3061 10452
rect 2871 10379 2877 10413
rect 2911 10379 2949 10413
rect 2983 10379 3021 10413
rect 3055 10379 3061 10413
rect 2871 10340 3061 10379
rect 2871 10306 2877 10340
rect 2911 10306 2949 10340
rect 2983 10306 3021 10340
rect 3055 10306 3061 10340
rect 2871 10267 3061 10306
rect 2871 10233 2877 10267
rect 2911 10233 2949 10267
rect 2983 10233 3021 10267
rect 3055 10233 3061 10267
rect 2871 10194 3061 10233
rect 2871 10160 2877 10194
rect 2911 10160 2949 10194
rect 2983 10160 3021 10194
rect 3055 10160 3061 10194
rect 2871 10121 3061 10160
rect 2871 10087 2877 10121
rect 2911 10087 2949 10121
rect 2983 10087 3021 10121
rect 3055 10087 3061 10121
rect 2871 10048 3061 10087
rect 2871 10014 2877 10048
rect 2911 10014 2949 10048
rect 2983 10014 3021 10048
rect 3055 10014 3061 10048
rect 2871 9975 3061 10014
rect 2871 9941 2877 9975
rect 2911 9941 2949 9975
rect 2983 9941 3021 9975
rect 3055 9941 3061 9975
rect 2871 9902 3061 9941
rect 2871 9868 2877 9902
rect 2911 9868 2949 9902
rect 2983 9868 3021 9902
rect 3055 9868 3061 9902
rect 2871 9829 3061 9868
rect 2871 9795 2877 9829
rect 2911 9795 2949 9829
rect 2983 9795 3021 9829
rect 3055 9795 3061 9829
rect 2871 9756 3061 9795
rect 2871 9722 2877 9756
rect 2911 9722 2949 9756
rect 2983 9722 3021 9756
rect 3055 9722 3061 9756
rect 2871 9683 3061 9722
rect 2871 9649 2877 9683
rect 2911 9649 2949 9683
rect 2983 9649 3021 9683
rect 3055 9649 3061 9683
rect 2871 9610 3061 9649
rect 2871 9576 2877 9610
rect 2911 9576 2949 9610
rect 2983 9576 3021 9610
rect 3055 9576 3061 9610
rect 2871 9537 3061 9576
rect 2871 9503 2877 9537
rect 2911 9503 2949 9537
rect 2983 9503 3021 9537
rect 3055 9503 3061 9537
rect 2871 9491 3061 9503
rect 3361 10947 3491 10953
rect 3413 10895 3439 10947
rect 3361 10881 3491 10895
rect 3413 10829 3439 10881
rect 3361 10815 3491 10829
rect 3413 10763 3439 10815
rect 3361 10749 3491 10763
rect 3413 10697 3439 10749
rect 3361 10683 3491 10697
rect 3413 10631 3439 10683
rect 3361 10617 3491 10631
rect 3413 10565 3439 10617
rect 3361 10551 3491 10565
rect 3413 10499 3439 10551
rect 3361 10485 3491 10499
rect 3413 10433 3439 10485
rect 3361 10419 3491 10433
rect 3413 10367 3439 10419
rect 3361 10353 3491 10367
rect 3413 10301 3439 10353
rect 3361 10286 3491 10301
rect 3413 10234 3439 10286
rect 3361 10219 3491 10234
rect 3413 10167 3439 10219
rect 3361 10152 3491 10167
rect 3413 10100 3439 10152
rect 3361 10085 3491 10100
rect 3413 10033 3439 10085
rect 3361 10018 3491 10033
rect 3413 9966 3439 10018
rect 3361 9951 3491 9966
rect 3413 9899 3439 9951
rect 3361 9884 3491 9899
rect 3413 9832 3439 9884
rect 3361 9817 3491 9832
rect 3413 9765 3439 9817
rect 3361 9750 3491 9765
rect 3413 9698 3439 9750
rect 3361 9683 3491 9698
rect 3413 9631 3439 9683
rect 3361 9616 3491 9631
rect 3413 9564 3439 9616
rect 3361 9549 3491 9564
rect 3413 9497 3439 9549
rect 3361 9491 3491 9497
rect 3791 10817 3797 11562
rect 3975 10817 3981 11562
rect 4711 13362 4901 14103
rect 4711 13290 4717 13362
rect 4895 13290 4901 13362
rect 4711 13238 4712 13290
rect 4900 13238 4901 13290
rect 4711 13226 4717 13238
rect 4895 13226 4901 13238
rect 4711 13174 4712 13226
rect 4900 13174 4901 13226
rect 4711 13162 4717 13174
rect 4895 13162 4901 13174
rect 4711 13110 4712 13162
rect 4900 13110 4901 13162
rect 4711 13098 4717 13110
rect 4895 13098 4901 13110
rect 4711 13046 4712 13098
rect 4900 13046 4901 13098
rect 4711 13034 4717 13046
rect 4895 13034 4901 13046
rect 4711 12982 4712 13034
rect 4900 12982 4901 13034
rect 4711 12970 4717 12982
rect 4895 12970 4901 12982
rect 4711 12918 4712 12970
rect 4900 12918 4901 12970
rect 4711 12906 4717 12918
rect 4895 12906 4901 12918
rect 4711 12854 4712 12906
rect 4900 12854 4901 12906
rect 4711 12842 4717 12854
rect 4895 12842 4901 12854
rect 4711 12790 4712 12842
rect 4900 12790 4901 12842
rect 4711 12778 4717 12790
rect 4895 12778 4901 12790
rect 4711 12726 4712 12778
rect 4900 12726 4901 12778
rect 4711 12714 4717 12726
rect 4895 12714 4901 12726
rect 4711 12662 4712 12714
rect 4900 12662 4901 12714
rect 4711 12650 4717 12662
rect 4895 12650 4901 12662
rect 4711 12598 4712 12650
rect 4900 12598 4901 12650
rect 4711 12586 4717 12598
rect 4895 12586 4901 12598
rect 4711 12534 4712 12586
rect 4900 12534 4901 12586
rect 4711 12522 4717 12534
rect 4895 12522 4901 12534
rect 4711 12470 4712 12522
rect 4900 12470 4901 12522
rect 4711 12458 4717 12470
rect 4895 12458 4901 12470
rect 4711 12406 4712 12458
rect 4900 12406 4901 12458
rect 4711 12394 4717 12406
rect 4895 12394 4901 12406
rect 4711 12342 4712 12394
rect 4900 12342 4901 12394
rect 4711 12329 4717 12342
rect 4895 12329 4901 12342
rect 4711 12277 4712 12329
rect 4900 12277 4901 12329
rect 4711 12264 4717 12277
rect 4895 12264 4901 12277
rect 4711 12212 4712 12264
rect 4900 12212 4901 12264
rect 4711 12199 4717 12212
rect 4895 12199 4901 12212
rect 4711 12147 4712 12199
rect 4900 12147 4901 12199
rect 4711 12134 4717 12147
rect 4895 12134 4901 12147
rect 4711 12082 4712 12134
rect 4900 12082 4901 12134
rect 4711 12069 4717 12082
rect 4895 12069 4901 12082
rect 4711 12017 4712 12069
rect 4900 12017 4901 12069
rect 4711 12004 4717 12017
rect 4895 12004 4901 12017
rect 4711 11952 4712 12004
rect 4900 11952 4901 12004
rect 4711 11939 4717 11952
rect 4895 11939 4901 11952
rect 4711 11887 4712 11939
rect 4900 11887 4901 11939
rect 4711 11874 4717 11887
rect 4895 11874 4901 11887
rect 4711 11822 4712 11874
rect 4900 11822 4901 11874
rect 4711 11809 4717 11822
rect 4895 11809 4901 11822
rect 4711 11757 4712 11809
rect 4900 11757 4901 11809
rect 4711 11744 4717 11757
rect 4895 11744 4901 11757
rect 4711 11692 4712 11744
rect 4900 11692 4901 11744
rect 4711 11679 4717 11692
rect 4895 11679 4901 11692
rect 4711 11627 4712 11679
rect 4900 11627 4901 11679
rect 4711 11614 4717 11627
rect 4895 11614 4901 11627
rect 4711 11562 4712 11614
rect 4900 11562 4901 11614
rect 3791 10778 3981 10817
rect 3791 10744 3797 10778
rect 3831 10744 3869 10778
rect 3903 10744 3941 10778
rect 3975 10744 3981 10778
rect 3791 10705 3981 10744
rect 3791 10671 3797 10705
rect 3831 10671 3869 10705
rect 3903 10671 3941 10705
rect 3975 10671 3981 10705
rect 3791 10632 3981 10671
rect 3791 10598 3797 10632
rect 3831 10598 3869 10632
rect 3903 10598 3941 10632
rect 3975 10598 3981 10632
rect 3791 10559 3981 10598
rect 3791 10525 3797 10559
rect 3831 10525 3869 10559
rect 3903 10525 3941 10559
rect 3975 10525 3981 10559
rect 3791 10486 3981 10525
rect 3791 10452 3797 10486
rect 3831 10452 3869 10486
rect 3903 10452 3941 10486
rect 3975 10452 3981 10486
rect 3791 10413 3981 10452
rect 3791 10379 3797 10413
rect 3831 10379 3869 10413
rect 3903 10379 3941 10413
rect 3975 10379 3981 10413
rect 3791 10340 3981 10379
rect 3791 10306 3797 10340
rect 3831 10306 3869 10340
rect 3903 10306 3941 10340
rect 3975 10306 3981 10340
rect 3791 10267 3981 10306
rect 3791 10233 3797 10267
rect 3831 10233 3869 10267
rect 3903 10233 3941 10267
rect 3975 10233 3981 10267
rect 3791 10194 3981 10233
rect 3791 10160 3797 10194
rect 3831 10160 3869 10194
rect 3903 10160 3941 10194
rect 3975 10160 3981 10194
rect 3791 10121 3981 10160
rect 3791 10087 3797 10121
rect 3831 10087 3869 10121
rect 3903 10087 3941 10121
rect 3975 10087 3981 10121
rect 3791 10048 3981 10087
rect 3791 10014 3797 10048
rect 3831 10014 3869 10048
rect 3903 10014 3941 10048
rect 3975 10014 3981 10048
rect 3791 9975 3981 10014
rect 3791 9941 3797 9975
rect 3831 9941 3869 9975
rect 3903 9941 3941 9975
rect 3975 9941 3981 9975
rect 3791 9902 3981 9941
rect 3791 9868 3797 9902
rect 3831 9868 3869 9902
rect 3903 9868 3941 9902
rect 3975 9868 3981 9902
rect 3791 9829 3981 9868
rect 3791 9795 3797 9829
rect 3831 9795 3869 9829
rect 3903 9795 3941 9829
rect 3975 9795 3981 9829
rect 3791 9756 3981 9795
rect 3791 9722 3797 9756
rect 3831 9722 3869 9756
rect 3903 9722 3941 9756
rect 3975 9722 3981 9756
rect 3791 9683 3981 9722
rect 3791 9649 3797 9683
rect 3831 9649 3869 9683
rect 3903 9649 3941 9683
rect 3975 9649 3981 9683
rect 3791 9610 3981 9649
rect 3791 9576 3797 9610
rect 3831 9576 3869 9610
rect 3903 9576 3941 9610
rect 3975 9576 3981 9610
rect 3791 9537 3981 9576
rect 3791 9503 3797 9537
rect 3831 9503 3869 9537
rect 3903 9503 3941 9537
rect 3975 9503 3981 9537
rect 3791 9491 3981 9503
rect 4281 11225 4411 11231
rect 4333 11173 4359 11225
rect 4281 11161 4411 11173
rect 4333 11109 4359 11161
rect 4281 11097 4411 11109
rect 4333 11045 4359 11097
rect 4281 11033 4411 11045
rect 4333 10981 4359 11033
rect 4281 10969 4411 10981
rect 4333 10917 4359 10969
rect 4281 10905 4411 10917
rect 4333 10853 4359 10905
rect 4281 10841 4411 10853
rect 4333 10789 4359 10841
rect 4281 10777 4411 10789
rect 4333 10725 4359 10777
rect 4281 10713 4411 10725
rect 4333 10661 4359 10713
rect 4281 10649 4411 10661
rect 4333 10597 4359 10649
rect 4281 10585 4411 10597
rect 4333 10533 4359 10585
rect 4281 10521 4411 10533
rect 4333 10469 4359 10521
rect 4281 10457 4411 10469
rect 4333 10405 4359 10457
rect 4281 10393 4411 10405
rect 4333 10341 4359 10393
rect 4281 10329 4411 10341
rect 4333 10277 4359 10329
rect 4281 10264 4411 10277
rect 4333 10212 4359 10264
rect 4281 10199 4411 10212
rect 4333 10147 4359 10199
rect 4281 10134 4411 10147
rect 4333 10082 4359 10134
rect 4281 10069 4411 10082
rect 4333 10017 4359 10069
rect 4281 10004 4411 10017
rect 4333 9952 4359 10004
rect 4281 9939 4411 9952
rect 4333 9887 4359 9939
rect 4281 9874 4411 9887
rect 4333 9822 4359 9874
rect 4281 9809 4411 9822
rect 4333 9757 4359 9809
rect 4281 9744 4411 9757
rect 4333 9692 4359 9744
rect 4281 9679 4411 9692
rect 4333 9627 4359 9679
rect 4281 9614 4411 9627
rect 4333 9562 4359 9614
rect 4281 9549 4411 9562
rect 4333 9497 4359 9549
rect 4281 9491 4411 9497
rect 4711 10160 4717 11562
rect 4895 10160 4901 11562
rect 4711 10121 4901 10160
rect 4711 10087 4717 10121
rect 4751 10087 4789 10121
rect 4823 10087 4861 10121
rect 4895 10087 4901 10121
rect 4711 10048 4901 10087
rect 4711 10014 4717 10048
rect 4751 10014 4789 10048
rect 4823 10014 4861 10048
rect 4895 10014 4901 10048
rect 4711 9975 4901 10014
rect 4711 9941 4717 9975
rect 4751 9941 4789 9975
rect 4823 9941 4861 9975
rect 4895 9941 4901 9975
rect 4711 9902 4901 9941
rect 4711 9868 4717 9902
rect 4751 9868 4789 9902
rect 4823 9868 4861 9902
rect 4895 9868 4901 9902
rect 4711 9829 4901 9868
rect 4711 9795 4717 9829
rect 4751 9795 4789 9829
rect 4823 9795 4861 9829
rect 4895 9795 4901 9829
rect 4711 9756 4901 9795
rect 4711 9722 4717 9756
rect 4751 9722 4789 9756
rect 4823 9722 4861 9756
rect 4895 9722 4901 9756
rect 4711 9683 4901 9722
rect 4711 9649 4717 9683
rect 4751 9649 4789 9683
rect 4823 9649 4861 9683
rect 4895 9649 4901 9683
rect 4711 9610 4901 9649
rect 4711 9576 4717 9610
rect 4751 9576 4789 9610
rect 4823 9576 4861 9610
rect 4895 9576 4901 9610
rect 4711 9537 4901 9576
rect 4711 9503 4717 9537
rect 4751 9503 4789 9537
rect 4823 9503 4861 9537
rect 4895 9503 4901 9537
rect 4711 9491 4901 9503
rect 5201 20425 5331 23297
rect 5253 20373 5279 20425
rect 5201 20361 5331 20373
rect 5253 20309 5279 20361
rect 5201 20297 5331 20309
rect 5253 20245 5279 20297
rect 5201 20233 5331 20245
rect 5253 20181 5279 20233
rect 5201 20169 5331 20181
rect 5253 20117 5279 20169
rect 5201 20105 5331 20117
rect 5253 20053 5279 20105
rect 5201 20041 5331 20053
rect 5253 19989 5279 20041
rect 5201 19977 5331 19989
rect 5253 19925 5279 19977
rect 5201 19913 5331 19925
rect 5253 19861 5279 19913
rect 5201 19849 5331 19861
rect 5253 19797 5279 19849
rect 5201 19785 5331 19797
rect 5253 19733 5279 19785
rect 5201 19721 5331 19733
rect 5253 19669 5279 19721
rect 5201 19657 5331 19669
rect 5253 19605 5279 19657
rect 5201 19593 5331 19605
rect 5253 19541 5279 19593
rect 5201 19529 5331 19541
rect 5253 19477 5279 19529
rect 5201 19464 5331 19477
rect 5253 19412 5279 19464
rect 5201 19399 5331 19412
rect 5253 19347 5279 19399
rect 5201 19334 5331 19347
rect 5253 19282 5279 19334
rect 5201 19269 5331 19282
rect 5253 19217 5279 19269
rect 5201 19204 5331 19217
rect 5253 19152 5279 19204
rect 5201 19139 5331 19152
rect 5253 19087 5279 19139
rect 5201 19074 5331 19087
rect 5253 19022 5279 19074
rect 5201 19009 5331 19022
rect 5253 18957 5279 19009
rect 5201 18944 5331 18957
rect 5253 18892 5279 18944
rect 5201 18879 5331 18892
rect 5253 18827 5279 18879
rect 5201 18814 5331 18827
rect 5253 18762 5279 18814
rect 5201 18749 5331 18762
rect 5253 18697 5279 18749
rect 5201 15825 5331 18697
rect 5253 15773 5279 15825
rect 5201 15761 5331 15773
rect 5253 15709 5279 15761
rect 5201 15697 5331 15709
rect 5253 15645 5279 15697
rect 5201 15633 5331 15645
rect 5253 15581 5279 15633
rect 5201 15569 5331 15581
rect 5253 15517 5279 15569
rect 5201 15505 5331 15517
rect 5253 15453 5279 15505
rect 5201 15441 5331 15453
rect 5253 15389 5279 15441
rect 5201 15377 5331 15389
rect 5253 15325 5279 15377
rect 5201 15313 5331 15325
rect 5253 15261 5279 15313
rect 5201 15249 5331 15261
rect 5253 15197 5279 15249
rect 5201 15185 5331 15197
rect 5253 15133 5279 15185
rect 5201 15121 5331 15133
rect 5253 15069 5279 15121
rect 5201 15057 5331 15069
rect 5253 15005 5279 15057
rect 5201 14993 5331 15005
rect 5253 14941 5279 14993
rect 5201 14929 5331 14941
rect 5253 14877 5279 14929
rect 5201 14864 5331 14877
rect 5253 14812 5279 14864
rect 5201 14799 5331 14812
rect 5253 14747 5279 14799
rect 5201 14734 5331 14747
rect 5253 14682 5279 14734
rect 5201 14669 5331 14682
rect 5253 14617 5279 14669
rect 5201 14604 5331 14617
rect 5253 14552 5279 14604
rect 5201 14539 5331 14552
rect 5253 14487 5279 14539
rect 5201 14474 5331 14487
rect 5253 14422 5279 14474
rect 5201 14409 5331 14422
rect 5253 14357 5279 14409
rect 5201 14344 5331 14357
rect 5253 14292 5279 14344
rect 5201 14279 5331 14292
rect 5253 14227 5279 14279
rect 5201 14214 5331 14227
rect 5253 14162 5279 14214
rect 5201 14149 5331 14162
rect 5253 14097 5279 14149
rect 5201 11225 5331 14097
rect 5253 11173 5279 11225
rect 5201 11161 5331 11173
rect 5253 11109 5279 11161
rect 5201 11097 5331 11109
rect 5253 11045 5279 11097
rect 5201 11033 5331 11045
rect 5253 10981 5279 11033
rect 5201 10969 5331 10981
rect 5253 10917 5279 10969
rect 5201 10905 5331 10917
rect 5253 10853 5279 10905
rect 5201 10841 5331 10853
rect 5253 10789 5279 10841
rect 5201 10777 5331 10789
rect 5253 10725 5279 10777
rect 5201 10713 5331 10725
rect 5253 10661 5279 10713
rect 5201 10649 5331 10661
rect 5253 10597 5279 10649
rect 5201 10585 5331 10597
rect 5253 10533 5279 10585
rect 5201 10521 5331 10533
rect 5253 10469 5279 10521
rect 5201 10457 5331 10469
rect 5253 10405 5279 10457
rect 5201 10393 5331 10405
rect 5253 10341 5279 10393
rect 5201 10329 5331 10341
rect 5253 10277 5279 10329
rect 5201 10264 5331 10277
rect 5253 10212 5279 10264
rect 5201 10199 5331 10212
rect 5253 10147 5279 10199
rect 5201 10134 5331 10147
rect 5253 10082 5279 10134
rect 5201 10069 5331 10082
rect 5253 10017 5279 10069
rect 5201 10004 5331 10017
rect 5253 9952 5279 10004
rect 5201 9939 5331 9952
rect 5253 9887 5279 9939
rect 5201 9874 5331 9887
rect 5253 9822 5279 9874
rect 5201 9809 5331 9822
rect 5253 9757 5279 9809
rect 5201 9744 5331 9757
rect 5253 9692 5279 9744
rect 5201 9679 5331 9692
rect 5253 9627 5279 9679
rect 5201 9614 5331 9627
rect 5253 9562 5279 9614
rect 5201 9549 5331 9562
rect 5253 9497 5279 9549
rect 5201 9491 5331 9497
rect 5631 37962 5821 38003
rect 5631 37928 5637 37962
rect 5671 37928 5709 37962
rect 5743 37928 5781 37962
rect 5815 37928 5821 37962
rect 5631 37887 5821 37928
rect 5631 37853 5637 37887
rect 5671 37853 5709 37887
rect 5743 37853 5781 37887
rect 5815 37853 5821 37887
rect 5631 37812 5821 37853
rect 5631 37778 5637 37812
rect 5671 37778 5709 37812
rect 5743 37778 5781 37812
rect 5815 37778 5821 37812
rect 5631 37737 5821 37778
rect 5631 37703 5637 37737
rect 5671 37703 5709 37737
rect 5743 37703 5781 37737
rect 5815 37703 5821 37737
rect 5631 37662 5821 37703
rect 5631 37628 5637 37662
rect 5671 37628 5709 37662
rect 5743 37628 5781 37662
rect 5815 37628 5821 37662
rect 5631 37587 5821 37628
rect 5631 37553 5637 37587
rect 5671 37553 5709 37587
rect 5743 37553 5781 37587
rect 5815 37553 5821 37587
rect 5631 37512 5821 37553
rect 5631 37478 5637 37512
rect 5671 37478 5709 37512
rect 5743 37478 5781 37512
rect 5815 37478 5821 37512
rect 5631 37437 5821 37478
rect 5631 37403 5637 37437
rect 5671 37403 5709 37437
rect 5743 37403 5781 37437
rect 5815 37403 5821 37437
rect 5631 37362 5821 37403
rect 5631 37328 5637 37362
rect 5671 37328 5709 37362
rect 5743 37328 5781 37362
rect 5815 37328 5821 37362
rect 5631 37287 5821 37328
rect 5631 37253 5637 37287
rect 5671 37253 5709 37287
rect 5743 37253 5781 37287
rect 5815 37253 5821 37287
rect 5631 37212 5821 37253
rect 5631 37178 5637 37212
rect 5671 37178 5709 37212
rect 5743 37178 5781 37212
rect 5815 37178 5821 37212
rect 5631 37137 5821 37178
rect 5631 37103 5637 37137
rect 5671 37103 5709 37137
rect 5743 37103 5781 37137
rect 5815 37103 5821 37137
rect 5631 36353 5821 37103
rect 5631 36290 5637 36353
rect 5815 36290 5821 36353
rect 5631 36238 5632 36290
rect 5820 36238 5821 36290
rect 5631 36226 5637 36238
rect 5815 36226 5821 36238
rect 5631 36174 5632 36226
rect 5820 36174 5821 36226
rect 5631 36162 5637 36174
rect 5815 36162 5821 36174
rect 5631 36110 5632 36162
rect 5820 36110 5821 36162
rect 5631 36098 5637 36110
rect 5815 36098 5821 36110
rect 5631 36046 5632 36098
rect 5820 36046 5821 36098
rect 5631 36034 5637 36046
rect 5815 36034 5821 36046
rect 5631 35982 5632 36034
rect 5820 35982 5821 36034
rect 5631 35970 5637 35982
rect 5815 35970 5821 35982
rect 5631 35918 5632 35970
rect 5820 35918 5821 35970
rect 5631 35906 5637 35918
rect 5815 35906 5821 35918
rect 5631 35854 5632 35906
rect 5820 35854 5821 35906
rect 5631 35842 5637 35854
rect 5815 35842 5821 35854
rect 5631 35790 5632 35842
rect 5820 35790 5821 35842
rect 5631 35778 5637 35790
rect 5815 35778 5821 35790
rect 5631 35726 5632 35778
rect 5820 35726 5821 35778
rect 5631 35714 5637 35726
rect 5815 35714 5821 35726
rect 5631 35662 5632 35714
rect 5820 35662 5821 35714
rect 5631 35650 5637 35662
rect 5815 35650 5821 35662
rect 5631 35598 5632 35650
rect 5820 35598 5821 35650
rect 5631 35586 5637 35598
rect 5815 35586 5821 35598
rect 5631 35534 5632 35586
rect 5820 35534 5821 35586
rect 5631 35522 5637 35534
rect 5815 35522 5821 35534
rect 5631 35470 5632 35522
rect 5820 35470 5821 35522
rect 5631 35458 5637 35470
rect 5815 35458 5821 35470
rect 5631 35406 5632 35458
rect 5820 35406 5821 35458
rect 5631 35394 5637 35406
rect 5815 35394 5821 35406
rect 5631 35342 5632 35394
rect 5820 35342 5821 35394
rect 5631 35329 5637 35342
rect 5815 35329 5821 35342
rect 5631 35277 5632 35329
rect 5820 35277 5821 35329
rect 5631 35264 5637 35277
rect 5815 35264 5821 35277
rect 5631 35212 5632 35264
rect 5820 35212 5821 35264
rect 5631 35199 5637 35212
rect 5815 35199 5821 35212
rect 5631 35147 5632 35199
rect 5820 35147 5821 35199
rect 5631 35134 5637 35147
rect 5815 35134 5821 35147
rect 5631 35082 5632 35134
rect 5820 35082 5821 35134
rect 5631 35069 5637 35082
rect 5815 35069 5821 35082
rect 5631 35017 5632 35069
rect 5820 35017 5821 35069
rect 5631 35004 5637 35017
rect 5815 35004 5821 35017
rect 5631 34952 5632 35004
rect 5820 34952 5821 35004
rect 5631 34939 5637 34952
rect 5815 34939 5821 34952
rect 5631 34887 5632 34939
rect 5820 34887 5821 34939
rect 5631 34874 5637 34887
rect 5815 34874 5821 34887
rect 5631 34822 5632 34874
rect 5820 34822 5821 34874
rect 5631 34809 5637 34822
rect 5815 34809 5821 34822
rect 5631 34757 5632 34809
rect 5820 34757 5821 34809
rect 5631 34744 5637 34757
rect 5815 34744 5821 34757
rect 5631 34692 5632 34744
rect 5820 34692 5821 34744
rect 5631 34679 5637 34692
rect 5815 34679 5821 34692
rect 5631 34627 5632 34679
rect 5820 34627 5821 34679
rect 5631 34614 5637 34627
rect 5815 34614 5821 34627
rect 5631 34562 5632 34614
rect 5820 34562 5821 34614
rect 5631 32503 5637 34562
rect 5815 32503 5821 34562
rect 5631 31753 5821 32503
rect 5631 31690 5637 31753
rect 5815 31690 5821 31753
rect 5631 31638 5632 31690
rect 5820 31638 5821 31690
rect 5631 31626 5637 31638
rect 5815 31626 5821 31638
rect 5631 31574 5632 31626
rect 5820 31574 5821 31626
rect 5631 31562 5637 31574
rect 5815 31562 5821 31574
rect 5631 31510 5632 31562
rect 5820 31510 5821 31562
rect 5631 31498 5637 31510
rect 5815 31498 5821 31510
rect 5631 31446 5632 31498
rect 5820 31446 5821 31498
rect 5631 31434 5637 31446
rect 5815 31434 5821 31446
rect 5631 31382 5632 31434
rect 5820 31382 5821 31434
rect 5631 31370 5637 31382
rect 5815 31370 5821 31382
rect 5631 31318 5632 31370
rect 5820 31318 5821 31370
rect 5631 31306 5637 31318
rect 5815 31306 5821 31318
rect 5631 31254 5632 31306
rect 5820 31254 5821 31306
rect 5631 31242 5637 31254
rect 5815 31242 5821 31254
rect 5631 31190 5632 31242
rect 5820 31190 5821 31242
rect 5631 31178 5637 31190
rect 5815 31178 5821 31190
rect 5631 31126 5632 31178
rect 5820 31126 5821 31178
rect 5631 31114 5637 31126
rect 5815 31114 5821 31126
rect 5631 31062 5632 31114
rect 5820 31062 5821 31114
rect 5631 31050 5637 31062
rect 5815 31050 5821 31062
rect 5631 30998 5632 31050
rect 5820 30998 5821 31050
rect 5631 30986 5637 30998
rect 5815 30986 5821 30998
rect 5631 30934 5632 30986
rect 5820 30934 5821 30986
rect 5631 30922 5637 30934
rect 5815 30922 5821 30934
rect 5631 30870 5632 30922
rect 5820 30870 5821 30922
rect 5631 30858 5637 30870
rect 5815 30858 5821 30870
rect 5631 30806 5632 30858
rect 5820 30806 5821 30858
rect 5631 30794 5637 30806
rect 5815 30794 5821 30806
rect 5631 30742 5632 30794
rect 5820 30742 5821 30794
rect 5631 30729 5637 30742
rect 5815 30729 5821 30742
rect 5631 30677 5632 30729
rect 5820 30677 5821 30729
rect 5631 30664 5637 30677
rect 5815 30664 5821 30677
rect 5631 30612 5632 30664
rect 5820 30612 5821 30664
rect 5631 30599 5637 30612
rect 5815 30599 5821 30612
rect 5631 30547 5632 30599
rect 5820 30547 5821 30599
rect 5631 30534 5637 30547
rect 5815 30534 5821 30547
rect 5631 30482 5632 30534
rect 5820 30482 5821 30534
rect 5631 30469 5637 30482
rect 5815 30469 5821 30482
rect 5631 30417 5632 30469
rect 5820 30417 5821 30469
rect 5631 30404 5637 30417
rect 5815 30404 5821 30417
rect 5631 30352 5632 30404
rect 5820 30352 5821 30404
rect 5631 30339 5637 30352
rect 5815 30339 5821 30352
rect 5631 30287 5632 30339
rect 5820 30287 5821 30339
rect 5631 30274 5637 30287
rect 5815 30274 5821 30287
rect 5631 30222 5632 30274
rect 5820 30222 5821 30274
rect 5631 30209 5637 30222
rect 5815 30209 5821 30222
rect 5631 30157 5632 30209
rect 5820 30157 5821 30209
rect 5631 30144 5637 30157
rect 5815 30144 5821 30157
rect 5631 30092 5632 30144
rect 5820 30092 5821 30144
rect 5631 30079 5637 30092
rect 5815 30079 5821 30092
rect 5631 30027 5632 30079
rect 5820 30027 5821 30079
rect 5631 30014 5637 30027
rect 5815 30014 5821 30027
rect 5631 29962 5632 30014
rect 5820 29962 5821 30014
rect 5631 27903 5637 29962
rect 5815 27903 5821 29962
rect 5631 27162 5821 27903
rect 5631 27090 5637 27162
rect 5815 27090 5821 27162
rect 5631 27038 5632 27090
rect 5820 27038 5821 27090
rect 5631 27026 5637 27038
rect 5815 27026 5821 27038
rect 5631 26974 5632 27026
rect 5820 26974 5821 27026
rect 5631 26962 5637 26974
rect 5815 26962 5821 26974
rect 5631 26910 5632 26962
rect 5820 26910 5821 26962
rect 5631 26898 5637 26910
rect 5815 26898 5821 26910
rect 5631 26846 5632 26898
rect 5820 26846 5821 26898
rect 5631 26834 5637 26846
rect 5815 26834 5821 26846
rect 5631 26782 5632 26834
rect 5820 26782 5821 26834
rect 5631 26770 5637 26782
rect 5815 26770 5821 26782
rect 5631 26718 5632 26770
rect 5820 26718 5821 26770
rect 5631 26706 5637 26718
rect 5815 26706 5821 26718
rect 5631 26654 5632 26706
rect 5820 26654 5821 26706
rect 5631 26642 5637 26654
rect 5815 26642 5821 26654
rect 5631 26590 5632 26642
rect 5820 26590 5821 26642
rect 5631 26578 5637 26590
rect 5815 26578 5821 26590
rect 5631 26526 5632 26578
rect 5820 26526 5821 26578
rect 5631 26514 5637 26526
rect 5815 26514 5821 26526
rect 5631 26462 5632 26514
rect 5820 26462 5821 26514
rect 5631 26450 5637 26462
rect 5815 26450 5821 26462
rect 5631 26398 5632 26450
rect 5820 26398 5821 26450
rect 5631 26386 5637 26398
rect 5815 26386 5821 26398
rect 5631 26334 5632 26386
rect 5820 26334 5821 26386
rect 5631 26322 5637 26334
rect 5815 26322 5821 26334
rect 5631 26270 5632 26322
rect 5820 26270 5821 26322
rect 5631 26258 5637 26270
rect 5815 26258 5821 26270
rect 5631 26206 5632 26258
rect 5820 26206 5821 26258
rect 5631 26194 5637 26206
rect 5815 26194 5821 26206
rect 5631 26142 5632 26194
rect 5820 26142 5821 26194
rect 5631 26129 5637 26142
rect 5815 26129 5821 26142
rect 5631 26077 5632 26129
rect 5820 26077 5821 26129
rect 5631 26064 5637 26077
rect 5815 26064 5821 26077
rect 5631 26012 5632 26064
rect 5820 26012 5821 26064
rect 5631 25999 5637 26012
rect 5815 25999 5821 26012
rect 5631 25947 5632 25999
rect 5820 25947 5821 25999
rect 5631 25934 5637 25947
rect 5815 25934 5821 25947
rect 5631 25882 5632 25934
rect 5820 25882 5821 25934
rect 5631 25869 5637 25882
rect 5815 25869 5821 25882
rect 5631 25817 5632 25869
rect 5820 25817 5821 25869
rect 5631 25804 5637 25817
rect 5815 25804 5821 25817
rect 5631 25752 5632 25804
rect 5820 25752 5821 25804
rect 5631 25739 5637 25752
rect 5815 25739 5821 25752
rect 5631 25687 5632 25739
rect 5820 25687 5821 25739
rect 5631 25674 5637 25687
rect 5815 25674 5821 25687
rect 5631 25622 5632 25674
rect 5820 25622 5821 25674
rect 5631 25609 5637 25622
rect 5815 25609 5821 25622
rect 5631 25557 5632 25609
rect 5820 25557 5821 25609
rect 5631 25544 5637 25557
rect 5815 25544 5821 25557
rect 5631 25492 5632 25544
rect 5820 25492 5821 25544
rect 5631 25479 5637 25492
rect 5815 25479 5821 25492
rect 5631 25427 5632 25479
rect 5820 25427 5821 25479
rect 5631 25414 5637 25427
rect 5815 25414 5821 25427
rect 5631 25362 5632 25414
rect 5820 25362 5821 25414
rect 5631 23960 5637 25362
rect 5815 23960 5821 25362
rect 5631 23921 5821 23960
rect 5631 23887 5637 23921
rect 5671 23887 5709 23921
rect 5743 23887 5781 23921
rect 5815 23887 5821 23921
rect 5631 23848 5821 23887
rect 5631 23814 5637 23848
rect 5671 23814 5709 23848
rect 5743 23814 5781 23848
rect 5815 23814 5821 23848
rect 5631 23775 5821 23814
rect 5631 23741 5637 23775
rect 5671 23741 5709 23775
rect 5743 23741 5781 23775
rect 5815 23741 5821 23775
rect 5631 23702 5821 23741
rect 5631 23668 5637 23702
rect 5671 23668 5709 23702
rect 5743 23668 5781 23702
rect 5815 23668 5821 23702
rect 5631 23629 5821 23668
rect 5631 23595 5637 23629
rect 5671 23595 5709 23629
rect 5743 23595 5781 23629
rect 5815 23595 5821 23629
rect 5631 23556 5821 23595
rect 5631 23522 5637 23556
rect 5671 23522 5709 23556
rect 5743 23522 5781 23556
rect 5815 23522 5821 23556
rect 5631 23483 5821 23522
rect 5631 23449 5637 23483
rect 5671 23449 5709 23483
rect 5743 23449 5781 23483
rect 5815 23449 5821 23483
rect 5631 23410 5821 23449
rect 5631 23376 5637 23410
rect 5671 23376 5709 23410
rect 5743 23376 5781 23410
rect 5815 23376 5821 23410
rect 5631 23337 5821 23376
rect 5631 23303 5637 23337
rect 5671 23303 5709 23337
rect 5743 23303 5781 23337
rect 5815 23303 5821 23337
rect 5631 22571 5821 23303
rect 5631 22490 5637 22571
rect 5815 22490 5821 22571
rect 5631 22438 5632 22490
rect 5820 22438 5821 22490
rect 5631 22426 5637 22438
rect 5815 22426 5821 22438
rect 5631 22374 5632 22426
rect 5820 22374 5821 22426
rect 5631 22362 5637 22374
rect 5815 22362 5821 22374
rect 5631 22310 5632 22362
rect 5820 22310 5821 22362
rect 5631 22298 5637 22310
rect 5815 22298 5821 22310
rect 5631 22246 5632 22298
rect 5820 22246 5821 22298
rect 5631 22234 5637 22246
rect 5815 22234 5821 22246
rect 5631 22182 5632 22234
rect 5820 22182 5821 22234
rect 5631 22170 5637 22182
rect 5815 22170 5821 22182
rect 5631 22118 5632 22170
rect 5820 22118 5821 22170
rect 5631 22106 5637 22118
rect 5815 22106 5821 22118
rect 5631 22054 5632 22106
rect 5820 22054 5821 22106
rect 5631 22042 5637 22054
rect 5815 22042 5821 22054
rect 5631 21990 5632 22042
rect 5820 21990 5821 22042
rect 5631 21978 5637 21990
rect 5815 21978 5821 21990
rect 5631 21926 5632 21978
rect 5820 21926 5821 21978
rect 5631 21914 5637 21926
rect 5815 21914 5821 21926
rect 5631 21862 5632 21914
rect 5820 21862 5821 21914
rect 5631 21850 5637 21862
rect 5815 21850 5821 21862
rect 5631 21798 5632 21850
rect 5820 21798 5821 21850
rect 5631 21786 5637 21798
rect 5815 21786 5821 21798
rect 5631 21734 5632 21786
rect 5820 21734 5821 21786
rect 5631 21722 5637 21734
rect 5815 21722 5821 21734
rect 5631 21670 5632 21722
rect 5820 21670 5821 21722
rect 5631 21658 5637 21670
rect 5815 21658 5821 21670
rect 5631 21606 5632 21658
rect 5820 21606 5821 21658
rect 5631 21594 5637 21606
rect 5815 21594 5821 21606
rect 5631 21542 5632 21594
rect 5820 21542 5821 21594
rect 5631 21529 5637 21542
rect 5815 21529 5821 21542
rect 5631 21477 5632 21529
rect 5820 21477 5821 21529
rect 5631 21464 5637 21477
rect 5815 21464 5821 21477
rect 5631 21412 5632 21464
rect 5820 21412 5821 21464
rect 5631 21399 5637 21412
rect 5815 21399 5821 21412
rect 5631 21347 5632 21399
rect 5820 21347 5821 21399
rect 5631 21334 5637 21347
rect 5815 21334 5821 21347
rect 5631 21282 5632 21334
rect 5820 21282 5821 21334
rect 5631 21269 5637 21282
rect 5815 21269 5821 21282
rect 5631 21217 5632 21269
rect 5820 21217 5821 21269
rect 5631 21204 5637 21217
rect 5815 21204 5821 21217
rect 5631 21152 5632 21204
rect 5820 21152 5821 21204
rect 5631 21139 5637 21152
rect 5815 21139 5821 21152
rect 5631 21087 5632 21139
rect 5820 21087 5821 21139
rect 5631 21074 5637 21087
rect 5815 21074 5821 21087
rect 5631 21022 5632 21074
rect 5820 21022 5821 21074
rect 5631 21009 5637 21022
rect 5815 21009 5821 21022
rect 5631 20957 5632 21009
rect 5820 20957 5821 21009
rect 5631 20944 5637 20957
rect 5815 20944 5821 20957
rect 5631 20892 5632 20944
rect 5820 20892 5821 20944
rect 5631 20879 5637 20892
rect 5815 20879 5821 20892
rect 5631 20827 5632 20879
rect 5820 20827 5821 20879
rect 5631 20814 5637 20827
rect 5815 20814 5821 20827
rect 5631 20762 5632 20814
rect 5820 20762 5821 20814
rect 5631 20017 5637 20762
rect 5815 20017 5821 20762
rect 5631 19978 5821 20017
rect 5631 19944 5637 19978
rect 5671 19944 5709 19978
rect 5743 19944 5781 19978
rect 5815 19944 5821 19978
rect 5631 19905 5821 19944
rect 5631 19871 5637 19905
rect 5671 19871 5709 19905
rect 5743 19871 5781 19905
rect 5815 19871 5821 19905
rect 5631 19832 5821 19871
rect 5631 19798 5637 19832
rect 5671 19798 5709 19832
rect 5743 19798 5781 19832
rect 5815 19798 5821 19832
rect 5631 19759 5821 19798
rect 5631 19725 5637 19759
rect 5671 19725 5709 19759
rect 5743 19725 5781 19759
rect 5815 19725 5821 19759
rect 5631 19686 5821 19725
rect 5631 19652 5637 19686
rect 5671 19652 5709 19686
rect 5743 19652 5781 19686
rect 5815 19652 5821 19686
rect 5631 19613 5821 19652
rect 5631 19579 5637 19613
rect 5671 19579 5709 19613
rect 5743 19579 5781 19613
rect 5815 19579 5821 19613
rect 5631 19540 5821 19579
rect 5631 19506 5637 19540
rect 5671 19506 5709 19540
rect 5743 19506 5781 19540
rect 5815 19506 5821 19540
rect 5631 19467 5821 19506
rect 5631 19433 5637 19467
rect 5671 19433 5709 19467
rect 5743 19433 5781 19467
rect 5815 19433 5821 19467
rect 5631 19394 5821 19433
rect 5631 19360 5637 19394
rect 5671 19360 5709 19394
rect 5743 19360 5781 19394
rect 5815 19360 5821 19394
rect 5631 19321 5821 19360
rect 5631 19287 5637 19321
rect 5671 19287 5709 19321
rect 5743 19287 5781 19321
rect 5815 19287 5821 19321
rect 5631 19248 5821 19287
rect 5631 19214 5637 19248
rect 5671 19214 5709 19248
rect 5743 19214 5781 19248
rect 5815 19214 5821 19248
rect 5631 19175 5821 19214
rect 5631 19141 5637 19175
rect 5671 19141 5709 19175
rect 5743 19141 5781 19175
rect 5815 19141 5821 19175
rect 5631 19102 5821 19141
rect 5631 19068 5637 19102
rect 5671 19068 5709 19102
rect 5743 19068 5781 19102
rect 5815 19068 5821 19102
rect 5631 19029 5821 19068
rect 5631 18995 5637 19029
rect 5671 18995 5709 19029
rect 5743 18995 5781 19029
rect 5815 18995 5821 19029
rect 5631 18956 5821 18995
rect 5631 18922 5637 18956
rect 5671 18922 5709 18956
rect 5743 18922 5781 18956
rect 5815 18922 5821 18956
rect 5631 18883 5821 18922
rect 5631 18849 5637 18883
rect 5671 18849 5709 18883
rect 5743 18849 5781 18883
rect 5815 18849 5821 18883
rect 5631 18810 5821 18849
rect 5631 18776 5637 18810
rect 5671 18776 5709 18810
rect 5743 18776 5781 18810
rect 5815 18776 5821 18810
rect 5631 18737 5821 18776
rect 5631 18703 5637 18737
rect 5671 18703 5709 18737
rect 5743 18703 5781 18737
rect 5815 18703 5821 18737
rect 5631 17962 5821 18703
rect 5631 17890 5637 17962
rect 5815 17890 5821 17962
rect 5631 17838 5632 17890
rect 5820 17838 5821 17890
rect 5631 17826 5637 17838
rect 5815 17826 5821 17838
rect 5631 17774 5632 17826
rect 5820 17774 5821 17826
rect 5631 17762 5637 17774
rect 5815 17762 5821 17774
rect 5631 17710 5632 17762
rect 5820 17710 5821 17762
rect 5631 17698 5637 17710
rect 5815 17698 5821 17710
rect 5631 17646 5632 17698
rect 5820 17646 5821 17698
rect 5631 17634 5637 17646
rect 5815 17634 5821 17646
rect 5631 17582 5632 17634
rect 5820 17582 5821 17634
rect 5631 17570 5637 17582
rect 5815 17570 5821 17582
rect 5631 17518 5632 17570
rect 5820 17518 5821 17570
rect 5631 17506 5637 17518
rect 5815 17506 5821 17518
rect 5631 17454 5632 17506
rect 5820 17454 5821 17506
rect 5631 17442 5637 17454
rect 5815 17442 5821 17454
rect 5631 17390 5632 17442
rect 5820 17390 5821 17442
rect 5631 17378 5637 17390
rect 5815 17378 5821 17390
rect 5631 17326 5632 17378
rect 5820 17326 5821 17378
rect 5631 17314 5637 17326
rect 5815 17314 5821 17326
rect 5631 17262 5632 17314
rect 5820 17262 5821 17314
rect 5631 17250 5637 17262
rect 5815 17250 5821 17262
rect 5631 17198 5632 17250
rect 5820 17198 5821 17250
rect 5631 17186 5637 17198
rect 5815 17186 5821 17198
rect 5631 17134 5632 17186
rect 5820 17134 5821 17186
rect 5631 17122 5637 17134
rect 5815 17122 5821 17134
rect 5631 17070 5632 17122
rect 5820 17070 5821 17122
rect 5631 17058 5637 17070
rect 5815 17058 5821 17070
rect 5631 17006 5632 17058
rect 5820 17006 5821 17058
rect 5631 16994 5637 17006
rect 5815 16994 5821 17006
rect 5631 16942 5632 16994
rect 5820 16942 5821 16994
rect 5631 16929 5637 16942
rect 5815 16929 5821 16942
rect 5631 16877 5632 16929
rect 5820 16877 5821 16929
rect 5631 16864 5637 16877
rect 5815 16864 5821 16877
rect 5631 16812 5632 16864
rect 5820 16812 5821 16864
rect 5631 16799 5637 16812
rect 5815 16799 5821 16812
rect 5631 16747 5632 16799
rect 5820 16747 5821 16799
rect 5631 16734 5637 16747
rect 5815 16734 5821 16747
rect 5631 16682 5632 16734
rect 5820 16682 5821 16734
rect 5631 16669 5637 16682
rect 5815 16669 5821 16682
rect 5631 16617 5632 16669
rect 5820 16617 5821 16669
rect 5631 16604 5637 16617
rect 5815 16604 5821 16617
rect 5631 16552 5632 16604
rect 5820 16552 5821 16604
rect 5631 16539 5637 16552
rect 5815 16539 5821 16552
rect 5631 16487 5632 16539
rect 5820 16487 5821 16539
rect 5631 16474 5637 16487
rect 5815 16474 5821 16487
rect 5631 16422 5632 16474
rect 5820 16422 5821 16474
rect 5631 16409 5637 16422
rect 5815 16409 5821 16422
rect 5631 16357 5632 16409
rect 5820 16357 5821 16409
rect 5631 16344 5637 16357
rect 5815 16344 5821 16357
rect 5631 16292 5632 16344
rect 5820 16292 5821 16344
rect 5631 16279 5637 16292
rect 5815 16279 5821 16292
rect 5631 16227 5632 16279
rect 5820 16227 5821 16279
rect 5631 16214 5637 16227
rect 5815 16214 5821 16227
rect 5631 16162 5632 16214
rect 5820 16162 5821 16214
rect 5631 14760 5637 16162
rect 5815 14760 5821 16162
rect 5631 14721 5821 14760
rect 5631 14687 5637 14721
rect 5671 14687 5709 14721
rect 5743 14687 5781 14721
rect 5815 14687 5821 14721
rect 5631 14648 5821 14687
rect 5631 14614 5637 14648
rect 5671 14614 5709 14648
rect 5743 14614 5781 14648
rect 5815 14614 5821 14648
rect 5631 14575 5821 14614
rect 5631 14541 5637 14575
rect 5671 14541 5709 14575
rect 5743 14541 5781 14575
rect 5815 14541 5821 14575
rect 5631 14502 5821 14541
rect 5631 14468 5637 14502
rect 5671 14468 5709 14502
rect 5743 14468 5781 14502
rect 5815 14468 5821 14502
rect 5631 14429 5821 14468
rect 5631 14395 5637 14429
rect 5671 14395 5709 14429
rect 5743 14395 5781 14429
rect 5815 14395 5821 14429
rect 5631 14356 5821 14395
rect 5631 14322 5637 14356
rect 5671 14322 5709 14356
rect 5743 14322 5781 14356
rect 5815 14322 5821 14356
rect 5631 14283 5821 14322
rect 5631 14249 5637 14283
rect 5671 14249 5709 14283
rect 5743 14249 5781 14283
rect 5815 14249 5821 14283
rect 5631 14210 5821 14249
rect 5631 14176 5637 14210
rect 5671 14176 5709 14210
rect 5743 14176 5781 14210
rect 5815 14176 5821 14210
rect 5631 14137 5821 14176
rect 5631 14103 5637 14137
rect 5671 14103 5709 14137
rect 5743 14103 5781 14137
rect 5815 14103 5821 14137
rect 5631 13362 5821 14103
rect 5631 13290 5637 13362
rect 5815 13290 5821 13362
rect 5631 13238 5632 13290
rect 5820 13238 5821 13290
rect 5631 13226 5637 13238
rect 5815 13226 5821 13238
rect 5631 13174 5632 13226
rect 5820 13174 5821 13226
rect 5631 13162 5637 13174
rect 5815 13162 5821 13174
rect 5631 13110 5632 13162
rect 5820 13110 5821 13162
rect 5631 13098 5637 13110
rect 5815 13098 5821 13110
rect 5631 13046 5632 13098
rect 5820 13046 5821 13098
rect 5631 13034 5637 13046
rect 5815 13034 5821 13046
rect 5631 12982 5632 13034
rect 5820 12982 5821 13034
rect 5631 12970 5637 12982
rect 5815 12970 5821 12982
rect 5631 12918 5632 12970
rect 5820 12918 5821 12970
rect 5631 12906 5637 12918
rect 5815 12906 5821 12918
rect 5631 12854 5632 12906
rect 5820 12854 5821 12906
rect 5631 12842 5637 12854
rect 5815 12842 5821 12854
rect 5631 12790 5632 12842
rect 5820 12790 5821 12842
rect 5631 12778 5637 12790
rect 5815 12778 5821 12790
rect 5631 12726 5632 12778
rect 5820 12726 5821 12778
rect 5631 12714 5637 12726
rect 5815 12714 5821 12726
rect 5631 12662 5632 12714
rect 5820 12662 5821 12714
rect 5631 12650 5637 12662
rect 5815 12650 5821 12662
rect 5631 12598 5632 12650
rect 5820 12598 5821 12650
rect 5631 12586 5637 12598
rect 5815 12586 5821 12598
rect 5631 12534 5632 12586
rect 5820 12534 5821 12586
rect 5631 12522 5637 12534
rect 5815 12522 5821 12534
rect 5631 12470 5632 12522
rect 5820 12470 5821 12522
rect 5631 12458 5637 12470
rect 5815 12458 5821 12470
rect 5631 12406 5632 12458
rect 5820 12406 5821 12458
rect 5631 12394 5637 12406
rect 5815 12394 5821 12406
rect 5631 12342 5632 12394
rect 5820 12342 5821 12394
rect 5631 12329 5637 12342
rect 5815 12329 5821 12342
rect 5631 12277 5632 12329
rect 5820 12277 5821 12329
rect 5631 12264 5637 12277
rect 5815 12264 5821 12277
rect 5631 12212 5632 12264
rect 5820 12212 5821 12264
rect 5631 12199 5637 12212
rect 5815 12199 5821 12212
rect 5631 12147 5632 12199
rect 5820 12147 5821 12199
rect 5631 12134 5637 12147
rect 5815 12134 5821 12147
rect 5631 12082 5632 12134
rect 5820 12082 5821 12134
rect 5631 12069 5637 12082
rect 5815 12069 5821 12082
rect 5631 12017 5632 12069
rect 5820 12017 5821 12069
rect 5631 12004 5637 12017
rect 5815 12004 5821 12017
rect 5631 11952 5632 12004
rect 5820 11952 5821 12004
rect 5631 11939 5637 11952
rect 5815 11939 5821 11952
rect 5631 11887 5632 11939
rect 5820 11887 5821 11939
rect 5631 11874 5637 11887
rect 5815 11874 5821 11887
rect 5631 11822 5632 11874
rect 5820 11822 5821 11874
rect 5631 11809 5637 11822
rect 5815 11809 5821 11822
rect 5631 11757 5632 11809
rect 5820 11757 5821 11809
rect 5631 11744 5637 11757
rect 5815 11744 5821 11757
rect 5631 11692 5632 11744
rect 5820 11692 5821 11744
rect 5631 11679 5637 11692
rect 5815 11679 5821 11692
rect 5631 11627 5632 11679
rect 5820 11627 5821 11679
rect 5631 11614 5637 11627
rect 5815 11614 5821 11627
rect 5631 11562 5632 11614
rect 5820 11562 5821 11614
rect 5631 10160 5637 11562
rect 5815 10160 5821 11562
rect 5631 10121 5821 10160
rect 5631 10087 5637 10121
rect 5671 10087 5709 10121
rect 5743 10087 5781 10121
rect 5815 10087 5821 10121
rect 5631 10048 5821 10087
rect 5631 10014 5637 10048
rect 5671 10014 5709 10048
rect 5743 10014 5781 10048
rect 5815 10014 5821 10048
rect 5631 9975 5821 10014
rect 5631 9941 5637 9975
rect 5671 9941 5709 9975
rect 5743 9941 5781 9975
rect 5815 9941 5821 9975
rect 5631 9902 5821 9941
rect 5631 9868 5637 9902
rect 5671 9868 5709 9902
rect 5743 9868 5781 9902
rect 5815 9868 5821 9902
rect 5631 9829 5821 9868
rect 5631 9795 5637 9829
rect 5671 9795 5709 9829
rect 5743 9795 5781 9829
rect 5815 9795 5821 9829
rect 5631 9756 5821 9795
rect 5631 9722 5637 9756
rect 5671 9722 5709 9756
rect 5743 9722 5781 9756
rect 5815 9722 5821 9756
rect 5631 9683 5821 9722
rect 5631 9649 5637 9683
rect 5671 9649 5709 9683
rect 5743 9649 5781 9683
rect 5815 9649 5821 9683
rect 5631 9610 5821 9649
rect 5631 9576 5637 9610
rect 5671 9576 5709 9610
rect 5743 9576 5781 9610
rect 5815 9576 5821 9610
rect 5631 9537 5821 9576
rect 5631 9503 5637 9537
rect 5671 9503 5709 9537
rect 5743 9503 5781 9537
rect 5815 9503 5821 9537
rect 5631 9491 5821 9503
rect 6121 37997 6251 38003
rect 6173 37945 6199 37997
rect 6121 37929 6251 37945
rect 6173 37877 6199 37929
rect 6121 37861 6251 37877
rect 6173 37809 6199 37861
rect 6121 37793 6251 37809
rect 6173 37741 6199 37793
rect 6121 37725 6251 37741
rect 6173 37673 6199 37725
rect 6121 37657 6251 37673
rect 6173 37605 6199 37657
rect 6121 37589 6251 37605
rect 6173 37537 6199 37589
rect 6121 37521 6251 37537
rect 6173 37469 6199 37521
rect 6121 37453 6251 37469
rect 6173 37401 6199 37453
rect 6121 37385 6251 37401
rect 6173 37333 6199 37385
rect 6121 37318 6251 37333
rect 6173 37266 6199 37318
rect 6121 37251 6251 37266
rect 6173 37199 6199 37251
rect 6121 37184 6251 37199
rect 6173 37132 6199 37184
rect 6121 37117 6251 37132
rect 6173 37065 6199 37117
rect 6121 34225 6251 37065
rect 6173 34173 6199 34225
rect 6121 34161 6251 34173
rect 6173 34109 6199 34161
rect 6121 34097 6251 34109
rect 6173 34045 6199 34097
rect 6121 34033 6251 34045
rect 6173 33981 6199 34033
rect 6121 33969 6251 33981
rect 6173 33917 6199 33969
rect 6121 33905 6251 33917
rect 6173 33853 6199 33905
rect 6121 33841 6251 33853
rect 6173 33789 6199 33841
rect 6121 33777 6251 33789
rect 6173 33725 6199 33777
rect 6121 33713 6251 33725
rect 6173 33661 6199 33713
rect 6121 33649 6251 33661
rect 6173 33597 6199 33649
rect 6121 33585 6251 33597
rect 6173 33533 6199 33585
rect 6121 33521 6251 33533
rect 6173 33469 6199 33521
rect 6121 33457 6251 33469
rect 6173 33405 6199 33457
rect 6121 33393 6251 33405
rect 6173 33341 6199 33393
rect 6121 33329 6251 33341
rect 6173 33277 6199 33329
rect 6121 33264 6251 33277
rect 6173 33212 6199 33264
rect 6121 33199 6251 33212
rect 6173 33147 6199 33199
rect 6121 33134 6251 33147
rect 6173 33082 6199 33134
rect 6121 33069 6251 33082
rect 6173 33017 6199 33069
rect 6121 33004 6251 33017
rect 6173 32952 6199 33004
rect 6121 32939 6251 32952
rect 6173 32887 6199 32939
rect 6121 32874 6251 32887
rect 6173 32822 6199 32874
rect 6121 32809 6251 32822
rect 6173 32757 6199 32809
rect 6121 32744 6251 32757
rect 6173 32692 6199 32744
rect 6121 32679 6251 32692
rect 6173 32627 6199 32679
rect 6121 32614 6251 32627
rect 6173 32562 6199 32614
rect 6121 32549 6251 32562
rect 6173 32497 6199 32549
rect 6121 29625 6251 32497
rect 6173 29573 6199 29625
rect 6121 29561 6251 29573
rect 6173 29509 6199 29561
rect 6121 29497 6251 29509
rect 6173 29445 6199 29497
rect 6121 29433 6251 29445
rect 6173 29381 6199 29433
rect 6121 29369 6251 29381
rect 6173 29317 6199 29369
rect 6121 29305 6251 29317
rect 6173 29253 6199 29305
rect 6121 29241 6251 29253
rect 6173 29189 6199 29241
rect 6121 29177 6251 29189
rect 6173 29125 6199 29177
rect 6121 29113 6251 29125
rect 6173 29061 6199 29113
rect 6121 29049 6251 29061
rect 6173 28997 6199 29049
rect 6121 28985 6251 28997
rect 6173 28933 6199 28985
rect 6121 28921 6251 28933
rect 6173 28869 6199 28921
rect 6121 28857 6251 28869
rect 6173 28805 6199 28857
rect 6121 28793 6251 28805
rect 6173 28741 6199 28793
rect 6121 28729 6251 28741
rect 6173 28677 6199 28729
rect 6121 28664 6251 28677
rect 6173 28612 6199 28664
rect 6121 28599 6251 28612
rect 6173 28547 6199 28599
rect 6121 28534 6251 28547
rect 6173 28482 6199 28534
rect 6121 28469 6251 28482
rect 6173 28417 6199 28469
rect 6121 28404 6251 28417
rect 6173 28352 6199 28404
rect 6121 28339 6251 28352
rect 6173 28287 6199 28339
rect 6121 28274 6251 28287
rect 6173 28222 6199 28274
rect 6121 28209 6251 28222
rect 6173 28157 6199 28209
rect 6121 28144 6251 28157
rect 6173 28092 6199 28144
rect 6121 28079 6251 28092
rect 6173 28027 6199 28079
rect 6121 28014 6251 28027
rect 6173 27962 6199 28014
rect 6121 27949 6251 27962
rect 6173 27897 6199 27949
rect 6121 25025 6251 27897
rect 6173 24973 6199 25025
rect 6121 24961 6251 24973
rect 6173 24909 6199 24961
rect 6121 24897 6251 24909
rect 6173 24845 6199 24897
rect 6121 24833 6251 24845
rect 6173 24781 6199 24833
rect 6121 24769 6251 24781
rect 6173 24717 6199 24769
rect 6121 24705 6251 24717
rect 6173 24653 6199 24705
rect 6121 24641 6251 24653
rect 6173 24589 6199 24641
rect 6121 24577 6251 24589
rect 6173 24525 6199 24577
rect 6121 24513 6251 24525
rect 6173 24461 6199 24513
rect 6121 24449 6251 24461
rect 6173 24397 6199 24449
rect 6121 24385 6251 24397
rect 6173 24333 6199 24385
rect 6121 24321 6251 24333
rect 6173 24269 6199 24321
rect 6121 24257 6251 24269
rect 6173 24205 6199 24257
rect 6121 24193 6251 24205
rect 6173 24141 6199 24193
rect 6121 24129 6251 24141
rect 6173 24077 6199 24129
rect 6121 24064 6251 24077
rect 6173 24012 6199 24064
rect 6121 23999 6251 24012
rect 6173 23947 6199 23999
rect 6121 23934 6251 23947
rect 6173 23882 6199 23934
rect 6121 23869 6251 23882
rect 6173 23817 6199 23869
rect 6121 23804 6251 23817
rect 6173 23752 6199 23804
rect 6121 23739 6251 23752
rect 6173 23687 6199 23739
rect 6121 23674 6251 23687
rect 6173 23622 6199 23674
rect 6121 23609 6251 23622
rect 6173 23557 6199 23609
rect 6121 23544 6251 23557
rect 6173 23492 6199 23544
rect 6121 23479 6251 23492
rect 6173 23427 6199 23479
rect 6121 23414 6251 23427
rect 6173 23362 6199 23414
rect 6121 23349 6251 23362
rect 6173 23297 6199 23349
rect 6121 20425 6251 23297
rect 6173 20373 6199 20425
rect 6121 20361 6251 20373
rect 6173 20309 6199 20361
rect 6121 20297 6251 20309
rect 6173 20245 6199 20297
rect 6121 20233 6251 20245
rect 6173 20181 6199 20233
rect 6121 20169 6251 20181
rect 6173 20117 6199 20169
rect 6121 20105 6251 20117
rect 6173 20053 6199 20105
rect 6121 20041 6251 20053
rect 6173 19989 6199 20041
rect 6121 19977 6251 19989
rect 6173 19925 6199 19977
rect 6121 19913 6251 19925
rect 6173 19861 6199 19913
rect 6121 19849 6251 19861
rect 6173 19797 6199 19849
rect 6121 19785 6251 19797
rect 6173 19733 6199 19785
rect 6121 19721 6251 19733
rect 6173 19669 6199 19721
rect 6121 19657 6251 19669
rect 6173 19605 6199 19657
rect 6121 19593 6251 19605
rect 6173 19541 6199 19593
rect 6121 19529 6251 19541
rect 6173 19477 6199 19529
rect 6121 19464 6251 19477
rect 6173 19412 6199 19464
rect 6121 19399 6251 19412
rect 6173 19347 6199 19399
rect 6121 19334 6251 19347
rect 6173 19282 6199 19334
rect 6121 19269 6251 19282
rect 6173 19217 6199 19269
rect 6121 19204 6251 19217
rect 6173 19152 6199 19204
rect 6121 19139 6251 19152
rect 6173 19087 6199 19139
rect 6121 19074 6251 19087
rect 6173 19022 6199 19074
rect 6121 19009 6251 19022
rect 6173 18957 6199 19009
rect 6121 18944 6251 18957
rect 6173 18892 6199 18944
rect 6121 18879 6251 18892
rect 6173 18827 6199 18879
rect 6121 18814 6251 18827
rect 6173 18762 6199 18814
rect 6121 18749 6251 18762
rect 6173 18697 6199 18749
rect 6121 15825 6251 18697
rect 6173 15773 6199 15825
rect 6121 15761 6251 15773
rect 6173 15709 6199 15761
rect 6121 15697 6251 15709
rect 6173 15645 6199 15697
rect 6121 15633 6251 15645
rect 6173 15581 6199 15633
rect 6121 15569 6251 15581
rect 6173 15517 6199 15569
rect 6121 15505 6251 15517
rect 6173 15453 6199 15505
rect 6121 15441 6251 15453
rect 6173 15389 6199 15441
rect 6121 15377 6251 15389
rect 6173 15325 6199 15377
rect 6121 15313 6251 15325
rect 6173 15261 6199 15313
rect 6121 15249 6251 15261
rect 6173 15197 6199 15249
rect 6121 15185 6251 15197
rect 6173 15133 6199 15185
rect 6121 15121 6251 15133
rect 6173 15069 6199 15121
rect 6121 15057 6251 15069
rect 6173 15005 6199 15057
rect 6121 14993 6251 15005
rect 6173 14941 6199 14993
rect 6121 14929 6251 14941
rect 6173 14877 6199 14929
rect 6121 14864 6251 14877
rect 6173 14812 6199 14864
rect 6121 14799 6251 14812
rect 6173 14747 6199 14799
rect 6121 14734 6251 14747
rect 6173 14682 6199 14734
rect 6121 14669 6251 14682
rect 6173 14617 6199 14669
rect 6121 14604 6251 14617
rect 6173 14552 6199 14604
rect 6121 14539 6251 14552
rect 6173 14487 6199 14539
rect 6121 14474 6251 14487
rect 6173 14422 6199 14474
rect 6121 14409 6251 14422
rect 6173 14357 6199 14409
rect 6121 14344 6251 14357
rect 6173 14292 6199 14344
rect 6121 14279 6251 14292
rect 6173 14227 6199 14279
rect 6121 14214 6251 14227
rect 6173 14162 6199 14214
rect 6121 14149 6251 14162
rect 6173 14097 6199 14149
rect 6121 11225 6251 14097
rect 6173 11173 6199 11225
rect 6121 11161 6251 11173
rect 6173 11109 6199 11161
rect 6121 11097 6251 11109
rect 6173 11045 6199 11097
rect 6121 11033 6251 11045
rect 6173 10981 6199 11033
rect 6121 10969 6251 10981
rect 6173 10917 6199 10969
rect 6121 10905 6251 10917
rect 6173 10853 6199 10905
rect 6121 10841 6251 10853
rect 6173 10789 6199 10841
rect 6121 10777 6251 10789
rect 6173 10725 6199 10777
rect 6121 10713 6251 10725
rect 6173 10661 6199 10713
rect 6121 10649 6251 10661
rect 6173 10597 6199 10649
rect 6121 10585 6251 10597
rect 6173 10533 6199 10585
rect 6121 10521 6251 10533
rect 6173 10469 6199 10521
rect 6121 10457 6251 10469
rect 6173 10405 6199 10457
rect 6121 10393 6251 10405
rect 6173 10341 6199 10393
rect 6121 10329 6251 10341
rect 6173 10277 6199 10329
rect 6121 10264 6251 10277
rect 6173 10212 6199 10264
rect 6121 10199 6251 10212
rect 6173 10147 6199 10199
rect 6121 10134 6251 10147
rect 6173 10082 6199 10134
rect 6121 10069 6251 10082
rect 6173 10017 6199 10069
rect 6121 10004 6251 10017
rect 6173 9952 6199 10004
rect 6121 9939 6251 9952
rect 6173 9887 6199 9939
rect 6121 9874 6251 9887
rect 6173 9822 6199 9874
rect 6121 9809 6251 9822
rect 6173 9757 6199 9809
rect 6121 9744 6251 9757
rect 6173 9692 6199 9744
rect 6121 9679 6251 9692
rect 6173 9627 6199 9679
rect 6121 9614 6251 9627
rect 6173 9562 6199 9614
rect 6121 9549 6251 9562
rect 6173 9497 6199 9549
rect 6121 9491 6251 9497
rect 6551 37962 6741 38003
rect 6551 37928 6557 37962
rect 6591 37928 6629 37962
rect 6663 37928 6701 37962
rect 6735 37928 6741 37962
rect 6551 37887 6741 37928
rect 6551 37853 6557 37887
rect 6591 37853 6629 37887
rect 6663 37853 6701 37887
rect 6735 37853 6741 37887
rect 6551 37812 6741 37853
rect 6551 37778 6557 37812
rect 6591 37778 6629 37812
rect 6663 37778 6701 37812
rect 6735 37778 6741 37812
rect 6551 37737 6741 37778
rect 6551 37703 6557 37737
rect 6591 37703 6629 37737
rect 6663 37703 6701 37737
rect 6735 37703 6741 37737
rect 6551 37662 6741 37703
rect 6551 37628 6557 37662
rect 6591 37628 6629 37662
rect 6663 37628 6701 37662
rect 6735 37628 6741 37662
rect 6551 37587 6741 37628
rect 6551 37553 6557 37587
rect 6591 37553 6629 37587
rect 6663 37553 6701 37587
rect 6735 37553 6741 37587
rect 6551 37512 6741 37553
rect 6551 37478 6557 37512
rect 6591 37478 6629 37512
rect 6663 37478 6701 37512
rect 6735 37478 6741 37512
rect 6551 37437 6741 37478
rect 6551 37403 6557 37437
rect 6591 37403 6629 37437
rect 6663 37403 6701 37437
rect 6735 37403 6741 37437
rect 6551 37362 6741 37403
rect 6551 37328 6557 37362
rect 6591 37328 6629 37362
rect 6663 37328 6701 37362
rect 6735 37328 6741 37362
rect 6551 37287 6741 37328
rect 6551 37253 6557 37287
rect 6591 37253 6629 37287
rect 6663 37253 6701 37287
rect 6735 37253 6741 37287
rect 6551 37212 6741 37253
rect 6551 37178 6557 37212
rect 6591 37178 6629 37212
rect 6663 37178 6701 37212
rect 6735 37178 6741 37212
rect 6551 37137 6741 37178
rect 6551 37103 6557 37137
rect 6591 37103 6629 37137
rect 6663 37103 6701 37137
rect 6735 37103 6741 37137
rect 6551 36353 6741 37103
rect 6551 36290 6557 36353
rect 6735 36290 6741 36353
rect 6551 36238 6552 36290
rect 6740 36238 6741 36290
rect 6551 36226 6557 36238
rect 6735 36226 6741 36238
rect 6551 36174 6552 36226
rect 6740 36174 6741 36226
rect 6551 36162 6557 36174
rect 6735 36162 6741 36174
rect 6551 36110 6552 36162
rect 6740 36110 6741 36162
rect 6551 36098 6557 36110
rect 6735 36098 6741 36110
rect 6551 36046 6552 36098
rect 6740 36046 6741 36098
rect 6551 36034 6557 36046
rect 6735 36034 6741 36046
rect 6551 35982 6552 36034
rect 6740 35982 6741 36034
rect 6551 35970 6557 35982
rect 6735 35970 6741 35982
rect 6551 35918 6552 35970
rect 6740 35918 6741 35970
rect 6551 35906 6557 35918
rect 6735 35906 6741 35918
rect 6551 35854 6552 35906
rect 6740 35854 6741 35906
rect 6551 35842 6557 35854
rect 6735 35842 6741 35854
rect 6551 35790 6552 35842
rect 6740 35790 6741 35842
rect 6551 35778 6557 35790
rect 6735 35778 6741 35790
rect 6551 35726 6552 35778
rect 6740 35726 6741 35778
rect 6551 35714 6557 35726
rect 6735 35714 6741 35726
rect 6551 35662 6552 35714
rect 6740 35662 6741 35714
rect 6551 35650 6557 35662
rect 6735 35650 6741 35662
rect 6551 35598 6552 35650
rect 6740 35598 6741 35650
rect 6551 35586 6557 35598
rect 6735 35586 6741 35598
rect 6551 35534 6552 35586
rect 6740 35534 6741 35586
rect 6551 35522 6557 35534
rect 6735 35522 6741 35534
rect 6551 35470 6552 35522
rect 6740 35470 6741 35522
rect 6551 35458 6557 35470
rect 6735 35458 6741 35470
rect 6551 35406 6552 35458
rect 6740 35406 6741 35458
rect 6551 35394 6557 35406
rect 6735 35394 6741 35406
rect 6551 35342 6552 35394
rect 6740 35342 6741 35394
rect 6551 35329 6557 35342
rect 6735 35329 6741 35342
rect 6551 35277 6552 35329
rect 6740 35277 6741 35329
rect 6551 35264 6557 35277
rect 6735 35264 6741 35277
rect 6551 35212 6552 35264
rect 6740 35212 6741 35264
rect 6551 35199 6557 35212
rect 6735 35199 6741 35212
rect 6551 35147 6552 35199
rect 6740 35147 6741 35199
rect 6551 35134 6557 35147
rect 6735 35134 6741 35147
rect 6551 35082 6552 35134
rect 6740 35082 6741 35134
rect 6551 35069 6557 35082
rect 6735 35069 6741 35082
rect 6551 35017 6552 35069
rect 6740 35017 6741 35069
rect 6551 35004 6557 35017
rect 6735 35004 6741 35017
rect 6551 34952 6552 35004
rect 6740 34952 6741 35004
rect 6551 34939 6557 34952
rect 6735 34939 6741 34952
rect 6551 34887 6552 34939
rect 6740 34887 6741 34939
rect 6551 34874 6557 34887
rect 6735 34874 6741 34887
rect 6551 34822 6552 34874
rect 6740 34822 6741 34874
rect 6551 34809 6557 34822
rect 6735 34809 6741 34822
rect 6551 34757 6552 34809
rect 6740 34757 6741 34809
rect 6551 34744 6557 34757
rect 6735 34744 6741 34757
rect 6551 34692 6552 34744
rect 6740 34692 6741 34744
rect 6551 34679 6557 34692
rect 6735 34679 6741 34692
rect 6551 34627 6552 34679
rect 6740 34627 6741 34679
rect 6551 34614 6557 34627
rect 6735 34614 6741 34627
rect 6551 34562 6552 34614
rect 6740 34562 6741 34614
rect 6551 32503 6557 34562
rect 6735 32503 6741 34562
rect 6551 31753 6741 32503
rect 6551 31690 6557 31753
rect 6735 31690 6741 31753
rect 6551 31638 6552 31690
rect 6740 31638 6741 31690
rect 6551 31626 6557 31638
rect 6735 31626 6741 31638
rect 6551 31574 6552 31626
rect 6740 31574 6741 31626
rect 6551 31562 6557 31574
rect 6735 31562 6741 31574
rect 6551 31510 6552 31562
rect 6740 31510 6741 31562
rect 6551 31498 6557 31510
rect 6735 31498 6741 31510
rect 6551 31446 6552 31498
rect 6740 31446 6741 31498
rect 6551 31434 6557 31446
rect 6735 31434 6741 31446
rect 6551 31382 6552 31434
rect 6740 31382 6741 31434
rect 6551 31370 6557 31382
rect 6735 31370 6741 31382
rect 6551 31318 6552 31370
rect 6740 31318 6741 31370
rect 6551 31306 6557 31318
rect 6735 31306 6741 31318
rect 6551 31254 6552 31306
rect 6740 31254 6741 31306
rect 6551 31242 6557 31254
rect 6735 31242 6741 31254
rect 6551 31190 6552 31242
rect 6740 31190 6741 31242
rect 6551 31178 6557 31190
rect 6735 31178 6741 31190
rect 6551 31126 6552 31178
rect 6740 31126 6741 31178
rect 6551 31114 6557 31126
rect 6735 31114 6741 31126
rect 6551 31062 6552 31114
rect 6740 31062 6741 31114
rect 6551 31050 6557 31062
rect 6735 31050 6741 31062
rect 6551 30998 6552 31050
rect 6740 30998 6741 31050
rect 6551 30986 6557 30998
rect 6735 30986 6741 30998
rect 6551 30934 6552 30986
rect 6740 30934 6741 30986
rect 6551 30922 6557 30934
rect 6735 30922 6741 30934
rect 6551 30870 6552 30922
rect 6740 30870 6741 30922
rect 6551 30858 6557 30870
rect 6735 30858 6741 30870
rect 6551 30806 6552 30858
rect 6740 30806 6741 30858
rect 6551 30794 6557 30806
rect 6735 30794 6741 30806
rect 6551 30742 6552 30794
rect 6740 30742 6741 30794
rect 6551 30729 6557 30742
rect 6735 30729 6741 30742
rect 6551 30677 6552 30729
rect 6740 30677 6741 30729
rect 6551 30664 6557 30677
rect 6735 30664 6741 30677
rect 6551 30612 6552 30664
rect 6740 30612 6741 30664
rect 6551 30599 6557 30612
rect 6735 30599 6741 30612
rect 6551 30547 6552 30599
rect 6740 30547 6741 30599
rect 6551 30534 6557 30547
rect 6735 30534 6741 30547
rect 6551 30482 6552 30534
rect 6740 30482 6741 30534
rect 6551 30469 6557 30482
rect 6735 30469 6741 30482
rect 6551 30417 6552 30469
rect 6740 30417 6741 30469
rect 6551 30404 6557 30417
rect 6735 30404 6741 30417
rect 6551 30352 6552 30404
rect 6740 30352 6741 30404
rect 6551 30339 6557 30352
rect 6735 30339 6741 30352
rect 6551 30287 6552 30339
rect 6740 30287 6741 30339
rect 6551 30274 6557 30287
rect 6735 30274 6741 30287
rect 6551 30222 6552 30274
rect 6740 30222 6741 30274
rect 6551 30209 6557 30222
rect 6735 30209 6741 30222
rect 6551 30157 6552 30209
rect 6740 30157 6741 30209
rect 6551 30144 6557 30157
rect 6735 30144 6741 30157
rect 6551 30092 6552 30144
rect 6740 30092 6741 30144
rect 6551 30079 6557 30092
rect 6735 30079 6741 30092
rect 6551 30027 6552 30079
rect 6740 30027 6741 30079
rect 6551 30014 6557 30027
rect 6735 30014 6741 30027
rect 6551 29962 6552 30014
rect 6740 29962 6741 30014
rect 6551 27903 6557 29962
rect 6735 27903 6741 29962
rect 6551 27153 6741 27903
rect 6551 27090 6557 27153
rect 6735 27090 6741 27153
rect 6551 27038 6552 27090
rect 6740 27038 6741 27090
rect 6551 27026 6557 27038
rect 6735 27026 6741 27038
rect 6551 26974 6552 27026
rect 6740 26974 6741 27026
rect 6551 26962 6557 26974
rect 6735 26962 6741 26974
rect 6551 26910 6552 26962
rect 6740 26910 6741 26962
rect 6551 26898 6557 26910
rect 6735 26898 6741 26910
rect 6551 26846 6552 26898
rect 6740 26846 6741 26898
rect 6551 26834 6557 26846
rect 6735 26834 6741 26846
rect 6551 26782 6552 26834
rect 6740 26782 6741 26834
rect 6551 26770 6557 26782
rect 6735 26770 6741 26782
rect 6551 26718 6552 26770
rect 6740 26718 6741 26770
rect 6551 26706 6557 26718
rect 6735 26706 6741 26718
rect 6551 26654 6552 26706
rect 6740 26654 6741 26706
rect 6551 26642 6557 26654
rect 6735 26642 6741 26654
rect 6551 26590 6552 26642
rect 6740 26590 6741 26642
rect 6551 26578 6557 26590
rect 6735 26578 6741 26590
rect 6551 26526 6552 26578
rect 6740 26526 6741 26578
rect 6551 26514 6557 26526
rect 6735 26514 6741 26526
rect 6551 26462 6552 26514
rect 6740 26462 6741 26514
rect 6551 26450 6557 26462
rect 6735 26450 6741 26462
rect 6551 26398 6552 26450
rect 6740 26398 6741 26450
rect 6551 26386 6557 26398
rect 6735 26386 6741 26398
rect 6551 26334 6552 26386
rect 6740 26334 6741 26386
rect 6551 26322 6557 26334
rect 6735 26322 6741 26334
rect 6551 26270 6552 26322
rect 6740 26270 6741 26322
rect 6551 26258 6557 26270
rect 6735 26258 6741 26270
rect 6551 26206 6552 26258
rect 6740 26206 6741 26258
rect 6551 26194 6557 26206
rect 6735 26194 6741 26206
rect 6551 26142 6552 26194
rect 6740 26142 6741 26194
rect 6551 26129 6557 26142
rect 6735 26129 6741 26142
rect 6551 26077 6552 26129
rect 6740 26077 6741 26129
rect 6551 26064 6557 26077
rect 6735 26064 6741 26077
rect 6551 26012 6552 26064
rect 6740 26012 6741 26064
rect 6551 25999 6557 26012
rect 6735 25999 6741 26012
rect 6551 25947 6552 25999
rect 6740 25947 6741 25999
rect 6551 25934 6557 25947
rect 6735 25934 6741 25947
rect 6551 25882 6552 25934
rect 6740 25882 6741 25934
rect 6551 25869 6557 25882
rect 6735 25869 6741 25882
rect 6551 25817 6552 25869
rect 6740 25817 6741 25869
rect 6551 25804 6557 25817
rect 6735 25804 6741 25817
rect 6551 25752 6552 25804
rect 6740 25752 6741 25804
rect 6551 25739 6557 25752
rect 6735 25739 6741 25752
rect 6551 25687 6552 25739
rect 6740 25687 6741 25739
rect 6551 25674 6557 25687
rect 6735 25674 6741 25687
rect 6551 25622 6552 25674
rect 6740 25622 6741 25674
rect 6551 25609 6557 25622
rect 6735 25609 6741 25622
rect 6551 25557 6552 25609
rect 6740 25557 6741 25609
rect 6551 25544 6557 25557
rect 6735 25544 6741 25557
rect 6551 25492 6552 25544
rect 6740 25492 6741 25544
rect 6551 25479 6557 25492
rect 6735 25479 6741 25492
rect 6551 25427 6552 25479
rect 6740 25427 6741 25479
rect 6551 25414 6557 25427
rect 6735 25414 6741 25427
rect 6551 25362 6552 25414
rect 6740 25362 6741 25414
rect 6551 23303 6557 25362
rect 6735 23303 6741 25362
rect 6551 22562 6741 23303
rect 6551 22490 6557 22562
rect 6735 22490 6741 22562
rect 6551 22438 6552 22490
rect 6740 22438 6741 22490
rect 6551 22426 6557 22438
rect 6735 22426 6741 22438
rect 6551 22374 6552 22426
rect 6740 22374 6741 22426
rect 6551 22362 6557 22374
rect 6735 22362 6741 22374
rect 6551 22310 6552 22362
rect 6740 22310 6741 22362
rect 6551 22298 6557 22310
rect 6735 22298 6741 22310
rect 6551 22246 6552 22298
rect 6740 22246 6741 22298
rect 6551 22234 6557 22246
rect 6735 22234 6741 22246
rect 6551 22182 6552 22234
rect 6740 22182 6741 22234
rect 6551 22170 6557 22182
rect 6735 22170 6741 22182
rect 6551 22118 6552 22170
rect 6740 22118 6741 22170
rect 6551 22106 6557 22118
rect 6735 22106 6741 22118
rect 6551 22054 6552 22106
rect 6740 22054 6741 22106
rect 6551 22042 6557 22054
rect 6735 22042 6741 22054
rect 6551 21990 6552 22042
rect 6740 21990 6741 22042
rect 6551 21978 6557 21990
rect 6735 21978 6741 21990
rect 6551 21926 6552 21978
rect 6740 21926 6741 21978
rect 6551 21914 6557 21926
rect 6735 21914 6741 21926
rect 6551 21862 6552 21914
rect 6740 21862 6741 21914
rect 6551 21850 6557 21862
rect 6735 21850 6741 21862
rect 6551 21798 6552 21850
rect 6740 21798 6741 21850
rect 6551 21786 6557 21798
rect 6735 21786 6741 21798
rect 6551 21734 6552 21786
rect 6740 21734 6741 21786
rect 6551 21722 6557 21734
rect 6735 21722 6741 21734
rect 6551 21670 6552 21722
rect 6740 21670 6741 21722
rect 6551 21658 6557 21670
rect 6735 21658 6741 21670
rect 6551 21606 6552 21658
rect 6740 21606 6741 21658
rect 6551 21594 6557 21606
rect 6735 21594 6741 21606
rect 6551 21542 6552 21594
rect 6740 21542 6741 21594
rect 6551 21529 6557 21542
rect 6735 21529 6741 21542
rect 6551 21477 6552 21529
rect 6740 21477 6741 21529
rect 6551 21464 6557 21477
rect 6735 21464 6741 21477
rect 6551 21412 6552 21464
rect 6740 21412 6741 21464
rect 6551 21399 6557 21412
rect 6735 21399 6741 21412
rect 6551 21347 6552 21399
rect 6740 21347 6741 21399
rect 6551 21334 6557 21347
rect 6735 21334 6741 21347
rect 6551 21282 6552 21334
rect 6740 21282 6741 21334
rect 6551 21269 6557 21282
rect 6735 21269 6741 21282
rect 6551 21217 6552 21269
rect 6740 21217 6741 21269
rect 6551 21204 6557 21217
rect 6735 21204 6741 21217
rect 6551 21152 6552 21204
rect 6740 21152 6741 21204
rect 6551 21139 6557 21152
rect 6735 21139 6741 21152
rect 6551 21087 6552 21139
rect 6740 21087 6741 21139
rect 6551 21074 6557 21087
rect 6735 21074 6741 21087
rect 6551 21022 6552 21074
rect 6740 21022 6741 21074
rect 6551 21009 6557 21022
rect 6735 21009 6741 21022
rect 6551 20957 6552 21009
rect 6740 20957 6741 21009
rect 6551 20944 6557 20957
rect 6735 20944 6741 20957
rect 6551 20892 6552 20944
rect 6740 20892 6741 20944
rect 6551 20879 6557 20892
rect 6735 20879 6741 20892
rect 6551 20827 6552 20879
rect 6740 20827 6741 20879
rect 6551 20814 6557 20827
rect 6735 20814 6741 20827
rect 6551 20762 6552 20814
rect 6740 20762 6741 20814
rect 6551 19360 6557 20762
rect 6735 19360 6741 20762
rect 6551 19321 6741 19360
rect 6551 19287 6557 19321
rect 6591 19287 6629 19321
rect 6663 19287 6701 19321
rect 6735 19287 6741 19321
rect 6551 19248 6741 19287
rect 6551 19214 6557 19248
rect 6591 19214 6629 19248
rect 6663 19214 6701 19248
rect 6735 19214 6741 19248
rect 6551 19175 6741 19214
rect 6551 19141 6557 19175
rect 6591 19141 6629 19175
rect 6663 19141 6701 19175
rect 6735 19141 6741 19175
rect 6551 19102 6741 19141
rect 6551 19068 6557 19102
rect 6591 19068 6629 19102
rect 6663 19068 6701 19102
rect 6735 19068 6741 19102
rect 6551 19029 6741 19068
rect 6551 18995 6557 19029
rect 6591 18995 6629 19029
rect 6663 18995 6701 19029
rect 6735 18995 6741 19029
rect 6551 18956 6741 18995
rect 6551 18922 6557 18956
rect 6591 18922 6629 18956
rect 6663 18922 6701 18956
rect 6735 18922 6741 18956
rect 6551 18883 6741 18922
rect 6551 18849 6557 18883
rect 6591 18849 6629 18883
rect 6663 18849 6701 18883
rect 6735 18849 6741 18883
rect 6551 18810 6741 18849
rect 6551 18776 6557 18810
rect 6591 18776 6629 18810
rect 6663 18776 6701 18810
rect 6735 18776 6741 18810
rect 6551 18737 6741 18776
rect 6551 18703 6557 18737
rect 6591 18703 6629 18737
rect 6663 18703 6701 18737
rect 6735 18703 6741 18737
rect 6551 17953 6741 18703
rect 6551 17890 6557 17953
rect 6735 17890 6741 17953
rect 6551 17838 6552 17890
rect 6740 17838 6741 17890
rect 6551 17826 6557 17838
rect 6735 17826 6741 17838
rect 6551 17774 6552 17826
rect 6740 17774 6741 17826
rect 6551 17762 6557 17774
rect 6735 17762 6741 17774
rect 6551 17710 6552 17762
rect 6740 17710 6741 17762
rect 6551 17698 6557 17710
rect 6735 17698 6741 17710
rect 6551 17646 6552 17698
rect 6740 17646 6741 17698
rect 6551 17634 6557 17646
rect 6735 17634 6741 17646
rect 6551 17582 6552 17634
rect 6740 17582 6741 17634
rect 6551 17570 6557 17582
rect 6735 17570 6741 17582
rect 6551 17518 6552 17570
rect 6740 17518 6741 17570
rect 6551 17506 6557 17518
rect 6735 17506 6741 17518
rect 6551 17454 6552 17506
rect 6740 17454 6741 17506
rect 6551 17442 6557 17454
rect 6735 17442 6741 17454
rect 6551 17390 6552 17442
rect 6740 17390 6741 17442
rect 6551 17378 6557 17390
rect 6735 17378 6741 17390
rect 6551 17326 6552 17378
rect 6740 17326 6741 17378
rect 6551 17314 6557 17326
rect 6735 17314 6741 17326
rect 6551 17262 6552 17314
rect 6740 17262 6741 17314
rect 6551 17250 6557 17262
rect 6735 17250 6741 17262
rect 6551 17198 6552 17250
rect 6740 17198 6741 17250
rect 6551 17186 6557 17198
rect 6735 17186 6741 17198
rect 6551 17134 6552 17186
rect 6740 17134 6741 17186
rect 6551 17122 6557 17134
rect 6735 17122 6741 17134
rect 6551 17070 6552 17122
rect 6740 17070 6741 17122
rect 6551 17058 6557 17070
rect 6735 17058 6741 17070
rect 6551 17006 6552 17058
rect 6740 17006 6741 17058
rect 6551 16994 6557 17006
rect 6735 16994 6741 17006
rect 6551 16942 6552 16994
rect 6740 16942 6741 16994
rect 6551 16929 6557 16942
rect 6735 16929 6741 16942
rect 6551 16877 6552 16929
rect 6740 16877 6741 16929
rect 6551 16864 6557 16877
rect 6735 16864 6741 16877
rect 6551 16812 6552 16864
rect 6740 16812 6741 16864
rect 6551 16799 6557 16812
rect 6735 16799 6741 16812
rect 6551 16747 6552 16799
rect 6740 16747 6741 16799
rect 6551 16734 6557 16747
rect 6735 16734 6741 16747
rect 6551 16682 6552 16734
rect 6740 16682 6741 16734
rect 6551 16669 6557 16682
rect 6735 16669 6741 16682
rect 6551 16617 6552 16669
rect 6740 16617 6741 16669
rect 6551 16604 6557 16617
rect 6735 16604 6741 16617
rect 6551 16552 6552 16604
rect 6740 16552 6741 16604
rect 6551 16539 6557 16552
rect 6735 16539 6741 16552
rect 6551 16487 6552 16539
rect 6740 16487 6741 16539
rect 6551 16474 6557 16487
rect 6735 16474 6741 16487
rect 6551 16422 6552 16474
rect 6740 16422 6741 16474
rect 6551 16409 6557 16422
rect 6735 16409 6741 16422
rect 6551 16357 6552 16409
rect 6740 16357 6741 16409
rect 6551 16344 6557 16357
rect 6735 16344 6741 16357
rect 6551 16292 6552 16344
rect 6740 16292 6741 16344
rect 6551 16279 6557 16292
rect 6735 16279 6741 16292
rect 6551 16227 6552 16279
rect 6740 16227 6741 16279
rect 6551 16214 6557 16227
rect 6735 16214 6741 16227
rect 6551 16162 6552 16214
rect 6740 16162 6741 16214
rect 6551 14103 6557 16162
rect 6735 14103 6741 16162
rect 6551 13362 6741 14103
rect 6551 13290 6557 13362
rect 6735 13290 6741 13362
rect 6551 13238 6552 13290
rect 6740 13238 6741 13290
rect 6551 13226 6557 13238
rect 6735 13226 6741 13238
rect 6551 13174 6552 13226
rect 6740 13174 6741 13226
rect 6551 13162 6557 13174
rect 6735 13162 6741 13174
rect 6551 13110 6552 13162
rect 6740 13110 6741 13162
rect 6551 13098 6557 13110
rect 6735 13098 6741 13110
rect 6551 13046 6552 13098
rect 6740 13046 6741 13098
rect 6551 13034 6557 13046
rect 6735 13034 6741 13046
rect 6551 12982 6552 13034
rect 6740 12982 6741 13034
rect 6551 12970 6557 12982
rect 6735 12970 6741 12982
rect 6551 12918 6552 12970
rect 6740 12918 6741 12970
rect 6551 12906 6557 12918
rect 6735 12906 6741 12918
rect 6551 12854 6552 12906
rect 6740 12854 6741 12906
rect 6551 12842 6557 12854
rect 6735 12842 6741 12854
rect 6551 12790 6552 12842
rect 6740 12790 6741 12842
rect 6551 12778 6557 12790
rect 6735 12778 6741 12790
rect 6551 12726 6552 12778
rect 6740 12726 6741 12778
rect 6551 12714 6557 12726
rect 6735 12714 6741 12726
rect 6551 12662 6552 12714
rect 6740 12662 6741 12714
rect 6551 12650 6557 12662
rect 6735 12650 6741 12662
rect 6551 12598 6552 12650
rect 6740 12598 6741 12650
rect 6551 12586 6557 12598
rect 6735 12586 6741 12598
rect 6551 12534 6552 12586
rect 6740 12534 6741 12586
rect 6551 12522 6557 12534
rect 6735 12522 6741 12534
rect 6551 12470 6552 12522
rect 6740 12470 6741 12522
rect 6551 12458 6557 12470
rect 6735 12458 6741 12470
rect 6551 12406 6552 12458
rect 6740 12406 6741 12458
rect 6551 12394 6557 12406
rect 6735 12394 6741 12406
rect 6551 12342 6552 12394
rect 6740 12342 6741 12394
rect 6551 12329 6557 12342
rect 6735 12329 6741 12342
rect 6551 12277 6552 12329
rect 6740 12277 6741 12329
rect 6551 12264 6557 12277
rect 6735 12264 6741 12277
rect 6551 12212 6552 12264
rect 6740 12212 6741 12264
rect 6551 12199 6557 12212
rect 6735 12199 6741 12212
rect 6551 12147 6552 12199
rect 6740 12147 6741 12199
rect 6551 12134 6557 12147
rect 6735 12134 6741 12147
rect 6551 12082 6552 12134
rect 6740 12082 6741 12134
rect 6551 12069 6557 12082
rect 6735 12069 6741 12082
rect 6551 12017 6552 12069
rect 6740 12017 6741 12069
rect 6551 12004 6557 12017
rect 6735 12004 6741 12017
rect 6551 11952 6552 12004
rect 6740 11952 6741 12004
rect 6551 11939 6557 11952
rect 6735 11939 6741 11952
rect 6551 11887 6552 11939
rect 6740 11887 6741 11939
rect 6551 11874 6557 11887
rect 6735 11874 6741 11887
rect 6551 11822 6552 11874
rect 6740 11822 6741 11874
rect 6551 11809 6557 11822
rect 6735 11809 6741 11822
rect 6551 11757 6552 11809
rect 6740 11757 6741 11809
rect 6551 11744 6557 11757
rect 6735 11744 6741 11757
rect 6551 11692 6552 11744
rect 6740 11692 6741 11744
rect 6551 11679 6557 11692
rect 6735 11679 6741 11692
rect 6551 11627 6552 11679
rect 6740 11627 6741 11679
rect 6551 11614 6557 11627
rect 6735 11614 6741 11627
rect 6551 11562 6552 11614
rect 6740 11562 6741 11614
rect 6551 10160 6557 11562
rect 6735 10160 6741 11562
rect 6551 10121 6741 10160
rect 6551 10087 6557 10121
rect 6591 10087 6629 10121
rect 6663 10087 6701 10121
rect 6735 10087 6741 10121
rect 6551 10048 6741 10087
rect 6551 10014 6557 10048
rect 6591 10014 6629 10048
rect 6663 10014 6701 10048
rect 6735 10014 6741 10048
rect 6551 9975 6741 10014
rect 6551 9941 6557 9975
rect 6591 9941 6629 9975
rect 6663 9941 6701 9975
rect 6735 9941 6741 9975
rect 6551 9902 6741 9941
rect 6551 9868 6557 9902
rect 6591 9868 6629 9902
rect 6663 9868 6701 9902
rect 6735 9868 6741 9902
rect 6551 9829 6741 9868
rect 6551 9795 6557 9829
rect 6591 9795 6629 9829
rect 6663 9795 6701 9829
rect 6735 9795 6741 9829
rect 6551 9756 6741 9795
rect 6551 9722 6557 9756
rect 6591 9722 6629 9756
rect 6663 9722 6701 9756
rect 6735 9722 6741 9756
rect 6551 9683 6741 9722
rect 6551 9649 6557 9683
rect 6591 9649 6629 9683
rect 6663 9649 6701 9683
rect 6735 9649 6741 9683
rect 6551 9610 6741 9649
rect 6551 9576 6557 9610
rect 6591 9576 6629 9610
rect 6663 9576 6701 9610
rect 6735 9576 6741 9610
rect 6551 9537 6741 9576
rect 6551 9503 6557 9537
rect 6591 9503 6629 9537
rect 6663 9503 6701 9537
rect 6735 9503 6741 9537
rect 6551 9491 6741 9503
rect 7041 37997 7171 38003
rect 7093 37945 7119 37997
rect 7041 37929 7171 37945
rect 7093 37877 7119 37929
rect 7041 37861 7171 37877
rect 7093 37809 7119 37861
rect 7041 37793 7171 37809
rect 7093 37741 7119 37793
rect 7041 37725 7171 37741
rect 7093 37673 7119 37725
rect 7041 37657 7171 37673
rect 7093 37605 7119 37657
rect 7041 37589 7171 37605
rect 7093 37537 7119 37589
rect 7041 37521 7171 37537
rect 7093 37469 7119 37521
rect 7041 37453 7171 37469
rect 7093 37401 7119 37453
rect 7041 37385 7171 37401
rect 7093 37333 7119 37385
rect 7041 37318 7171 37333
rect 7093 37266 7119 37318
rect 7041 37251 7171 37266
rect 7093 37199 7119 37251
rect 7041 37184 7171 37199
rect 7093 37132 7119 37184
rect 7041 37117 7171 37132
rect 7093 37065 7119 37117
rect 7041 34225 7171 37065
rect 7093 34173 7119 34225
rect 7041 34161 7171 34173
rect 7093 34109 7119 34161
rect 7041 34097 7171 34109
rect 7093 34045 7119 34097
rect 7041 34033 7171 34045
rect 7093 33981 7119 34033
rect 7041 33969 7171 33981
rect 7093 33917 7119 33969
rect 7041 33905 7171 33917
rect 7093 33853 7119 33905
rect 7041 33841 7171 33853
rect 7093 33789 7119 33841
rect 7041 33777 7171 33789
rect 7093 33725 7119 33777
rect 7041 33713 7171 33725
rect 7093 33661 7119 33713
rect 7041 33649 7171 33661
rect 7093 33597 7119 33649
rect 7041 33585 7171 33597
rect 7093 33533 7119 33585
rect 7041 33521 7171 33533
rect 7093 33469 7119 33521
rect 7041 33457 7171 33469
rect 7093 33405 7119 33457
rect 7041 33393 7171 33405
rect 7093 33341 7119 33393
rect 7041 33329 7171 33341
rect 7093 33277 7119 33329
rect 7041 33264 7171 33277
rect 7093 33212 7119 33264
rect 7041 33199 7171 33212
rect 7093 33147 7119 33199
rect 7041 33134 7171 33147
rect 7093 33082 7119 33134
rect 7041 33069 7171 33082
rect 7093 33017 7119 33069
rect 7041 33004 7171 33017
rect 7093 32952 7119 33004
rect 7041 32939 7171 32952
rect 7093 32887 7119 32939
rect 7041 32874 7171 32887
rect 7093 32822 7119 32874
rect 7041 32809 7171 32822
rect 7093 32757 7119 32809
rect 7041 32744 7171 32757
rect 7093 32692 7119 32744
rect 7041 32679 7171 32692
rect 7093 32627 7119 32679
rect 7041 32614 7171 32627
rect 7093 32562 7119 32614
rect 7041 32549 7171 32562
rect 7093 32497 7119 32549
rect 7041 29625 7171 32497
rect 7093 29573 7119 29625
rect 7041 29561 7171 29573
rect 7093 29509 7119 29561
rect 7041 29497 7171 29509
rect 7093 29445 7119 29497
rect 7041 29433 7171 29445
rect 7093 29381 7119 29433
rect 7041 29369 7171 29381
rect 7093 29317 7119 29369
rect 7041 29305 7171 29317
rect 7093 29253 7119 29305
rect 7041 29241 7171 29253
rect 7093 29189 7119 29241
rect 7041 29177 7171 29189
rect 7093 29125 7119 29177
rect 7041 29113 7171 29125
rect 7093 29061 7119 29113
rect 7041 29049 7171 29061
rect 7093 28997 7119 29049
rect 7041 28985 7171 28997
rect 7093 28933 7119 28985
rect 7041 28921 7171 28933
rect 7093 28869 7119 28921
rect 7041 28857 7171 28869
rect 7093 28805 7119 28857
rect 7041 28793 7171 28805
rect 7093 28741 7119 28793
rect 7041 28729 7171 28741
rect 7093 28677 7119 28729
rect 7041 28664 7171 28677
rect 7093 28612 7119 28664
rect 7041 28599 7171 28612
rect 7093 28547 7119 28599
rect 7041 28534 7171 28547
rect 7093 28482 7119 28534
rect 7041 28469 7171 28482
rect 7093 28417 7119 28469
rect 7041 28404 7171 28417
rect 7093 28352 7119 28404
rect 7041 28339 7171 28352
rect 7093 28287 7119 28339
rect 7041 28274 7171 28287
rect 7093 28222 7119 28274
rect 7041 28209 7171 28222
rect 7093 28157 7119 28209
rect 7041 28144 7171 28157
rect 7093 28092 7119 28144
rect 7041 28079 7171 28092
rect 7093 28027 7119 28079
rect 7041 28014 7171 28027
rect 7093 27962 7119 28014
rect 7041 27949 7171 27962
rect 7093 27897 7119 27949
rect 7041 25025 7171 27897
rect 7093 24973 7119 25025
rect 7041 24961 7171 24973
rect 7093 24909 7119 24961
rect 7041 24897 7171 24909
rect 7093 24845 7119 24897
rect 7041 24833 7171 24845
rect 7093 24781 7119 24833
rect 7041 24769 7171 24781
rect 7093 24717 7119 24769
rect 7041 24705 7171 24717
rect 7093 24653 7119 24705
rect 7041 24641 7171 24653
rect 7093 24589 7119 24641
rect 7041 24577 7171 24589
rect 7093 24525 7119 24577
rect 7041 24513 7171 24525
rect 7093 24461 7119 24513
rect 7041 24449 7171 24461
rect 7093 24397 7119 24449
rect 7041 24385 7171 24397
rect 7093 24333 7119 24385
rect 7041 24321 7171 24333
rect 7093 24269 7119 24321
rect 7041 24257 7171 24269
rect 7093 24205 7119 24257
rect 7041 24193 7171 24205
rect 7093 24141 7119 24193
rect 7041 24129 7171 24141
rect 7093 24077 7119 24129
rect 7041 24064 7171 24077
rect 7093 24012 7119 24064
rect 7041 23999 7171 24012
rect 7093 23947 7119 23999
rect 7041 23934 7171 23947
rect 7093 23882 7119 23934
rect 7041 23869 7171 23882
rect 7093 23817 7119 23869
rect 7041 23804 7171 23817
rect 7093 23752 7119 23804
rect 7041 23739 7171 23752
rect 7093 23687 7119 23739
rect 7041 23674 7171 23687
rect 7093 23622 7119 23674
rect 7041 23609 7171 23622
rect 7093 23557 7119 23609
rect 7041 23544 7171 23557
rect 7093 23492 7119 23544
rect 7041 23479 7171 23492
rect 7093 23427 7119 23479
rect 7041 23414 7171 23427
rect 7093 23362 7119 23414
rect 7041 23349 7171 23362
rect 7093 23297 7119 23349
rect 7041 20425 7171 23297
rect 7093 20373 7119 20425
rect 7041 20361 7171 20373
rect 7093 20309 7119 20361
rect 7041 20297 7171 20309
rect 7093 20245 7119 20297
rect 7041 20233 7171 20245
rect 7093 20181 7119 20233
rect 7041 20169 7171 20181
rect 7093 20117 7119 20169
rect 7041 20105 7171 20117
rect 7093 20053 7119 20105
rect 7041 20041 7171 20053
rect 7093 19989 7119 20041
rect 7041 19977 7171 19989
rect 7093 19925 7119 19977
rect 7041 19913 7171 19925
rect 7093 19861 7119 19913
rect 7041 19849 7171 19861
rect 7093 19797 7119 19849
rect 7041 19785 7171 19797
rect 7093 19733 7119 19785
rect 7041 19721 7171 19733
rect 7093 19669 7119 19721
rect 7041 19657 7171 19669
rect 7093 19605 7119 19657
rect 7041 19593 7171 19605
rect 7093 19541 7119 19593
rect 7041 19529 7171 19541
rect 7093 19477 7119 19529
rect 7041 19464 7171 19477
rect 7093 19412 7119 19464
rect 7041 19399 7171 19412
rect 7093 19347 7119 19399
rect 7041 19334 7171 19347
rect 7093 19282 7119 19334
rect 7041 19269 7171 19282
rect 7093 19217 7119 19269
rect 7041 19204 7171 19217
rect 7093 19152 7119 19204
rect 7041 19139 7171 19152
rect 7093 19087 7119 19139
rect 7041 19074 7171 19087
rect 7093 19022 7119 19074
rect 7041 19009 7171 19022
rect 7093 18957 7119 19009
rect 7041 18944 7171 18957
rect 7093 18892 7119 18944
rect 7041 18879 7171 18892
rect 7093 18827 7119 18879
rect 7041 18814 7171 18827
rect 7093 18762 7119 18814
rect 7041 18749 7171 18762
rect 7093 18697 7119 18749
rect 7041 15825 7171 18697
rect 7093 15773 7119 15825
rect 7041 15761 7171 15773
rect 7093 15709 7119 15761
rect 7041 15697 7171 15709
rect 7093 15645 7119 15697
rect 7041 15633 7171 15645
rect 7093 15581 7119 15633
rect 7041 15569 7171 15581
rect 7093 15517 7119 15569
rect 7041 15505 7171 15517
rect 7093 15453 7119 15505
rect 7041 15441 7171 15453
rect 7093 15389 7119 15441
rect 7041 15377 7171 15389
rect 7093 15325 7119 15377
rect 7041 15313 7171 15325
rect 7093 15261 7119 15313
rect 7041 15249 7171 15261
rect 7093 15197 7119 15249
rect 7041 15185 7171 15197
rect 7093 15133 7119 15185
rect 7041 15121 7171 15133
rect 7093 15069 7119 15121
rect 7041 15057 7171 15069
rect 7093 15005 7119 15057
rect 7041 14993 7171 15005
rect 7093 14941 7119 14993
rect 7041 14929 7171 14941
rect 7093 14877 7119 14929
rect 7041 14864 7171 14877
rect 7093 14812 7119 14864
rect 7041 14799 7171 14812
rect 7093 14747 7119 14799
rect 7041 14734 7171 14747
rect 7093 14682 7119 14734
rect 7041 14669 7171 14682
rect 7093 14617 7119 14669
rect 7041 14604 7171 14617
rect 7093 14552 7119 14604
rect 7041 14539 7171 14552
rect 7093 14487 7119 14539
rect 7041 14474 7171 14487
rect 7093 14422 7119 14474
rect 7041 14409 7171 14422
rect 7093 14357 7119 14409
rect 7041 14344 7171 14357
rect 7093 14292 7119 14344
rect 7041 14279 7171 14292
rect 7093 14227 7119 14279
rect 7041 14214 7171 14227
rect 7093 14162 7119 14214
rect 7041 14149 7171 14162
rect 7093 14097 7119 14149
rect 7041 11225 7171 14097
rect 7093 11173 7119 11225
rect 7041 11161 7171 11173
rect 7093 11109 7119 11161
rect 7041 11097 7171 11109
rect 7093 11045 7119 11097
rect 7041 11033 7171 11045
rect 7093 10981 7119 11033
rect 7041 10969 7171 10981
rect 7093 10917 7119 10969
rect 7041 10905 7171 10917
rect 7093 10853 7119 10905
rect 7041 10841 7171 10853
rect 7093 10789 7119 10841
rect 7041 10777 7171 10789
rect 7093 10725 7119 10777
rect 7041 10713 7171 10725
rect 7093 10661 7119 10713
rect 7041 10649 7171 10661
rect 7093 10597 7119 10649
rect 7041 10585 7171 10597
rect 7093 10533 7119 10585
rect 7041 10521 7171 10533
rect 7093 10469 7119 10521
rect 7041 10457 7171 10469
rect 7093 10405 7119 10457
rect 7041 10393 7171 10405
rect 7093 10341 7119 10393
rect 7041 10329 7171 10341
rect 7093 10277 7119 10329
rect 7041 10264 7171 10277
rect 7093 10212 7119 10264
rect 7041 10199 7171 10212
rect 7093 10147 7119 10199
rect 7041 10134 7171 10147
rect 7093 10082 7119 10134
rect 7041 10069 7171 10082
rect 7093 10017 7119 10069
rect 7041 10004 7171 10017
rect 7093 9952 7119 10004
rect 7041 9939 7171 9952
rect 7093 9887 7119 9939
rect 7041 9874 7171 9887
rect 7093 9822 7119 9874
rect 7041 9809 7171 9822
rect 7093 9757 7119 9809
rect 7041 9744 7171 9757
rect 7093 9692 7119 9744
rect 7041 9679 7171 9692
rect 7093 9627 7119 9679
rect 7041 9614 7171 9627
rect 7093 9562 7119 9614
rect 7041 9549 7171 9562
rect 7093 9497 7119 9549
rect 7041 9491 7171 9497
rect 7471 37962 7661 38003
rect 7471 37928 7477 37962
rect 7511 37928 7549 37962
rect 7583 37928 7621 37962
rect 7655 37928 7661 37962
rect 7471 37887 7661 37928
rect 7471 37853 7477 37887
rect 7511 37853 7549 37887
rect 7583 37853 7621 37887
rect 7655 37853 7661 37887
rect 7471 37812 7661 37853
rect 7471 37778 7477 37812
rect 7511 37778 7549 37812
rect 7583 37778 7621 37812
rect 7655 37778 7661 37812
rect 7471 37737 7661 37778
rect 7471 37703 7477 37737
rect 7511 37703 7549 37737
rect 7583 37703 7621 37737
rect 7655 37703 7661 37737
rect 7471 37662 7661 37703
rect 7471 37628 7477 37662
rect 7511 37628 7549 37662
rect 7583 37628 7621 37662
rect 7655 37628 7661 37662
rect 7471 37587 7661 37628
rect 7471 37553 7477 37587
rect 7511 37553 7549 37587
rect 7583 37553 7621 37587
rect 7655 37553 7661 37587
rect 7471 37512 7661 37553
rect 7471 37478 7477 37512
rect 7511 37478 7549 37512
rect 7583 37478 7621 37512
rect 7655 37478 7661 37512
rect 7471 37437 7661 37478
rect 7471 37403 7477 37437
rect 7511 37403 7549 37437
rect 7583 37403 7621 37437
rect 7655 37403 7661 37437
rect 7471 37362 7661 37403
rect 7471 37328 7477 37362
rect 7511 37328 7549 37362
rect 7583 37328 7621 37362
rect 7655 37328 7661 37362
rect 7471 37287 7661 37328
rect 7471 37253 7477 37287
rect 7511 37253 7549 37287
rect 7583 37253 7621 37287
rect 7655 37253 7661 37287
rect 7471 37212 7661 37253
rect 7471 37178 7477 37212
rect 7511 37178 7549 37212
rect 7583 37178 7621 37212
rect 7655 37178 7661 37212
rect 7471 37137 7661 37178
rect 7471 37103 7477 37137
rect 7511 37103 7549 37137
rect 7583 37103 7621 37137
rect 7655 37103 7661 37137
rect 7471 36353 7661 37103
rect 7471 36290 7477 36353
rect 7655 36290 7661 36353
rect 7471 36238 7472 36290
rect 7660 36238 7661 36290
rect 7471 36226 7477 36238
rect 7655 36226 7661 36238
rect 7471 36174 7472 36226
rect 7660 36174 7661 36226
rect 7471 36162 7477 36174
rect 7655 36162 7661 36174
rect 7471 36110 7472 36162
rect 7660 36110 7661 36162
rect 7471 36098 7477 36110
rect 7655 36098 7661 36110
rect 7471 36046 7472 36098
rect 7660 36046 7661 36098
rect 7471 36034 7477 36046
rect 7655 36034 7661 36046
rect 7471 35982 7472 36034
rect 7660 35982 7661 36034
rect 7471 35970 7477 35982
rect 7655 35970 7661 35982
rect 7471 35918 7472 35970
rect 7660 35918 7661 35970
rect 7471 35906 7477 35918
rect 7655 35906 7661 35918
rect 7471 35854 7472 35906
rect 7660 35854 7661 35906
rect 7471 35842 7477 35854
rect 7655 35842 7661 35854
rect 7471 35790 7472 35842
rect 7660 35790 7661 35842
rect 7471 35778 7477 35790
rect 7655 35778 7661 35790
rect 7471 35726 7472 35778
rect 7660 35726 7661 35778
rect 7471 35714 7477 35726
rect 7655 35714 7661 35726
rect 7471 35662 7472 35714
rect 7660 35662 7661 35714
rect 7471 35650 7477 35662
rect 7655 35650 7661 35662
rect 7471 35598 7472 35650
rect 7660 35598 7661 35650
rect 7471 35586 7477 35598
rect 7655 35586 7661 35598
rect 7471 35534 7472 35586
rect 7660 35534 7661 35586
rect 7471 35522 7477 35534
rect 7655 35522 7661 35534
rect 7471 35470 7472 35522
rect 7660 35470 7661 35522
rect 7471 35458 7477 35470
rect 7655 35458 7661 35470
rect 7471 35406 7472 35458
rect 7660 35406 7661 35458
rect 7471 35394 7477 35406
rect 7655 35394 7661 35406
rect 7471 35342 7472 35394
rect 7660 35342 7661 35394
rect 7471 35329 7477 35342
rect 7655 35329 7661 35342
rect 7471 35277 7472 35329
rect 7660 35277 7661 35329
rect 7471 35264 7477 35277
rect 7655 35264 7661 35277
rect 7471 35212 7472 35264
rect 7660 35212 7661 35264
rect 7471 35199 7477 35212
rect 7655 35199 7661 35212
rect 7471 35147 7472 35199
rect 7660 35147 7661 35199
rect 7471 35134 7477 35147
rect 7655 35134 7661 35147
rect 7471 35082 7472 35134
rect 7660 35082 7661 35134
rect 7471 35069 7477 35082
rect 7655 35069 7661 35082
rect 7471 35017 7472 35069
rect 7660 35017 7661 35069
rect 7471 35004 7477 35017
rect 7655 35004 7661 35017
rect 7471 34952 7472 35004
rect 7660 34952 7661 35004
rect 7471 34939 7477 34952
rect 7655 34939 7661 34952
rect 7471 34887 7472 34939
rect 7660 34887 7661 34939
rect 7471 34874 7477 34887
rect 7655 34874 7661 34887
rect 7471 34822 7472 34874
rect 7660 34822 7661 34874
rect 7471 34809 7477 34822
rect 7655 34809 7661 34822
rect 7471 34757 7472 34809
rect 7660 34757 7661 34809
rect 7471 34744 7477 34757
rect 7655 34744 7661 34757
rect 7471 34692 7472 34744
rect 7660 34692 7661 34744
rect 7471 34679 7477 34692
rect 7655 34679 7661 34692
rect 7471 34627 7472 34679
rect 7660 34627 7661 34679
rect 7471 34614 7477 34627
rect 7655 34614 7661 34627
rect 7471 34562 7472 34614
rect 7660 34562 7661 34614
rect 7471 32503 7477 34562
rect 7655 32503 7661 34562
rect 7471 31753 7661 32503
rect 7471 31690 7477 31753
rect 7655 31690 7661 31753
rect 7471 31638 7472 31690
rect 7660 31638 7661 31690
rect 7471 31626 7477 31638
rect 7655 31626 7661 31638
rect 7471 31574 7472 31626
rect 7660 31574 7661 31626
rect 7471 31562 7477 31574
rect 7655 31562 7661 31574
rect 7471 31510 7472 31562
rect 7660 31510 7661 31562
rect 7471 31498 7477 31510
rect 7655 31498 7661 31510
rect 7471 31446 7472 31498
rect 7660 31446 7661 31498
rect 7471 31434 7477 31446
rect 7655 31434 7661 31446
rect 7471 31382 7472 31434
rect 7660 31382 7661 31434
rect 7471 31370 7477 31382
rect 7655 31370 7661 31382
rect 7471 31318 7472 31370
rect 7660 31318 7661 31370
rect 7471 31306 7477 31318
rect 7655 31306 7661 31318
rect 7471 31254 7472 31306
rect 7660 31254 7661 31306
rect 7471 31242 7477 31254
rect 7655 31242 7661 31254
rect 7471 31190 7472 31242
rect 7660 31190 7661 31242
rect 7471 31178 7477 31190
rect 7655 31178 7661 31190
rect 7471 31126 7472 31178
rect 7660 31126 7661 31178
rect 7471 31114 7477 31126
rect 7655 31114 7661 31126
rect 7471 31062 7472 31114
rect 7660 31062 7661 31114
rect 7471 31050 7477 31062
rect 7655 31050 7661 31062
rect 7471 30998 7472 31050
rect 7660 30998 7661 31050
rect 7471 30986 7477 30998
rect 7655 30986 7661 30998
rect 7471 30934 7472 30986
rect 7660 30934 7661 30986
rect 7471 30922 7477 30934
rect 7655 30922 7661 30934
rect 7471 30870 7472 30922
rect 7660 30870 7661 30922
rect 7471 30858 7477 30870
rect 7655 30858 7661 30870
rect 7471 30806 7472 30858
rect 7660 30806 7661 30858
rect 7471 30794 7477 30806
rect 7655 30794 7661 30806
rect 7471 30742 7472 30794
rect 7660 30742 7661 30794
rect 7471 30729 7477 30742
rect 7655 30729 7661 30742
rect 7471 30677 7472 30729
rect 7660 30677 7661 30729
rect 7471 30664 7477 30677
rect 7655 30664 7661 30677
rect 7471 30612 7472 30664
rect 7660 30612 7661 30664
rect 7471 30599 7477 30612
rect 7655 30599 7661 30612
rect 7471 30547 7472 30599
rect 7660 30547 7661 30599
rect 7471 30534 7477 30547
rect 7655 30534 7661 30547
rect 7471 30482 7472 30534
rect 7660 30482 7661 30534
rect 7471 30469 7477 30482
rect 7655 30469 7661 30482
rect 7471 30417 7472 30469
rect 7660 30417 7661 30469
rect 7471 30404 7477 30417
rect 7655 30404 7661 30417
rect 7471 30352 7472 30404
rect 7660 30352 7661 30404
rect 7471 30339 7477 30352
rect 7655 30339 7661 30352
rect 7471 30287 7472 30339
rect 7660 30287 7661 30339
rect 7471 30274 7477 30287
rect 7655 30274 7661 30287
rect 7471 30222 7472 30274
rect 7660 30222 7661 30274
rect 7471 30209 7477 30222
rect 7655 30209 7661 30222
rect 7471 30157 7472 30209
rect 7660 30157 7661 30209
rect 7471 30144 7477 30157
rect 7655 30144 7661 30157
rect 7471 30092 7472 30144
rect 7660 30092 7661 30144
rect 7471 30079 7477 30092
rect 7655 30079 7661 30092
rect 7471 30027 7472 30079
rect 7660 30027 7661 30079
rect 7471 30014 7477 30027
rect 7655 30014 7661 30027
rect 7471 29962 7472 30014
rect 7660 29962 7661 30014
rect 7471 27903 7477 29962
rect 7655 27903 7661 29962
rect 7471 27153 7661 27903
rect 7471 27090 7477 27153
rect 7655 27090 7661 27153
rect 7471 27038 7472 27090
rect 7660 27038 7661 27090
rect 7471 27026 7477 27038
rect 7655 27026 7661 27038
rect 7471 26974 7472 27026
rect 7660 26974 7661 27026
rect 7471 26962 7477 26974
rect 7655 26962 7661 26974
rect 7471 26910 7472 26962
rect 7660 26910 7661 26962
rect 7471 26898 7477 26910
rect 7655 26898 7661 26910
rect 7471 26846 7472 26898
rect 7660 26846 7661 26898
rect 7471 26834 7477 26846
rect 7655 26834 7661 26846
rect 7471 26782 7472 26834
rect 7660 26782 7661 26834
rect 7471 26770 7477 26782
rect 7655 26770 7661 26782
rect 7471 26718 7472 26770
rect 7660 26718 7661 26770
rect 7471 26706 7477 26718
rect 7655 26706 7661 26718
rect 7471 26654 7472 26706
rect 7660 26654 7661 26706
rect 7471 26642 7477 26654
rect 7655 26642 7661 26654
rect 7471 26590 7472 26642
rect 7660 26590 7661 26642
rect 7471 26578 7477 26590
rect 7655 26578 7661 26590
rect 7471 26526 7472 26578
rect 7660 26526 7661 26578
rect 7471 26514 7477 26526
rect 7655 26514 7661 26526
rect 7471 26462 7472 26514
rect 7660 26462 7661 26514
rect 7471 26450 7477 26462
rect 7655 26450 7661 26462
rect 7471 26398 7472 26450
rect 7660 26398 7661 26450
rect 7471 26386 7477 26398
rect 7655 26386 7661 26398
rect 7471 26334 7472 26386
rect 7660 26334 7661 26386
rect 7471 26322 7477 26334
rect 7655 26322 7661 26334
rect 7471 26270 7472 26322
rect 7660 26270 7661 26322
rect 7471 26258 7477 26270
rect 7655 26258 7661 26270
rect 7471 26206 7472 26258
rect 7660 26206 7661 26258
rect 7471 26194 7477 26206
rect 7655 26194 7661 26206
rect 7471 26142 7472 26194
rect 7660 26142 7661 26194
rect 7471 26129 7477 26142
rect 7655 26129 7661 26142
rect 7471 26077 7472 26129
rect 7660 26077 7661 26129
rect 7471 26064 7477 26077
rect 7655 26064 7661 26077
rect 7471 26012 7472 26064
rect 7660 26012 7661 26064
rect 7471 25999 7477 26012
rect 7655 25999 7661 26012
rect 7471 25947 7472 25999
rect 7660 25947 7661 25999
rect 7471 25934 7477 25947
rect 7655 25934 7661 25947
rect 7471 25882 7472 25934
rect 7660 25882 7661 25934
rect 7471 25869 7477 25882
rect 7655 25869 7661 25882
rect 7471 25817 7472 25869
rect 7660 25817 7661 25869
rect 7471 25804 7477 25817
rect 7655 25804 7661 25817
rect 7471 25752 7472 25804
rect 7660 25752 7661 25804
rect 7471 25739 7477 25752
rect 7655 25739 7661 25752
rect 7471 25687 7472 25739
rect 7660 25687 7661 25739
rect 7471 25674 7477 25687
rect 7655 25674 7661 25687
rect 7471 25622 7472 25674
rect 7660 25622 7661 25674
rect 7471 25609 7477 25622
rect 7655 25609 7661 25622
rect 7471 25557 7472 25609
rect 7660 25557 7661 25609
rect 7471 25544 7477 25557
rect 7655 25544 7661 25557
rect 7471 25492 7472 25544
rect 7660 25492 7661 25544
rect 7471 25479 7477 25492
rect 7655 25479 7661 25492
rect 7471 25427 7472 25479
rect 7660 25427 7661 25479
rect 7471 25414 7477 25427
rect 7655 25414 7661 25427
rect 7471 25362 7472 25414
rect 7660 25362 7661 25414
rect 7471 23303 7477 25362
rect 7655 23303 7661 25362
rect 7471 22562 7661 23303
rect 7471 22490 7477 22562
rect 7655 22490 7661 22562
rect 7471 22438 7472 22490
rect 7660 22438 7661 22490
rect 7471 22426 7477 22438
rect 7655 22426 7661 22438
rect 7471 22374 7472 22426
rect 7660 22374 7661 22426
rect 7471 22362 7477 22374
rect 7655 22362 7661 22374
rect 7471 22310 7472 22362
rect 7660 22310 7661 22362
rect 7471 22298 7477 22310
rect 7655 22298 7661 22310
rect 7471 22246 7472 22298
rect 7660 22246 7661 22298
rect 7471 22234 7477 22246
rect 7655 22234 7661 22246
rect 7471 22182 7472 22234
rect 7660 22182 7661 22234
rect 7471 22170 7477 22182
rect 7655 22170 7661 22182
rect 7471 22118 7472 22170
rect 7660 22118 7661 22170
rect 7471 22106 7477 22118
rect 7655 22106 7661 22118
rect 7471 22054 7472 22106
rect 7660 22054 7661 22106
rect 7471 22042 7477 22054
rect 7655 22042 7661 22054
rect 7471 21990 7472 22042
rect 7660 21990 7661 22042
rect 7471 21978 7477 21990
rect 7655 21978 7661 21990
rect 7471 21926 7472 21978
rect 7660 21926 7661 21978
rect 7471 21914 7477 21926
rect 7655 21914 7661 21926
rect 7471 21862 7472 21914
rect 7660 21862 7661 21914
rect 7471 21850 7477 21862
rect 7655 21850 7661 21862
rect 7471 21798 7472 21850
rect 7660 21798 7661 21850
rect 7471 21786 7477 21798
rect 7655 21786 7661 21798
rect 7471 21734 7472 21786
rect 7660 21734 7661 21786
rect 7471 21722 7477 21734
rect 7655 21722 7661 21734
rect 7471 21670 7472 21722
rect 7660 21670 7661 21722
rect 7471 21658 7477 21670
rect 7655 21658 7661 21670
rect 7471 21606 7472 21658
rect 7660 21606 7661 21658
rect 7471 21594 7477 21606
rect 7655 21594 7661 21606
rect 7471 21542 7472 21594
rect 7660 21542 7661 21594
rect 7471 21529 7477 21542
rect 7655 21529 7661 21542
rect 7471 21477 7472 21529
rect 7660 21477 7661 21529
rect 7471 21464 7477 21477
rect 7655 21464 7661 21477
rect 7471 21412 7472 21464
rect 7660 21412 7661 21464
rect 7471 21399 7477 21412
rect 7655 21399 7661 21412
rect 7471 21347 7472 21399
rect 7660 21347 7661 21399
rect 7471 21334 7477 21347
rect 7655 21334 7661 21347
rect 7471 21282 7472 21334
rect 7660 21282 7661 21334
rect 7471 21269 7477 21282
rect 7655 21269 7661 21282
rect 7471 21217 7472 21269
rect 7660 21217 7661 21269
rect 7471 21204 7477 21217
rect 7655 21204 7661 21217
rect 7471 21152 7472 21204
rect 7660 21152 7661 21204
rect 7471 21139 7477 21152
rect 7655 21139 7661 21152
rect 7471 21087 7472 21139
rect 7660 21087 7661 21139
rect 7471 21074 7477 21087
rect 7655 21074 7661 21087
rect 7471 21022 7472 21074
rect 7660 21022 7661 21074
rect 7471 21009 7477 21022
rect 7655 21009 7661 21022
rect 7471 20957 7472 21009
rect 7660 20957 7661 21009
rect 7471 20944 7477 20957
rect 7655 20944 7661 20957
rect 7471 20892 7472 20944
rect 7660 20892 7661 20944
rect 7471 20879 7477 20892
rect 7655 20879 7661 20892
rect 7471 20827 7472 20879
rect 7660 20827 7661 20879
rect 7471 20814 7477 20827
rect 7655 20814 7661 20827
rect 7471 20762 7472 20814
rect 7660 20762 7661 20814
rect 7471 19360 7477 20762
rect 7655 19360 7661 20762
rect 7471 19321 7661 19360
rect 7471 19287 7477 19321
rect 7511 19287 7549 19321
rect 7583 19287 7621 19321
rect 7655 19287 7661 19321
rect 7471 19248 7661 19287
rect 7471 19214 7477 19248
rect 7511 19214 7549 19248
rect 7583 19214 7621 19248
rect 7655 19214 7661 19248
rect 7471 19175 7661 19214
rect 7471 19141 7477 19175
rect 7511 19141 7549 19175
rect 7583 19141 7621 19175
rect 7655 19141 7661 19175
rect 7471 19102 7661 19141
rect 7471 19068 7477 19102
rect 7511 19068 7549 19102
rect 7583 19068 7621 19102
rect 7655 19068 7661 19102
rect 7471 19029 7661 19068
rect 7471 18995 7477 19029
rect 7511 18995 7549 19029
rect 7583 18995 7621 19029
rect 7655 18995 7661 19029
rect 7471 18956 7661 18995
rect 7471 18922 7477 18956
rect 7511 18922 7549 18956
rect 7583 18922 7621 18956
rect 7655 18922 7661 18956
rect 7471 18883 7661 18922
rect 7471 18849 7477 18883
rect 7511 18849 7549 18883
rect 7583 18849 7621 18883
rect 7655 18849 7661 18883
rect 7471 18810 7661 18849
rect 7471 18776 7477 18810
rect 7511 18776 7549 18810
rect 7583 18776 7621 18810
rect 7655 18776 7661 18810
rect 7471 18737 7661 18776
rect 7471 18703 7477 18737
rect 7511 18703 7549 18737
rect 7583 18703 7621 18737
rect 7655 18703 7661 18737
rect 7471 17953 7661 18703
rect 7471 17890 7477 17953
rect 7655 17890 7661 17953
rect 7471 17838 7472 17890
rect 7660 17838 7661 17890
rect 7471 17826 7477 17838
rect 7655 17826 7661 17838
rect 7471 17774 7472 17826
rect 7660 17774 7661 17826
rect 7471 17762 7477 17774
rect 7655 17762 7661 17774
rect 7471 17710 7472 17762
rect 7660 17710 7661 17762
rect 7471 17698 7477 17710
rect 7655 17698 7661 17710
rect 7471 17646 7472 17698
rect 7660 17646 7661 17698
rect 7471 17634 7477 17646
rect 7655 17634 7661 17646
rect 7471 17582 7472 17634
rect 7660 17582 7661 17634
rect 7471 17570 7477 17582
rect 7655 17570 7661 17582
rect 7471 17518 7472 17570
rect 7660 17518 7661 17570
rect 7471 17506 7477 17518
rect 7655 17506 7661 17518
rect 7471 17454 7472 17506
rect 7660 17454 7661 17506
rect 7471 17442 7477 17454
rect 7655 17442 7661 17454
rect 7471 17390 7472 17442
rect 7660 17390 7661 17442
rect 7471 17378 7477 17390
rect 7655 17378 7661 17390
rect 7471 17326 7472 17378
rect 7660 17326 7661 17378
rect 7471 17314 7477 17326
rect 7655 17314 7661 17326
rect 7471 17262 7472 17314
rect 7660 17262 7661 17314
rect 7471 17250 7477 17262
rect 7655 17250 7661 17262
rect 7471 17198 7472 17250
rect 7660 17198 7661 17250
rect 7471 17186 7477 17198
rect 7655 17186 7661 17198
rect 7471 17134 7472 17186
rect 7660 17134 7661 17186
rect 7471 17122 7477 17134
rect 7655 17122 7661 17134
rect 7471 17070 7472 17122
rect 7660 17070 7661 17122
rect 7471 17058 7477 17070
rect 7655 17058 7661 17070
rect 7471 17006 7472 17058
rect 7660 17006 7661 17058
rect 7471 16994 7477 17006
rect 7655 16994 7661 17006
rect 7471 16942 7472 16994
rect 7660 16942 7661 16994
rect 7471 16929 7477 16942
rect 7655 16929 7661 16942
rect 7471 16877 7472 16929
rect 7660 16877 7661 16929
rect 7471 16864 7477 16877
rect 7655 16864 7661 16877
rect 7471 16812 7472 16864
rect 7660 16812 7661 16864
rect 7471 16799 7477 16812
rect 7655 16799 7661 16812
rect 7471 16747 7472 16799
rect 7660 16747 7661 16799
rect 7471 16734 7477 16747
rect 7655 16734 7661 16747
rect 7471 16682 7472 16734
rect 7660 16682 7661 16734
rect 7471 16669 7477 16682
rect 7655 16669 7661 16682
rect 7471 16617 7472 16669
rect 7660 16617 7661 16669
rect 7471 16604 7477 16617
rect 7655 16604 7661 16617
rect 7471 16552 7472 16604
rect 7660 16552 7661 16604
rect 7471 16539 7477 16552
rect 7655 16539 7661 16552
rect 7471 16487 7472 16539
rect 7660 16487 7661 16539
rect 7471 16474 7477 16487
rect 7655 16474 7661 16487
rect 7471 16422 7472 16474
rect 7660 16422 7661 16474
rect 7471 16409 7477 16422
rect 7655 16409 7661 16422
rect 7471 16357 7472 16409
rect 7660 16357 7661 16409
rect 7471 16344 7477 16357
rect 7655 16344 7661 16357
rect 7471 16292 7472 16344
rect 7660 16292 7661 16344
rect 7471 16279 7477 16292
rect 7655 16279 7661 16292
rect 7471 16227 7472 16279
rect 7660 16227 7661 16279
rect 7471 16214 7477 16227
rect 7655 16214 7661 16227
rect 7471 16162 7472 16214
rect 7660 16162 7661 16214
rect 7471 14103 7477 16162
rect 7655 14103 7661 16162
rect 7471 13362 7661 14103
rect 7471 13290 7477 13362
rect 7655 13290 7661 13362
rect 7471 13238 7472 13290
rect 7660 13238 7661 13290
rect 7471 13226 7477 13238
rect 7655 13226 7661 13238
rect 7471 13174 7472 13226
rect 7660 13174 7661 13226
rect 7471 13162 7477 13174
rect 7655 13162 7661 13174
rect 7471 13110 7472 13162
rect 7660 13110 7661 13162
rect 7471 13098 7477 13110
rect 7655 13098 7661 13110
rect 7471 13046 7472 13098
rect 7660 13046 7661 13098
rect 7471 13034 7477 13046
rect 7655 13034 7661 13046
rect 7471 12982 7472 13034
rect 7660 12982 7661 13034
rect 7471 12970 7477 12982
rect 7655 12970 7661 12982
rect 7471 12918 7472 12970
rect 7660 12918 7661 12970
rect 7471 12906 7477 12918
rect 7655 12906 7661 12918
rect 7471 12854 7472 12906
rect 7660 12854 7661 12906
rect 7471 12842 7477 12854
rect 7655 12842 7661 12854
rect 7471 12790 7472 12842
rect 7660 12790 7661 12842
rect 7471 12778 7477 12790
rect 7655 12778 7661 12790
rect 7471 12726 7472 12778
rect 7660 12726 7661 12778
rect 7471 12714 7477 12726
rect 7655 12714 7661 12726
rect 7471 12662 7472 12714
rect 7660 12662 7661 12714
rect 7471 12650 7477 12662
rect 7655 12650 7661 12662
rect 7471 12598 7472 12650
rect 7660 12598 7661 12650
rect 7471 12586 7477 12598
rect 7655 12586 7661 12598
rect 7471 12534 7472 12586
rect 7660 12534 7661 12586
rect 7471 12522 7477 12534
rect 7655 12522 7661 12534
rect 7471 12470 7472 12522
rect 7660 12470 7661 12522
rect 7471 12458 7477 12470
rect 7655 12458 7661 12470
rect 7471 12406 7472 12458
rect 7660 12406 7661 12458
rect 7471 12394 7477 12406
rect 7655 12394 7661 12406
rect 7471 12342 7472 12394
rect 7660 12342 7661 12394
rect 7471 12329 7477 12342
rect 7655 12329 7661 12342
rect 7471 12277 7472 12329
rect 7660 12277 7661 12329
rect 7471 12264 7477 12277
rect 7655 12264 7661 12277
rect 7471 12212 7472 12264
rect 7660 12212 7661 12264
rect 7471 12199 7477 12212
rect 7655 12199 7661 12212
rect 7471 12147 7472 12199
rect 7660 12147 7661 12199
rect 7471 12134 7477 12147
rect 7655 12134 7661 12147
rect 7471 12082 7472 12134
rect 7660 12082 7661 12134
rect 7471 12069 7477 12082
rect 7655 12069 7661 12082
rect 7471 12017 7472 12069
rect 7660 12017 7661 12069
rect 7471 12004 7477 12017
rect 7655 12004 7661 12017
rect 7471 11952 7472 12004
rect 7660 11952 7661 12004
rect 7471 11939 7477 11952
rect 7655 11939 7661 11952
rect 7471 11887 7472 11939
rect 7660 11887 7661 11939
rect 7471 11874 7477 11887
rect 7655 11874 7661 11887
rect 7471 11822 7472 11874
rect 7660 11822 7661 11874
rect 7471 11809 7477 11822
rect 7655 11809 7661 11822
rect 7471 11757 7472 11809
rect 7660 11757 7661 11809
rect 7471 11744 7477 11757
rect 7655 11744 7661 11757
rect 7471 11692 7472 11744
rect 7660 11692 7661 11744
rect 7471 11679 7477 11692
rect 7655 11679 7661 11692
rect 7471 11627 7472 11679
rect 7660 11627 7661 11679
rect 7471 11614 7477 11627
rect 7655 11614 7661 11627
rect 7471 11562 7472 11614
rect 7660 11562 7661 11614
rect 7471 10160 7477 11562
rect 7655 10160 7661 11562
rect 7471 10121 7661 10160
rect 7471 10087 7477 10121
rect 7511 10087 7549 10121
rect 7583 10087 7621 10121
rect 7655 10087 7661 10121
rect 7471 10048 7661 10087
rect 7471 10014 7477 10048
rect 7511 10014 7549 10048
rect 7583 10014 7621 10048
rect 7655 10014 7661 10048
rect 7471 9975 7661 10014
rect 7471 9941 7477 9975
rect 7511 9941 7549 9975
rect 7583 9941 7621 9975
rect 7655 9941 7661 9975
rect 7471 9902 7661 9941
rect 7471 9868 7477 9902
rect 7511 9868 7549 9902
rect 7583 9868 7621 9902
rect 7655 9868 7661 9902
rect 7471 9829 7661 9868
rect 7471 9795 7477 9829
rect 7511 9795 7549 9829
rect 7583 9795 7621 9829
rect 7655 9795 7661 9829
rect 7471 9756 7661 9795
rect 7471 9722 7477 9756
rect 7511 9722 7549 9756
rect 7583 9722 7621 9756
rect 7655 9722 7661 9756
rect 7471 9683 7661 9722
rect 7471 9649 7477 9683
rect 7511 9649 7549 9683
rect 7583 9649 7621 9683
rect 7655 9649 7661 9683
rect 7471 9610 7661 9649
rect 7471 9576 7477 9610
rect 7511 9576 7549 9610
rect 7583 9576 7621 9610
rect 7655 9576 7661 9610
rect 7471 9537 7661 9576
rect 7471 9503 7477 9537
rect 7511 9503 7549 9537
rect 7583 9503 7621 9537
rect 7655 9503 7661 9537
rect 7471 9491 7661 9503
rect 7961 37997 8091 38003
rect 8013 37945 8039 37997
rect 7961 37929 8091 37945
rect 8013 37877 8039 37929
rect 7961 37861 8091 37877
rect 8013 37809 8039 37861
rect 7961 37793 8091 37809
rect 8013 37741 8039 37793
rect 7961 37725 8091 37741
rect 8013 37673 8039 37725
rect 7961 37657 8091 37673
rect 8013 37605 8039 37657
rect 7961 37589 8091 37605
rect 8013 37537 8039 37589
rect 7961 37521 8091 37537
rect 8013 37469 8039 37521
rect 7961 37453 8091 37469
rect 8013 37401 8039 37453
rect 7961 37385 8091 37401
rect 8013 37333 8039 37385
rect 7961 37318 8091 37333
rect 8013 37266 8039 37318
rect 7961 37251 8091 37266
rect 8013 37199 8039 37251
rect 7961 37184 8091 37199
rect 8013 37132 8039 37184
rect 7961 37117 8091 37132
rect 8013 37065 8039 37117
rect 7961 34225 8091 37065
rect 8013 34173 8039 34225
rect 7961 34161 8091 34173
rect 8013 34109 8039 34161
rect 7961 34097 8091 34109
rect 8013 34045 8039 34097
rect 7961 34033 8091 34045
rect 8013 33981 8039 34033
rect 7961 33969 8091 33981
rect 8013 33917 8039 33969
rect 7961 33905 8091 33917
rect 8013 33853 8039 33905
rect 7961 33841 8091 33853
rect 8013 33789 8039 33841
rect 7961 33777 8091 33789
rect 8013 33725 8039 33777
rect 7961 33713 8091 33725
rect 8013 33661 8039 33713
rect 7961 33649 8091 33661
rect 8013 33597 8039 33649
rect 7961 33585 8091 33597
rect 8013 33533 8039 33585
rect 7961 33521 8091 33533
rect 8013 33469 8039 33521
rect 7961 33457 8091 33469
rect 8013 33405 8039 33457
rect 7961 33393 8091 33405
rect 8013 33341 8039 33393
rect 7961 33329 8091 33341
rect 8013 33277 8039 33329
rect 7961 33264 8091 33277
rect 8013 33212 8039 33264
rect 7961 33199 8091 33212
rect 8013 33147 8039 33199
rect 7961 33134 8091 33147
rect 8013 33082 8039 33134
rect 7961 33069 8091 33082
rect 8013 33017 8039 33069
rect 7961 33004 8091 33017
rect 8013 32952 8039 33004
rect 7961 32939 8091 32952
rect 8013 32887 8039 32939
rect 7961 32874 8091 32887
rect 8013 32822 8039 32874
rect 7961 32809 8091 32822
rect 8013 32757 8039 32809
rect 7961 32744 8091 32757
rect 8013 32692 8039 32744
rect 7961 32679 8091 32692
rect 8013 32627 8039 32679
rect 7961 32614 8091 32627
rect 8013 32562 8039 32614
rect 7961 32549 8091 32562
rect 8013 32497 8039 32549
rect 7961 29625 8091 32497
rect 8013 29573 8039 29625
rect 7961 29561 8091 29573
rect 8013 29509 8039 29561
rect 7961 29497 8091 29509
rect 8013 29445 8039 29497
rect 7961 29433 8091 29445
rect 8013 29381 8039 29433
rect 7961 29369 8091 29381
rect 8013 29317 8039 29369
rect 7961 29305 8091 29317
rect 8013 29253 8039 29305
rect 7961 29241 8091 29253
rect 8013 29189 8039 29241
rect 7961 29177 8091 29189
rect 8013 29125 8039 29177
rect 7961 29113 8091 29125
rect 8013 29061 8039 29113
rect 7961 29049 8091 29061
rect 8013 28997 8039 29049
rect 7961 28985 8091 28997
rect 8013 28933 8039 28985
rect 7961 28921 8091 28933
rect 8013 28869 8039 28921
rect 7961 28857 8091 28869
rect 8013 28805 8039 28857
rect 7961 28793 8091 28805
rect 8013 28741 8039 28793
rect 7961 28729 8091 28741
rect 8013 28677 8039 28729
rect 7961 28664 8091 28677
rect 8013 28612 8039 28664
rect 7961 28599 8091 28612
rect 8013 28547 8039 28599
rect 7961 28534 8091 28547
rect 8013 28482 8039 28534
rect 7961 28469 8091 28482
rect 8013 28417 8039 28469
rect 7961 28404 8091 28417
rect 8013 28352 8039 28404
rect 7961 28339 8091 28352
rect 8013 28287 8039 28339
rect 7961 28274 8091 28287
rect 8013 28222 8039 28274
rect 7961 28209 8091 28222
rect 8013 28157 8039 28209
rect 7961 28144 8091 28157
rect 8013 28092 8039 28144
rect 7961 28079 8091 28092
rect 8013 28027 8039 28079
rect 7961 28014 8091 28027
rect 8013 27962 8039 28014
rect 7961 27949 8091 27962
rect 8013 27897 8039 27949
rect 7961 25025 8091 27897
rect 8013 24973 8039 25025
rect 7961 24961 8091 24973
rect 8013 24909 8039 24961
rect 7961 24897 8091 24909
rect 8013 24845 8039 24897
rect 7961 24833 8091 24845
rect 8013 24781 8039 24833
rect 7961 24769 8091 24781
rect 8013 24717 8039 24769
rect 7961 24705 8091 24717
rect 8013 24653 8039 24705
rect 7961 24641 8091 24653
rect 8013 24589 8039 24641
rect 7961 24577 8091 24589
rect 8013 24525 8039 24577
rect 7961 24513 8091 24525
rect 8013 24461 8039 24513
rect 7961 24449 8091 24461
rect 8013 24397 8039 24449
rect 7961 24385 8091 24397
rect 8013 24333 8039 24385
rect 7961 24321 8091 24333
rect 8013 24269 8039 24321
rect 7961 24257 8091 24269
rect 8013 24205 8039 24257
rect 7961 24193 8091 24205
rect 8013 24141 8039 24193
rect 7961 24129 8091 24141
rect 8013 24077 8039 24129
rect 7961 24064 8091 24077
rect 8013 24012 8039 24064
rect 7961 23999 8091 24012
rect 8013 23947 8039 23999
rect 7961 23934 8091 23947
rect 8013 23882 8039 23934
rect 7961 23869 8091 23882
rect 8013 23817 8039 23869
rect 7961 23804 8091 23817
rect 8013 23752 8039 23804
rect 7961 23739 8091 23752
rect 8013 23687 8039 23739
rect 7961 23674 8091 23687
rect 8013 23622 8039 23674
rect 7961 23609 8091 23622
rect 8013 23557 8039 23609
rect 7961 23544 8091 23557
rect 8013 23492 8039 23544
rect 7961 23479 8091 23492
rect 8013 23427 8039 23479
rect 7961 23414 8091 23427
rect 8013 23362 8039 23414
rect 7961 23349 8091 23362
rect 8013 23297 8039 23349
rect 7961 20425 8091 23297
rect 8013 20373 8039 20425
rect 7961 20361 8091 20373
rect 8013 20309 8039 20361
rect 7961 20297 8091 20309
rect 8013 20245 8039 20297
rect 7961 20233 8091 20245
rect 8013 20181 8039 20233
rect 7961 20169 8091 20181
rect 8013 20117 8039 20169
rect 7961 20105 8091 20117
rect 8013 20053 8039 20105
rect 7961 20041 8091 20053
rect 8013 19989 8039 20041
rect 7961 19977 8091 19989
rect 8013 19925 8039 19977
rect 7961 19913 8091 19925
rect 8013 19861 8039 19913
rect 7961 19849 8091 19861
rect 8013 19797 8039 19849
rect 7961 19785 8091 19797
rect 8013 19733 8039 19785
rect 7961 19721 8091 19733
rect 8013 19669 8039 19721
rect 7961 19657 8091 19669
rect 8013 19605 8039 19657
rect 7961 19593 8091 19605
rect 8013 19541 8039 19593
rect 7961 19529 8091 19541
rect 8013 19477 8039 19529
rect 7961 19464 8091 19477
rect 8013 19412 8039 19464
rect 7961 19399 8091 19412
rect 8013 19347 8039 19399
rect 7961 19334 8091 19347
rect 8013 19282 8039 19334
rect 7961 19269 8091 19282
rect 8013 19217 8039 19269
rect 7961 19204 8091 19217
rect 8013 19152 8039 19204
rect 7961 19139 8091 19152
rect 8013 19087 8039 19139
rect 7961 19074 8091 19087
rect 8013 19022 8039 19074
rect 7961 19009 8091 19022
rect 8013 18957 8039 19009
rect 7961 18944 8091 18957
rect 8013 18892 8039 18944
rect 7961 18879 8091 18892
rect 8013 18827 8039 18879
rect 7961 18814 8091 18827
rect 8013 18762 8039 18814
rect 7961 18749 8091 18762
rect 8013 18697 8039 18749
rect 7961 15825 8091 18697
rect 8013 15773 8039 15825
rect 7961 15761 8091 15773
rect 8013 15709 8039 15761
rect 7961 15697 8091 15709
rect 8013 15645 8039 15697
rect 7961 15633 8091 15645
rect 8013 15581 8039 15633
rect 7961 15569 8091 15581
rect 8013 15517 8039 15569
rect 7961 15505 8091 15517
rect 8013 15453 8039 15505
rect 7961 15441 8091 15453
rect 8013 15389 8039 15441
rect 7961 15377 8091 15389
rect 8013 15325 8039 15377
rect 7961 15313 8091 15325
rect 8013 15261 8039 15313
rect 7961 15249 8091 15261
rect 8013 15197 8039 15249
rect 7961 15185 8091 15197
rect 8013 15133 8039 15185
rect 7961 15121 8091 15133
rect 8013 15069 8039 15121
rect 7961 15057 8091 15069
rect 8013 15005 8039 15057
rect 7961 14993 8091 15005
rect 8013 14941 8039 14993
rect 7961 14929 8091 14941
rect 8013 14877 8039 14929
rect 7961 14864 8091 14877
rect 8013 14812 8039 14864
rect 7961 14799 8091 14812
rect 8013 14747 8039 14799
rect 7961 14734 8091 14747
rect 8013 14682 8039 14734
rect 7961 14669 8091 14682
rect 8013 14617 8039 14669
rect 7961 14604 8091 14617
rect 8013 14552 8039 14604
rect 7961 14539 8091 14552
rect 8013 14487 8039 14539
rect 7961 14474 8091 14487
rect 8013 14422 8039 14474
rect 7961 14409 8091 14422
rect 8013 14357 8039 14409
rect 7961 14344 8091 14357
rect 8013 14292 8039 14344
rect 7961 14279 8091 14292
rect 8013 14227 8039 14279
rect 7961 14214 8091 14227
rect 8013 14162 8039 14214
rect 7961 14149 8091 14162
rect 8013 14097 8039 14149
rect 7961 11225 8091 14097
rect 8013 11173 8039 11225
rect 7961 11161 8091 11173
rect 8013 11109 8039 11161
rect 7961 11097 8091 11109
rect 8013 11045 8039 11097
rect 7961 11033 8091 11045
rect 8013 10981 8039 11033
rect 7961 10969 8091 10981
rect 8013 10917 8039 10969
rect 7961 10905 8091 10917
rect 8013 10853 8039 10905
rect 7961 10841 8091 10853
rect 8013 10789 8039 10841
rect 7961 10777 8091 10789
rect 8013 10725 8039 10777
rect 7961 10713 8091 10725
rect 8013 10661 8039 10713
rect 7961 10649 8091 10661
rect 8013 10597 8039 10649
rect 7961 10585 8091 10597
rect 8013 10533 8039 10585
rect 7961 10521 8091 10533
rect 8013 10469 8039 10521
rect 7961 10457 8091 10469
rect 8013 10405 8039 10457
rect 7961 10393 8091 10405
rect 8013 10341 8039 10393
rect 7961 10329 8091 10341
rect 8013 10277 8039 10329
rect 7961 10264 8091 10277
rect 8013 10212 8039 10264
rect 7961 10199 8091 10212
rect 8013 10147 8039 10199
rect 7961 10134 8091 10147
rect 8013 10082 8039 10134
rect 7961 10069 8091 10082
rect 8013 10017 8039 10069
rect 7961 10004 8091 10017
rect 8013 9952 8039 10004
rect 7961 9939 8091 9952
rect 8013 9887 8039 9939
rect 7961 9874 8091 9887
rect 8013 9822 8039 9874
rect 7961 9809 8091 9822
rect 8013 9757 8039 9809
rect 7961 9744 8091 9757
rect 8013 9692 8039 9744
rect 7961 9679 8091 9692
rect 8013 9627 8039 9679
rect 7961 9614 8091 9627
rect 8013 9562 8039 9614
rect 7961 9549 8091 9562
rect 8013 9497 8039 9549
rect 7961 9491 8091 9497
rect 8391 37962 8581 38003
rect 8391 37928 8397 37962
rect 8431 37928 8469 37962
rect 8503 37928 8541 37962
rect 8575 37928 8581 37962
rect 8391 37887 8581 37928
rect 8391 37853 8397 37887
rect 8431 37853 8469 37887
rect 8503 37853 8541 37887
rect 8575 37853 8581 37887
rect 8391 37812 8581 37853
rect 8391 37778 8397 37812
rect 8431 37778 8469 37812
rect 8503 37778 8541 37812
rect 8575 37778 8581 37812
rect 8391 37737 8581 37778
rect 8391 37703 8397 37737
rect 8431 37703 8469 37737
rect 8503 37703 8541 37737
rect 8575 37703 8581 37737
rect 8391 37662 8581 37703
rect 8391 37628 8397 37662
rect 8431 37628 8469 37662
rect 8503 37628 8541 37662
rect 8575 37628 8581 37662
rect 8391 37587 8581 37628
rect 8391 37553 8397 37587
rect 8431 37553 8469 37587
rect 8503 37553 8541 37587
rect 8575 37553 8581 37587
rect 8391 37512 8581 37553
rect 8391 37478 8397 37512
rect 8431 37478 8469 37512
rect 8503 37478 8541 37512
rect 8575 37478 8581 37512
rect 8391 37437 8581 37478
rect 8391 37403 8397 37437
rect 8431 37403 8469 37437
rect 8503 37403 8541 37437
rect 8575 37403 8581 37437
rect 8391 37362 8581 37403
rect 8391 37328 8397 37362
rect 8431 37328 8469 37362
rect 8503 37328 8541 37362
rect 8575 37328 8581 37362
rect 8391 37287 8581 37328
rect 8391 37253 8397 37287
rect 8431 37253 8469 37287
rect 8503 37253 8541 37287
rect 8575 37253 8581 37287
rect 8391 37212 8581 37253
rect 8391 37178 8397 37212
rect 8431 37178 8469 37212
rect 8503 37178 8541 37212
rect 8575 37178 8581 37212
rect 8391 37137 8581 37178
rect 8391 37103 8397 37137
rect 8431 37103 8469 37137
rect 8503 37103 8541 37137
rect 8575 37103 8581 37137
rect 8391 36353 8581 37103
rect 8391 36290 8397 36353
rect 8575 36290 8581 36353
rect 8391 36238 8392 36290
rect 8580 36238 8581 36290
rect 8391 36226 8397 36238
rect 8575 36226 8581 36238
rect 8391 36174 8392 36226
rect 8580 36174 8581 36226
rect 8391 36162 8397 36174
rect 8575 36162 8581 36174
rect 8391 36110 8392 36162
rect 8580 36110 8581 36162
rect 8391 36098 8397 36110
rect 8575 36098 8581 36110
rect 8391 36046 8392 36098
rect 8580 36046 8581 36098
rect 8391 36034 8397 36046
rect 8575 36034 8581 36046
rect 8391 35982 8392 36034
rect 8580 35982 8581 36034
rect 8391 35970 8397 35982
rect 8575 35970 8581 35982
rect 8391 35918 8392 35970
rect 8580 35918 8581 35970
rect 8391 35906 8397 35918
rect 8575 35906 8581 35918
rect 8391 35854 8392 35906
rect 8580 35854 8581 35906
rect 8391 35842 8397 35854
rect 8575 35842 8581 35854
rect 8391 35790 8392 35842
rect 8580 35790 8581 35842
rect 8391 35778 8397 35790
rect 8575 35778 8581 35790
rect 8391 35726 8392 35778
rect 8580 35726 8581 35778
rect 8391 35714 8397 35726
rect 8575 35714 8581 35726
rect 8391 35662 8392 35714
rect 8580 35662 8581 35714
rect 8391 35650 8397 35662
rect 8575 35650 8581 35662
rect 8391 35598 8392 35650
rect 8580 35598 8581 35650
rect 8391 35586 8397 35598
rect 8575 35586 8581 35598
rect 8391 35534 8392 35586
rect 8580 35534 8581 35586
rect 8391 35522 8397 35534
rect 8575 35522 8581 35534
rect 8391 35470 8392 35522
rect 8580 35470 8581 35522
rect 8391 35458 8397 35470
rect 8575 35458 8581 35470
rect 8391 35406 8392 35458
rect 8580 35406 8581 35458
rect 8391 35394 8397 35406
rect 8575 35394 8581 35406
rect 8391 35342 8392 35394
rect 8580 35342 8581 35394
rect 8391 35329 8397 35342
rect 8575 35329 8581 35342
rect 8391 35277 8392 35329
rect 8580 35277 8581 35329
rect 8391 35264 8397 35277
rect 8575 35264 8581 35277
rect 8391 35212 8392 35264
rect 8580 35212 8581 35264
rect 8391 35199 8397 35212
rect 8575 35199 8581 35212
rect 8391 35147 8392 35199
rect 8580 35147 8581 35199
rect 8391 35134 8397 35147
rect 8575 35134 8581 35147
rect 8391 35082 8392 35134
rect 8580 35082 8581 35134
rect 8391 35069 8397 35082
rect 8575 35069 8581 35082
rect 8391 35017 8392 35069
rect 8580 35017 8581 35069
rect 8391 35004 8397 35017
rect 8575 35004 8581 35017
rect 8391 34952 8392 35004
rect 8580 34952 8581 35004
rect 8391 34939 8397 34952
rect 8575 34939 8581 34952
rect 8391 34887 8392 34939
rect 8580 34887 8581 34939
rect 8391 34874 8397 34887
rect 8575 34874 8581 34887
rect 8391 34822 8392 34874
rect 8580 34822 8581 34874
rect 8391 34809 8397 34822
rect 8575 34809 8581 34822
rect 8391 34757 8392 34809
rect 8580 34757 8581 34809
rect 8391 34744 8397 34757
rect 8575 34744 8581 34757
rect 8391 34692 8392 34744
rect 8580 34692 8581 34744
rect 8391 34679 8397 34692
rect 8575 34679 8581 34692
rect 8391 34627 8392 34679
rect 8580 34627 8581 34679
rect 8391 34614 8397 34627
rect 8575 34614 8581 34627
rect 8391 34562 8392 34614
rect 8580 34562 8581 34614
rect 8391 32503 8397 34562
rect 8575 32503 8581 34562
rect 8391 31753 8581 32503
rect 8391 31690 8397 31753
rect 8575 31690 8581 31753
rect 8391 31638 8392 31690
rect 8580 31638 8581 31690
rect 8391 31626 8397 31638
rect 8575 31626 8581 31638
rect 8391 31574 8392 31626
rect 8580 31574 8581 31626
rect 8391 31562 8397 31574
rect 8575 31562 8581 31574
rect 8391 31510 8392 31562
rect 8580 31510 8581 31562
rect 8391 31498 8397 31510
rect 8575 31498 8581 31510
rect 8391 31446 8392 31498
rect 8580 31446 8581 31498
rect 8391 31434 8397 31446
rect 8575 31434 8581 31446
rect 8391 31382 8392 31434
rect 8580 31382 8581 31434
rect 8391 31370 8397 31382
rect 8575 31370 8581 31382
rect 8391 31318 8392 31370
rect 8580 31318 8581 31370
rect 8391 31306 8397 31318
rect 8575 31306 8581 31318
rect 8391 31254 8392 31306
rect 8580 31254 8581 31306
rect 8391 31242 8397 31254
rect 8575 31242 8581 31254
rect 8391 31190 8392 31242
rect 8580 31190 8581 31242
rect 8391 31178 8397 31190
rect 8575 31178 8581 31190
rect 8391 31126 8392 31178
rect 8580 31126 8581 31178
rect 8391 31114 8397 31126
rect 8575 31114 8581 31126
rect 8391 31062 8392 31114
rect 8580 31062 8581 31114
rect 8391 31050 8397 31062
rect 8575 31050 8581 31062
rect 8391 30998 8392 31050
rect 8580 30998 8581 31050
rect 8391 30986 8397 30998
rect 8575 30986 8581 30998
rect 8391 30934 8392 30986
rect 8580 30934 8581 30986
rect 8391 30922 8397 30934
rect 8575 30922 8581 30934
rect 8391 30870 8392 30922
rect 8580 30870 8581 30922
rect 8391 30858 8397 30870
rect 8575 30858 8581 30870
rect 8391 30806 8392 30858
rect 8580 30806 8581 30858
rect 8391 30794 8397 30806
rect 8575 30794 8581 30806
rect 8391 30742 8392 30794
rect 8580 30742 8581 30794
rect 8391 30729 8397 30742
rect 8575 30729 8581 30742
rect 8391 30677 8392 30729
rect 8580 30677 8581 30729
rect 8391 30664 8397 30677
rect 8575 30664 8581 30677
rect 8391 30612 8392 30664
rect 8580 30612 8581 30664
rect 8391 30599 8397 30612
rect 8575 30599 8581 30612
rect 8391 30547 8392 30599
rect 8580 30547 8581 30599
rect 8391 30534 8397 30547
rect 8575 30534 8581 30547
rect 8391 30482 8392 30534
rect 8580 30482 8581 30534
rect 8391 30469 8397 30482
rect 8575 30469 8581 30482
rect 8391 30417 8392 30469
rect 8580 30417 8581 30469
rect 8391 30404 8397 30417
rect 8575 30404 8581 30417
rect 8391 30352 8392 30404
rect 8580 30352 8581 30404
rect 8391 30339 8397 30352
rect 8575 30339 8581 30352
rect 8391 30287 8392 30339
rect 8580 30287 8581 30339
rect 8391 30274 8397 30287
rect 8575 30274 8581 30287
rect 8391 30222 8392 30274
rect 8580 30222 8581 30274
rect 8391 30209 8397 30222
rect 8575 30209 8581 30222
rect 8391 30157 8392 30209
rect 8580 30157 8581 30209
rect 8391 30144 8397 30157
rect 8575 30144 8581 30157
rect 8391 30092 8392 30144
rect 8580 30092 8581 30144
rect 8391 30079 8397 30092
rect 8575 30079 8581 30092
rect 8391 30027 8392 30079
rect 8580 30027 8581 30079
rect 8391 30014 8397 30027
rect 8575 30014 8581 30027
rect 8391 29962 8392 30014
rect 8580 29962 8581 30014
rect 8391 27903 8397 29962
rect 8575 27903 8581 29962
rect 8391 27153 8581 27903
rect 8391 27090 8397 27153
rect 8575 27090 8581 27153
rect 8391 27038 8392 27090
rect 8580 27038 8581 27090
rect 8391 27026 8397 27038
rect 8575 27026 8581 27038
rect 8391 26974 8392 27026
rect 8580 26974 8581 27026
rect 8391 26962 8397 26974
rect 8575 26962 8581 26974
rect 8391 26910 8392 26962
rect 8580 26910 8581 26962
rect 8391 26898 8397 26910
rect 8575 26898 8581 26910
rect 8391 26846 8392 26898
rect 8580 26846 8581 26898
rect 8391 26834 8397 26846
rect 8575 26834 8581 26846
rect 8391 26782 8392 26834
rect 8580 26782 8581 26834
rect 8391 26770 8397 26782
rect 8575 26770 8581 26782
rect 8391 26718 8392 26770
rect 8580 26718 8581 26770
rect 8391 26706 8397 26718
rect 8575 26706 8581 26718
rect 8391 26654 8392 26706
rect 8580 26654 8581 26706
rect 8391 26642 8397 26654
rect 8575 26642 8581 26654
rect 8391 26590 8392 26642
rect 8580 26590 8581 26642
rect 8391 26578 8397 26590
rect 8575 26578 8581 26590
rect 8391 26526 8392 26578
rect 8580 26526 8581 26578
rect 8391 26514 8397 26526
rect 8575 26514 8581 26526
rect 8391 26462 8392 26514
rect 8580 26462 8581 26514
rect 8391 26450 8397 26462
rect 8575 26450 8581 26462
rect 8391 26398 8392 26450
rect 8580 26398 8581 26450
rect 8391 26386 8397 26398
rect 8575 26386 8581 26398
rect 8391 26334 8392 26386
rect 8580 26334 8581 26386
rect 8391 26322 8397 26334
rect 8575 26322 8581 26334
rect 8391 26270 8392 26322
rect 8580 26270 8581 26322
rect 8391 26258 8397 26270
rect 8575 26258 8581 26270
rect 8391 26206 8392 26258
rect 8580 26206 8581 26258
rect 8391 26194 8397 26206
rect 8575 26194 8581 26206
rect 8391 26142 8392 26194
rect 8580 26142 8581 26194
rect 8391 26129 8397 26142
rect 8575 26129 8581 26142
rect 8391 26077 8392 26129
rect 8580 26077 8581 26129
rect 8391 26064 8397 26077
rect 8575 26064 8581 26077
rect 8391 26012 8392 26064
rect 8580 26012 8581 26064
rect 8391 25999 8397 26012
rect 8575 25999 8581 26012
rect 8391 25947 8392 25999
rect 8580 25947 8581 25999
rect 8391 25934 8397 25947
rect 8575 25934 8581 25947
rect 8391 25882 8392 25934
rect 8580 25882 8581 25934
rect 8391 25869 8397 25882
rect 8575 25869 8581 25882
rect 8391 25817 8392 25869
rect 8580 25817 8581 25869
rect 8391 25804 8397 25817
rect 8575 25804 8581 25817
rect 8391 25752 8392 25804
rect 8580 25752 8581 25804
rect 8391 25739 8397 25752
rect 8575 25739 8581 25752
rect 8391 25687 8392 25739
rect 8580 25687 8581 25739
rect 8391 25674 8397 25687
rect 8575 25674 8581 25687
rect 8391 25622 8392 25674
rect 8580 25622 8581 25674
rect 8391 25609 8397 25622
rect 8575 25609 8581 25622
rect 8391 25557 8392 25609
rect 8580 25557 8581 25609
rect 8391 25544 8397 25557
rect 8575 25544 8581 25557
rect 8391 25492 8392 25544
rect 8580 25492 8581 25544
rect 8391 25479 8397 25492
rect 8575 25479 8581 25492
rect 8391 25427 8392 25479
rect 8580 25427 8581 25479
rect 8391 25414 8397 25427
rect 8575 25414 8581 25427
rect 8391 25362 8392 25414
rect 8580 25362 8581 25414
rect 8391 23303 8397 25362
rect 8575 23303 8581 25362
rect 8391 22562 8581 23303
rect 8391 22490 8397 22562
rect 8575 22490 8581 22562
rect 8391 22438 8392 22490
rect 8580 22438 8581 22490
rect 8391 22426 8397 22438
rect 8575 22426 8581 22438
rect 8391 22374 8392 22426
rect 8580 22374 8581 22426
rect 8391 22362 8397 22374
rect 8575 22362 8581 22374
rect 8391 22310 8392 22362
rect 8580 22310 8581 22362
rect 8391 22298 8397 22310
rect 8575 22298 8581 22310
rect 8391 22246 8392 22298
rect 8580 22246 8581 22298
rect 8391 22234 8397 22246
rect 8575 22234 8581 22246
rect 8391 22182 8392 22234
rect 8580 22182 8581 22234
rect 8391 22170 8397 22182
rect 8575 22170 8581 22182
rect 8391 22118 8392 22170
rect 8580 22118 8581 22170
rect 8391 22106 8397 22118
rect 8575 22106 8581 22118
rect 8391 22054 8392 22106
rect 8580 22054 8581 22106
rect 8391 22042 8397 22054
rect 8575 22042 8581 22054
rect 8391 21990 8392 22042
rect 8580 21990 8581 22042
rect 8391 21978 8397 21990
rect 8575 21978 8581 21990
rect 8391 21926 8392 21978
rect 8580 21926 8581 21978
rect 8391 21914 8397 21926
rect 8575 21914 8581 21926
rect 8391 21862 8392 21914
rect 8580 21862 8581 21914
rect 8391 21850 8397 21862
rect 8575 21850 8581 21862
rect 8391 21798 8392 21850
rect 8580 21798 8581 21850
rect 8391 21786 8397 21798
rect 8575 21786 8581 21798
rect 8391 21734 8392 21786
rect 8580 21734 8581 21786
rect 8391 21722 8397 21734
rect 8575 21722 8581 21734
rect 8391 21670 8392 21722
rect 8580 21670 8581 21722
rect 8391 21658 8397 21670
rect 8575 21658 8581 21670
rect 8391 21606 8392 21658
rect 8580 21606 8581 21658
rect 8391 21594 8397 21606
rect 8575 21594 8581 21606
rect 8391 21542 8392 21594
rect 8580 21542 8581 21594
rect 8391 21529 8397 21542
rect 8575 21529 8581 21542
rect 8391 21477 8392 21529
rect 8580 21477 8581 21529
rect 8391 21464 8397 21477
rect 8575 21464 8581 21477
rect 8391 21412 8392 21464
rect 8580 21412 8581 21464
rect 8391 21399 8397 21412
rect 8575 21399 8581 21412
rect 8391 21347 8392 21399
rect 8580 21347 8581 21399
rect 8391 21334 8397 21347
rect 8575 21334 8581 21347
rect 8391 21282 8392 21334
rect 8580 21282 8581 21334
rect 8391 21269 8397 21282
rect 8575 21269 8581 21282
rect 8391 21217 8392 21269
rect 8580 21217 8581 21269
rect 8391 21204 8397 21217
rect 8575 21204 8581 21217
rect 8391 21152 8392 21204
rect 8580 21152 8581 21204
rect 8391 21139 8397 21152
rect 8575 21139 8581 21152
rect 8391 21087 8392 21139
rect 8580 21087 8581 21139
rect 8391 21074 8397 21087
rect 8575 21074 8581 21087
rect 8391 21022 8392 21074
rect 8580 21022 8581 21074
rect 8391 21009 8397 21022
rect 8575 21009 8581 21022
rect 8391 20957 8392 21009
rect 8580 20957 8581 21009
rect 8391 20944 8397 20957
rect 8575 20944 8581 20957
rect 8391 20892 8392 20944
rect 8580 20892 8581 20944
rect 8391 20879 8397 20892
rect 8575 20879 8581 20892
rect 8391 20827 8392 20879
rect 8580 20827 8581 20879
rect 8391 20814 8397 20827
rect 8575 20814 8581 20827
rect 8391 20762 8392 20814
rect 8580 20762 8581 20814
rect 8391 19360 8397 20762
rect 8575 19360 8581 20762
rect 8391 19321 8581 19360
rect 8391 19287 8397 19321
rect 8431 19287 8469 19321
rect 8503 19287 8541 19321
rect 8575 19287 8581 19321
rect 8391 19248 8581 19287
rect 8391 19214 8397 19248
rect 8431 19214 8469 19248
rect 8503 19214 8541 19248
rect 8575 19214 8581 19248
rect 8391 19175 8581 19214
rect 8391 19141 8397 19175
rect 8431 19141 8469 19175
rect 8503 19141 8541 19175
rect 8575 19141 8581 19175
rect 8391 19102 8581 19141
rect 8391 19068 8397 19102
rect 8431 19068 8469 19102
rect 8503 19068 8541 19102
rect 8575 19068 8581 19102
rect 8391 19029 8581 19068
rect 8391 18995 8397 19029
rect 8431 18995 8469 19029
rect 8503 18995 8541 19029
rect 8575 18995 8581 19029
rect 8391 18956 8581 18995
rect 8391 18922 8397 18956
rect 8431 18922 8469 18956
rect 8503 18922 8541 18956
rect 8575 18922 8581 18956
rect 8391 18883 8581 18922
rect 8391 18849 8397 18883
rect 8431 18849 8469 18883
rect 8503 18849 8541 18883
rect 8575 18849 8581 18883
rect 8391 18810 8581 18849
rect 8391 18776 8397 18810
rect 8431 18776 8469 18810
rect 8503 18776 8541 18810
rect 8575 18776 8581 18810
rect 8391 18737 8581 18776
rect 8391 18703 8397 18737
rect 8431 18703 8469 18737
rect 8503 18703 8541 18737
rect 8575 18703 8581 18737
rect 8391 17953 8581 18703
rect 8391 17890 8397 17953
rect 8575 17890 8581 17953
rect 8391 17838 8392 17890
rect 8580 17838 8581 17890
rect 8391 17826 8397 17838
rect 8575 17826 8581 17838
rect 8391 17774 8392 17826
rect 8580 17774 8581 17826
rect 8391 17762 8397 17774
rect 8575 17762 8581 17774
rect 8391 17710 8392 17762
rect 8580 17710 8581 17762
rect 8391 17698 8397 17710
rect 8575 17698 8581 17710
rect 8391 17646 8392 17698
rect 8580 17646 8581 17698
rect 8391 17634 8397 17646
rect 8575 17634 8581 17646
rect 8391 17582 8392 17634
rect 8580 17582 8581 17634
rect 8391 17570 8397 17582
rect 8575 17570 8581 17582
rect 8391 17518 8392 17570
rect 8580 17518 8581 17570
rect 8391 17506 8397 17518
rect 8575 17506 8581 17518
rect 8391 17454 8392 17506
rect 8580 17454 8581 17506
rect 8391 17442 8397 17454
rect 8575 17442 8581 17454
rect 8391 17390 8392 17442
rect 8580 17390 8581 17442
rect 8391 17378 8397 17390
rect 8575 17378 8581 17390
rect 8391 17326 8392 17378
rect 8580 17326 8581 17378
rect 8391 17314 8397 17326
rect 8575 17314 8581 17326
rect 8391 17262 8392 17314
rect 8580 17262 8581 17314
rect 8391 17250 8397 17262
rect 8575 17250 8581 17262
rect 8391 17198 8392 17250
rect 8580 17198 8581 17250
rect 8391 17186 8397 17198
rect 8575 17186 8581 17198
rect 8391 17134 8392 17186
rect 8580 17134 8581 17186
rect 8391 17122 8397 17134
rect 8575 17122 8581 17134
rect 8391 17070 8392 17122
rect 8580 17070 8581 17122
rect 8391 17058 8397 17070
rect 8575 17058 8581 17070
rect 8391 17006 8392 17058
rect 8580 17006 8581 17058
rect 8391 16994 8397 17006
rect 8575 16994 8581 17006
rect 8391 16942 8392 16994
rect 8580 16942 8581 16994
rect 8391 16929 8397 16942
rect 8575 16929 8581 16942
rect 8391 16877 8392 16929
rect 8580 16877 8581 16929
rect 8391 16864 8397 16877
rect 8575 16864 8581 16877
rect 8391 16812 8392 16864
rect 8580 16812 8581 16864
rect 8391 16799 8397 16812
rect 8575 16799 8581 16812
rect 8391 16747 8392 16799
rect 8580 16747 8581 16799
rect 8391 16734 8397 16747
rect 8575 16734 8581 16747
rect 8391 16682 8392 16734
rect 8580 16682 8581 16734
rect 8391 16669 8397 16682
rect 8575 16669 8581 16682
rect 8391 16617 8392 16669
rect 8580 16617 8581 16669
rect 8391 16604 8397 16617
rect 8575 16604 8581 16617
rect 8391 16552 8392 16604
rect 8580 16552 8581 16604
rect 8391 16539 8397 16552
rect 8575 16539 8581 16552
rect 8391 16487 8392 16539
rect 8580 16487 8581 16539
rect 8391 16474 8397 16487
rect 8575 16474 8581 16487
rect 8391 16422 8392 16474
rect 8580 16422 8581 16474
rect 8391 16409 8397 16422
rect 8575 16409 8581 16422
rect 8391 16357 8392 16409
rect 8580 16357 8581 16409
rect 8391 16344 8397 16357
rect 8575 16344 8581 16357
rect 8391 16292 8392 16344
rect 8580 16292 8581 16344
rect 8391 16279 8397 16292
rect 8575 16279 8581 16292
rect 8391 16227 8392 16279
rect 8580 16227 8581 16279
rect 8391 16214 8397 16227
rect 8575 16214 8581 16227
rect 8391 16162 8392 16214
rect 8580 16162 8581 16214
rect 8391 14103 8397 16162
rect 8575 14103 8581 16162
rect 8391 13362 8581 14103
rect 8391 13290 8397 13362
rect 8575 13290 8581 13362
rect 8391 13238 8392 13290
rect 8580 13238 8581 13290
rect 8391 13226 8397 13238
rect 8575 13226 8581 13238
rect 8391 13174 8392 13226
rect 8580 13174 8581 13226
rect 8391 13162 8397 13174
rect 8575 13162 8581 13174
rect 8391 13110 8392 13162
rect 8580 13110 8581 13162
rect 8391 13098 8397 13110
rect 8575 13098 8581 13110
rect 8391 13046 8392 13098
rect 8580 13046 8581 13098
rect 8391 13034 8397 13046
rect 8575 13034 8581 13046
rect 8391 12982 8392 13034
rect 8580 12982 8581 13034
rect 8391 12970 8397 12982
rect 8575 12970 8581 12982
rect 8391 12918 8392 12970
rect 8580 12918 8581 12970
rect 8391 12906 8397 12918
rect 8575 12906 8581 12918
rect 8391 12854 8392 12906
rect 8580 12854 8581 12906
rect 8391 12842 8397 12854
rect 8575 12842 8581 12854
rect 8391 12790 8392 12842
rect 8580 12790 8581 12842
rect 8391 12778 8397 12790
rect 8575 12778 8581 12790
rect 8391 12726 8392 12778
rect 8580 12726 8581 12778
rect 8391 12714 8397 12726
rect 8575 12714 8581 12726
rect 8391 12662 8392 12714
rect 8580 12662 8581 12714
rect 8391 12650 8397 12662
rect 8575 12650 8581 12662
rect 8391 12598 8392 12650
rect 8580 12598 8581 12650
rect 8391 12586 8397 12598
rect 8575 12586 8581 12598
rect 8391 12534 8392 12586
rect 8580 12534 8581 12586
rect 8391 12522 8397 12534
rect 8575 12522 8581 12534
rect 8391 12470 8392 12522
rect 8580 12470 8581 12522
rect 8391 12458 8397 12470
rect 8575 12458 8581 12470
rect 8391 12406 8392 12458
rect 8580 12406 8581 12458
rect 8391 12394 8397 12406
rect 8575 12394 8581 12406
rect 8391 12342 8392 12394
rect 8580 12342 8581 12394
rect 8391 12329 8397 12342
rect 8575 12329 8581 12342
rect 8391 12277 8392 12329
rect 8580 12277 8581 12329
rect 8391 12264 8397 12277
rect 8575 12264 8581 12277
rect 8391 12212 8392 12264
rect 8580 12212 8581 12264
rect 8391 12199 8397 12212
rect 8575 12199 8581 12212
rect 8391 12147 8392 12199
rect 8580 12147 8581 12199
rect 8391 12134 8397 12147
rect 8575 12134 8581 12147
rect 8391 12082 8392 12134
rect 8580 12082 8581 12134
rect 8391 12069 8397 12082
rect 8575 12069 8581 12082
rect 8391 12017 8392 12069
rect 8580 12017 8581 12069
rect 8391 12004 8397 12017
rect 8575 12004 8581 12017
rect 8391 11952 8392 12004
rect 8580 11952 8581 12004
rect 8391 11939 8397 11952
rect 8575 11939 8581 11952
rect 8391 11887 8392 11939
rect 8580 11887 8581 11939
rect 8391 11874 8397 11887
rect 8575 11874 8581 11887
rect 8391 11822 8392 11874
rect 8580 11822 8581 11874
rect 8391 11809 8397 11822
rect 8575 11809 8581 11822
rect 8391 11757 8392 11809
rect 8580 11757 8581 11809
rect 8391 11744 8397 11757
rect 8575 11744 8581 11757
rect 8391 11692 8392 11744
rect 8580 11692 8581 11744
rect 8391 11679 8397 11692
rect 8575 11679 8581 11692
rect 8391 11627 8392 11679
rect 8580 11627 8581 11679
rect 8391 11614 8397 11627
rect 8575 11614 8581 11627
rect 8391 11562 8392 11614
rect 8580 11562 8581 11614
rect 8391 10160 8397 11562
rect 8575 10160 8581 11562
rect 8391 10121 8581 10160
rect 8391 10087 8397 10121
rect 8431 10087 8469 10121
rect 8503 10087 8541 10121
rect 8575 10087 8581 10121
rect 8391 10048 8581 10087
rect 8391 10014 8397 10048
rect 8431 10014 8469 10048
rect 8503 10014 8541 10048
rect 8575 10014 8581 10048
rect 8391 9975 8581 10014
rect 8391 9941 8397 9975
rect 8431 9941 8469 9975
rect 8503 9941 8541 9975
rect 8575 9941 8581 9975
rect 8391 9902 8581 9941
rect 8391 9868 8397 9902
rect 8431 9868 8469 9902
rect 8503 9868 8541 9902
rect 8575 9868 8581 9902
rect 8391 9829 8581 9868
rect 8391 9795 8397 9829
rect 8431 9795 8469 9829
rect 8503 9795 8541 9829
rect 8575 9795 8581 9829
rect 8391 9756 8581 9795
rect 8391 9722 8397 9756
rect 8431 9722 8469 9756
rect 8503 9722 8541 9756
rect 8575 9722 8581 9756
rect 8391 9683 8581 9722
rect 8391 9649 8397 9683
rect 8431 9649 8469 9683
rect 8503 9649 8541 9683
rect 8575 9649 8581 9683
rect 8391 9610 8581 9649
rect 8391 9576 8397 9610
rect 8431 9576 8469 9610
rect 8503 9576 8541 9610
rect 8575 9576 8581 9610
rect 8391 9537 8581 9576
rect 8391 9503 8397 9537
rect 8431 9503 8469 9537
rect 8503 9503 8541 9537
rect 8575 9503 8581 9537
rect 8391 9491 8581 9503
rect 8881 37997 9011 38003
rect 8933 37945 8959 37997
rect 8881 37929 9011 37945
rect 8933 37877 8959 37929
rect 8881 37861 9011 37877
rect 8933 37809 8959 37861
rect 8881 37793 9011 37809
rect 8933 37741 8959 37793
rect 8881 37725 9011 37741
rect 8933 37673 8959 37725
rect 8881 37657 9011 37673
rect 8933 37605 8959 37657
rect 8881 37589 9011 37605
rect 8933 37537 8959 37589
rect 8881 37521 9011 37537
rect 8933 37469 8959 37521
rect 8881 37453 9011 37469
rect 8933 37401 8959 37453
rect 8881 37385 9011 37401
rect 8933 37333 8959 37385
rect 8881 37318 9011 37333
rect 8933 37266 8959 37318
rect 8881 37251 9011 37266
rect 8933 37199 8959 37251
rect 8881 37184 9011 37199
rect 8933 37132 8959 37184
rect 8881 37117 9011 37132
rect 8933 37065 8959 37117
rect 8881 34225 9011 37065
rect 8933 34173 8959 34225
rect 8881 34161 9011 34173
rect 8933 34109 8959 34161
rect 8881 34097 9011 34109
rect 8933 34045 8959 34097
rect 8881 34033 9011 34045
rect 8933 33981 8959 34033
rect 8881 33969 9011 33981
rect 8933 33917 8959 33969
rect 8881 33905 9011 33917
rect 8933 33853 8959 33905
rect 8881 33841 9011 33853
rect 8933 33789 8959 33841
rect 8881 33777 9011 33789
rect 8933 33725 8959 33777
rect 8881 33713 9011 33725
rect 8933 33661 8959 33713
rect 8881 33649 9011 33661
rect 8933 33597 8959 33649
rect 8881 33585 9011 33597
rect 8933 33533 8959 33585
rect 8881 33521 9011 33533
rect 8933 33469 8959 33521
rect 8881 33457 9011 33469
rect 8933 33405 8959 33457
rect 8881 33393 9011 33405
rect 8933 33341 8959 33393
rect 8881 33329 9011 33341
rect 8933 33277 8959 33329
rect 8881 33264 9011 33277
rect 8933 33212 8959 33264
rect 8881 33199 9011 33212
rect 8933 33147 8959 33199
rect 8881 33134 9011 33147
rect 8933 33082 8959 33134
rect 8881 33069 9011 33082
rect 8933 33017 8959 33069
rect 8881 33004 9011 33017
rect 8933 32952 8959 33004
rect 8881 32939 9011 32952
rect 8933 32887 8959 32939
rect 8881 32874 9011 32887
rect 8933 32822 8959 32874
rect 8881 32809 9011 32822
rect 8933 32757 8959 32809
rect 8881 32744 9011 32757
rect 8933 32692 8959 32744
rect 8881 32679 9011 32692
rect 8933 32627 8959 32679
rect 8881 32614 9011 32627
rect 8933 32562 8959 32614
rect 8881 32549 9011 32562
rect 8933 32497 8959 32549
rect 8881 29625 9011 32497
rect 8933 29573 8959 29625
rect 8881 29561 9011 29573
rect 8933 29509 8959 29561
rect 8881 29497 9011 29509
rect 8933 29445 8959 29497
rect 8881 29433 9011 29445
rect 8933 29381 8959 29433
rect 8881 29369 9011 29381
rect 8933 29317 8959 29369
rect 8881 29305 9011 29317
rect 8933 29253 8959 29305
rect 8881 29241 9011 29253
rect 8933 29189 8959 29241
rect 8881 29177 9011 29189
rect 8933 29125 8959 29177
rect 8881 29113 9011 29125
rect 8933 29061 8959 29113
rect 8881 29049 9011 29061
rect 8933 28997 8959 29049
rect 8881 28985 9011 28997
rect 8933 28933 8959 28985
rect 8881 28921 9011 28933
rect 8933 28869 8959 28921
rect 8881 28857 9011 28869
rect 8933 28805 8959 28857
rect 8881 28793 9011 28805
rect 8933 28741 8959 28793
rect 8881 28729 9011 28741
rect 8933 28677 8959 28729
rect 8881 28664 9011 28677
rect 8933 28612 8959 28664
rect 8881 28599 9011 28612
rect 8933 28547 8959 28599
rect 8881 28534 9011 28547
rect 8933 28482 8959 28534
rect 8881 28469 9011 28482
rect 8933 28417 8959 28469
rect 8881 28404 9011 28417
rect 8933 28352 8959 28404
rect 8881 28339 9011 28352
rect 8933 28287 8959 28339
rect 8881 28274 9011 28287
rect 8933 28222 8959 28274
rect 8881 28209 9011 28222
rect 8933 28157 8959 28209
rect 8881 28144 9011 28157
rect 8933 28092 8959 28144
rect 8881 28079 9011 28092
rect 8933 28027 8959 28079
rect 8881 28014 9011 28027
rect 8933 27962 8959 28014
rect 8881 27949 9011 27962
rect 8933 27897 8959 27949
rect 8881 25025 9011 27897
rect 8933 24973 8959 25025
rect 8881 24961 9011 24973
rect 8933 24909 8959 24961
rect 8881 24897 9011 24909
rect 8933 24845 8959 24897
rect 8881 24833 9011 24845
rect 8933 24781 8959 24833
rect 8881 24769 9011 24781
rect 8933 24717 8959 24769
rect 8881 24705 9011 24717
rect 8933 24653 8959 24705
rect 8881 24641 9011 24653
rect 8933 24589 8959 24641
rect 8881 24577 9011 24589
rect 8933 24525 8959 24577
rect 8881 24513 9011 24525
rect 8933 24461 8959 24513
rect 8881 24449 9011 24461
rect 8933 24397 8959 24449
rect 8881 24385 9011 24397
rect 8933 24333 8959 24385
rect 8881 24321 9011 24333
rect 8933 24269 8959 24321
rect 8881 24257 9011 24269
rect 8933 24205 8959 24257
rect 8881 24193 9011 24205
rect 8933 24141 8959 24193
rect 8881 24129 9011 24141
rect 8933 24077 8959 24129
rect 8881 24064 9011 24077
rect 8933 24012 8959 24064
rect 8881 23999 9011 24012
rect 8933 23947 8959 23999
rect 8881 23934 9011 23947
rect 8933 23882 8959 23934
rect 8881 23869 9011 23882
rect 8933 23817 8959 23869
rect 8881 23804 9011 23817
rect 8933 23752 8959 23804
rect 8881 23739 9011 23752
rect 8933 23687 8959 23739
rect 8881 23674 9011 23687
rect 8933 23622 8959 23674
rect 8881 23609 9011 23622
rect 8933 23557 8959 23609
rect 8881 23544 9011 23557
rect 8933 23492 8959 23544
rect 8881 23479 9011 23492
rect 8933 23427 8959 23479
rect 8881 23414 9011 23427
rect 8933 23362 8959 23414
rect 8881 23349 9011 23362
rect 8933 23297 8959 23349
rect 8881 20425 9011 23297
rect 8933 20373 8959 20425
rect 8881 20361 9011 20373
rect 8933 20309 8959 20361
rect 8881 20297 9011 20309
rect 8933 20245 8959 20297
rect 8881 20233 9011 20245
rect 8933 20181 8959 20233
rect 8881 20169 9011 20181
rect 8933 20117 8959 20169
rect 8881 20105 9011 20117
rect 8933 20053 8959 20105
rect 8881 20041 9011 20053
rect 8933 19989 8959 20041
rect 8881 19977 9011 19989
rect 8933 19925 8959 19977
rect 8881 19913 9011 19925
rect 8933 19861 8959 19913
rect 8881 19849 9011 19861
rect 8933 19797 8959 19849
rect 8881 19785 9011 19797
rect 8933 19733 8959 19785
rect 8881 19721 9011 19733
rect 8933 19669 8959 19721
rect 8881 19657 9011 19669
rect 8933 19605 8959 19657
rect 8881 19593 9011 19605
rect 8933 19541 8959 19593
rect 8881 19529 9011 19541
rect 8933 19477 8959 19529
rect 8881 19464 9011 19477
rect 8933 19412 8959 19464
rect 8881 19399 9011 19412
rect 8933 19347 8959 19399
rect 8881 19334 9011 19347
rect 8933 19282 8959 19334
rect 8881 19269 9011 19282
rect 8933 19217 8959 19269
rect 8881 19204 9011 19217
rect 8933 19152 8959 19204
rect 8881 19139 9011 19152
rect 8933 19087 8959 19139
rect 8881 19074 9011 19087
rect 8933 19022 8959 19074
rect 8881 19009 9011 19022
rect 8933 18957 8959 19009
rect 8881 18944 9011 18957
rect 8933 18892 8959 18944
rect 8881 18879 9011 18892
rect 8933 18827 8959 18879
rect 8881 18814 9011 18827
rect 8933 18762 8959 18814
rect 8881 18749 9011 18762
rect 8933 18697 8959 18749
rect 8881 15825 9011 18697
rect 8933 15773 8959 15825
rect 8881 15761 9011 15773
rect 8933 15709 8959 15761
rect 8881 15697 9011 15709
rect 8933 15645 8959 15697
rect 8881 15633 9011 15645
rect 8933 15581 8959 15633
rect 8881 15569 9011 15581
rect 8933 15517 8959 15569
rect 8881 15505 9011 15517
rect 8933 15453 8959 15505
rect 8881 15441 9011 15453
rect 8933 15389 8959 15441
rect 8881 15377 9011 15389
rect 8933 15325 8959 15377
rect 8881 15313 9011 15325
rect 8933 15261 8959 15313
rect 8881 15249 9011 15261
rect 8933 15197 8959 15249
rect 8881 15185 9011 15197
rect 8933 15133 8959 15185
rect 8881 15121 9011 15133
rect 8933 15069 8959 15121
rect 8881 15057 9011 15069
rect 8933 15005 8959 15057
rect 8881 14993 9011 15005
rect 8933 14941 8959 14993
rect 8881 14929 9011 14941
rect 8933 14877 8959 14929
rect 8881 14864 9011 14877
rect 8933 14812 8959 14864
rect 8881 14799 9011 14812
rect 8933 14747 8959 14799
rect 8881 14734 9011 14747
rect 8933 14682 8959 14734
rect 8881 14669 9011 14682
rect 8933 14617 8959 14669
rect 8881 14604 9011 14617
rect 8933 14552 8959 14604
rect 8881 14539 9011 14552
rect 8933 14487 8959 14539
rect 8881 14474 9011 14487
rect 8933 14422 8959 14474
rect 8881 14409 9011 14422
rect 8933 14357 8959 14409
rect 8881 14344 9011 14357
rect 8933 14292 8959 14344
rect 8881 14279 9011 14292
rect 8933 14227 8959 14279
rect 8881 14214 9011 14227
rect 8933 14162 8959 14214
rect 8881 14149 9011 14162
rect 8933 14097 8959 14149
rect 8881 11225 9011 14097
rect 8933 11173 8959 11225
rect 8881 11161 9011 11173
rect 8933 11109 8959 11161
rect 8881 11097 9011 11109
rect 8933 11045 8959 11097
rect 8881 11033 9011 11045
rect 8933 10981 8959 11033
rect 8881 10969 9011 10981
rect 8933 10917 8959 10969
rect 8881 10905 9011 10917
rect 8933 10853 8959 10905
rect 8881 10841 9011 10853
rect 8933 10789 8959 10841
rect 8881 10777 9011 10789
rect 8933 10725 8959 10777
rect 8881 10713 9011 10725
rect 8933 10661 8959 10713
rect 8881 10649 9011 10661
rect 8933 10597 8959 10649
rect 8881 10585 9011 10597
rect 8933 10533 8959 10585
rect 8881 10521 9011 10533
rect 8933 10469 8959 10521
rect 8881 10457 9011 10469
rect 8933 10405 8959 10457
rect 8881 10393 9011 10405
rect 8933 10341 8959 10393
rect 8881 10329 9011 10341
rect 8933 10277 8959 10329
rect 8881 10264 9011 10277
rect 8933 10212 8959 10264
rect 8881 10199 9011 10212
rect 8933 10147 8959 10199
rect 8881 10134 9011 10147
rect 8933 10082 8959 10134
rect 8881 10069 9011 10082
rect 8933 10017 8959 10069
rect 8881 10004 9011 10017
rect 8933 9952 8959 10004
rect 8881 9939 9011 9952
rect 8933 9887 8959 9939
rect 8881 9874 9011 9887
rect 8933 9822 8959 9874
rect 8881 9809 9011 9822
rect 8933 9757 8959 9809
rect 8881 9744 9011 9757
rect 8933 9692 8959 9744
rect 8881 9679 9011 9692
rect 8933 9627 8959 9679
rect 8881 9614 9011 9627
rect 8933 9562 8959 9614
rect 8881 9549 9011 9562
rect 8933 9497 8959 9549
rect 8881 9491 9011 9497
rect 9311 37962 9501 38003
rect 9311 37928 9317 37962
rect 9351 37928 9389 37962
rect 9423 37928 9461 37962
rect 9495 37928 9501 37962
rect 9311 37887 9501 37928
rect 9311 37853 9317 37887
rect 9351 37853 9389 37887
rect 9423 37853 9461 37887
rect 9495 37853 9501 37887
rect 9311 37812 9501 37853
rect 9311 37778 9317 37812
rect 9351 37778 9389 37812
rect 9423 37778 9461 37812
rect 9495 37778 9501 37812
rect 9311 37737 9501 37778
rect 9311 37703 9317 37737
rect 9351 37703 9389 37737
rect 9423 37703 9461 37737
rect 9495 37703 9501 37737
rect 9311 37662 9501 37703
rect 9311 37628 9317 37662
rect 9351 37628 9389 37662
rect 9423 37628 9461 37662
rect 9495 37628 9501 37662
rect 9311 37587 9501 37628
rect 9311 37553 9317 37587
rect 9351 37553 9389 37587
rect 9423 37553 9461 37587
rect 9495 37553 9501 37587
rect 9311 37512 9501 37553
rect 9311 37478 9317 37512
rect 9351 37478 9389 37512
rect 9423 37478 9461 37512
rect 9495 37478 9501 37512
rect 9311 37437 9501 37478
rect 9311 37403 9317 37437
rect 9351 37403 9389 37437
rect 9423 37403 9461 37437
rect 9495 37403 9501 37437
rect 9311 37362 9501 37403
rect 9311 37328 9317 37362
rect 9351 37328 9389 37362
rect 9423 37328 9461 37362
rect 9495 37328 9501 37362
rect 9311 37287 9501 37328
rect 9311 37253 9317 37287
rect 9351 37253 9389 37287
rect 9423 37253 9461 37287
rect 9495 37253 9501 37287
rect 9311 37212 9501 37253
rect 9311 37178 9317 37212
rect 9351 37178 9389 37212
rect 9423 37178 9461 37212
rect 9495 37178 9501 37212
rect 9311 37137 9501 37178
rect 9311 37103 9317 37137
rect 9351 37103 9389 37137
rect 9423 37103 9461 37137
rect 9495 37103 9501 37137
rect 9311 36353 9501 37103
rect 9311 36290 9317 36353
rect 9495 36290 9501 36353
rect 9311 36238 9312 36290
rect 9500 36238 9501 36290
rect 9311 36226 9317 36238
rect 9495 36226 9501 36238
rect 9311 36174 9312 36226
rect 9500 36174 9501 36226
rect 9311 36162 9317 36174
rect 9495 36162 9501 36174
rect 9311 36110 9312 36162
rect 9500 36110 9501 36162
rect 9311 36098 9317 36110
rect 9495 36098 9501 36110
rect 9311 36046 9312 36098
rect 9500 36046 9501 36098
rect 9311 36034 9317 36046
rect 9495 36034 9501 36046
rect 9311 35982 9312 36034
rect 9500 35982 9501 36034
rect 9311 35970 9317 35982
rect 9495 35970 9501 35982
rect 9311 35918 9312 35970
rect 9500 35918 9501 35970
rect 9311 35906 9317 35918
rect 9495 35906 9501 35918
rect 9311 35854 9312 35906
rect 9500 35854 9501 35906
rect 9311 35842 9317 35854
rect 9495 35842 9501 35854
rect 9311 35790 9312 35842
rect 9500 35790 9501 35842
rect 9311 35778 9317 35790
rect 9495 35778 9501 35790
rect 9311 35726 9312 35778
rect 9500 35726 9501 35778
rect 9311 35714 9317 35726
rect 9495 35714 9501 35726
rect 9311 35662 9312 35714
rect 9500 35662 9501 35714
rect 9311 35650 9317 35662
rect 9495 35650 9501 35662
rect 9311 35598 9312 35650
rect 9500 35598 9501 35650
rect 9311 35586 9317 35598
rect 9495 35586 9501 35598
rect 9311 35534 9312 35586
rect 9500 35534 9501 35586
rect 9311 35522 9317 35534
rect 9495 35522 9501 35534
rect 9311 35470 9312 35522
rect 9500 35470 9501 35522
rect 9311 35458 9317 35470
rect 9495 35458 9501 35470
rect 9311 35406 9312 35458
rect 9500 35406 9501 35458
rect 9311 35394 9317 35406
rect 9495 35394 9501 35406
rect 9311 35342 9312 35394
rect 9500 35342 9501 35394
rect 9311 35329 9317 35342
rect 9495 35329 9501 35342
rect 9311 35277 9312 35329
rect 9500 35277 9501 35329
rect 9311 35264 9317 35277
rect 9495 35264 9501 35277
rect 9311 35212 9312 35264
rect 9500 35212 9501 35264
rect 9311 35199 9317 35212
rect 9495 35199 9501 35212
rect 9311 35147 9312 35199
rect 9500 35147 9501 35199
rect 9311 35134 9317 35147
rect 9495 35134 9501 35147
rect 9311 35082 9312 35134
rect 9500 35082 9501 35134
rect 9311 35069 9317 35082
rect 9495 35069 9501 35082
rect 9311 35017 9312 35069
rect 9500 35017 9501 35069
rect 9311 35004 9317 35017
rect 9495 35004 9501 35017
rect 9311 34952 9312 35004
rect 9500 34952 9501 35004
rect 9311 34939 9317 34952
rect 9495 34939 9501 34952
rect 9311 34887 9312 34939
rect 9500 34887 9501 34939
rect 9311 34874 9317 34887
rect 9495 34874 9501 34887
rect 9311 34822 9312 34874
rect 9500 34822 9501 34874
rect 9311 34809 9317 34822
rect 9495 34809 9501 34822
rect 9311 34757 9312 34809
rect 9500 34757 9501 34809
rect 9311 34744 9317 34757
rect 9495 34744 9501 34757
rect 9311 34692 9312 34744
rect 9500 34692 9501 34744
rect 9311 34679 9317 34692
rect 9495 34679 9501 34692
rect 9311 34627 9312 34679
rect 9500 34627 9501 34679
rect 9311 34614 9317 34627
rect 9495 34614 9501 34627
rect 9311 34562 9312 34614
rect 9500 34562 9501 34614
rect 9311 32503 9317 34562
rect 9495 32503 9501 34562
rect 9311 31753 9501 32503
rect 9311 31690 9317 31753
rect 9495 31690 9501 31753
rect 9311 31638 9312 31690
rect 9500 31638 9501 31690
rect 9311 31626 9317 31638
rect 9495 31626 9501 31638
rect 9311 31574 9312 31626
rect 9500 31574 9501 31626
rect 9311 31562 9317 31574
rect 9495 31562 9501 31574
rect 9311 31510 9312 31562
rect 9500 31510 9501 31562
rect 9311 31498 9317 31510
rect 9495 31498 9501 31510
rect 9311 31446 9312 31498
rect 9500 31446 9501 31498
rect 9311 31434 9317 31446
rect 9495 31434 9501 31446
rect 9311 31382 9312 31434
rect 9500 31382 9501 31434
rect 9311 31370 9317 31382
rect 9495 31370 9501 31382
rect 9311 31318 9312 31370
rect 9500 31318 9501 31370
rect 9311 31306 9317 31318
rect 9495 31306 9501 31318
rect 9311 31254 9312 31306
rect 9500 31254 9501 31306
rect 9311 31242 9317 31254
rect 9495 31242 9501 31254
rect 9311 31190 9312 31242
rect 9500 31190 9501 31242
rect 9311 31178 9317 31190
rect 9495 31178 9501 31190
rect 9311 31126 9312 31178
rect 9500 31126 9501 31178
rect 9311 31114 9317 31126
rect 9495 31114 9501 31126
rect 9311 31062 9312 31114
rect 9500 31062 9501 31114
rect 9311 31050 9317 31062
rect 9495 31050 9501 31062
rect 9311 30998 9312 31050
rect 9500 30998 9501 31050
rect 9311 30986 9317 30998
rect 9495 30986 9501 30998
rect 9311 30934 9312 30986
rect 9500 30934 9501 30986
rect 9311 30922 9317 30934
rect 9495 30922 9501 30934
rect 9311 30870 9312 30922
rect 9500 30870 9501 30922
rect 9311 30858 9317 30870
rect 9495 30858 9501 30870
rect 9311 30806 9312 30858
rect 9500 30806 9501 30858
rect 9311 30794 9317 30806
rect 9495 30794 9501 30806
rect 9311 30742 9312 30794
rect 9500 30742 9501 30794
rect 9311 30729 9317 30742
rect 9495 30729 9501 30742
rect 9311 30677 9312 30729
rect 9500 30677 9501 30729
rect 9311 30664 9317 30677
rect 9495 30664 9501 30677
rect 9311 30612 9312 30664
rect 9500 30612 9501 30664
rect 9311 30599 9317 30612
rect 9495 30599 9501 30612
rect 9311 30547 9312 30599
rect 9500 30547 9501 30599
rect 9311 30534 9317 30547
rect 9495 30534 9501 30547
rect 9311 30482 9312 30534
rect 9500 30482 9501 30534
rect 9311 30469 9317 30482
rect 9495 30469 9501 30482
rect 9311 30417 9312 30469
rect 9500 30417 9501 30469
rect 9311 30404 9317 30417
rect 9495 30404 9501 30417
rect 9311 30352 9312 30404
rect 9500 30352 9501 30404
rect 9311 30339 9317 30352
rect 9495 30339 9501 30352
rect 9311 30287 9312 30339
rect 9500 30287 9501 30339
rect 9311 30274 9317 30287
rect 9495 30274 9501 30287
rect 9311 30222 9312 30274
rect 9500 30222 9501 30274
rect 9311 30209 9317 30222
rect 9495 30209 9501 30222
rect 9311 30157 9312 30209
rect 9500 30157 9501 30209
rect 9311 30144 9317 30157
rect 9495 30144 9501 30157
rect 9311 30092 9312 30144
rect 9500 30092 9501 30144
rect 9311 30079 9317 30092
rect 9495 30079 9501 30092
rect 9311 30027 9312 30079
rect 9500 30027 9501 30079
rect 9311 30014 9317 30027
rect 9495 30014 9501 30027
rect 9311 29962 9312 30014
rect 9500 29962 9501 30014
rect 9311 27903 9317 29962
rect 9495 27903 9501 29962
rect 9311 27153 9501 27903
rect 9311 27090 9317 27153
rect 9495 27090 9501 27153
rect 9311 27038 9312 27090
rect 9500 27038 9501 27090
rect 9311 27026 9317 27038
rect 9495 27026 9501 27038
rect 9311 26974 9312 27026
rect 9500 26974 9501 27026
rect 9311 26962 9317 26974
rect 9495 26962 9501 26974
rect 9311 26910 9312 26962
rect 9500 26910 9501 26962
rect 9311 26898 9317 26910
rect 9495 26898 9501 26910
rect 9311 26846 9312 26898
rect 9500 26846 9501 26898
rect 9311 26834 9317 26846
rect 9495 26834 9501 26846
rect 9311 26782 9312 26834
rect 9500 26782 9501 26834
rect 9311 26770 9317 26782
rect 9495 26770 9501 26782
rect 9311 26718 9312 26770
rect 9500 26718 9501 26770
rect 9311 26706 9317 26718
rect 9495 26706 9501 26718
rect 9311 26654 9312 26706
rect 9500 26654 9501 26706
rect 9311 26642 9317 26654
rect 9495 26642 9501 26654
rect 9311 26590 9312 26642
rect 9500 26590 9501 26642
rect 9311 26578 9317 26590
rect 9495 26578 9501 26590
rect 9311 26526 9312 26578
rect 9500 26526 9501 26578
rect 9311 26514 9317 26526
rect 9495 26514 9501 26526
rect 9311 26462 9312 26514
rect 9500 26462 9501 26514
rect 9311 26450 9317 26462
rect 9495 26450 9501 26462
rect 9311 26398 9312 26450
rect 9500 26398 9501 26450
rect 9311 26386 9317 26398
rect 9495 26386 9501 26398
rect 9311 26334 9312 26386
rect 9500 26334 9501 26386
rect 9311 26322 9317 26334
rect 9495 26322 9501 26334
rect 9311 26270 9312 26322
rect 9500 26270 9501 26322
rect 9311 26258 9317 26270
rect 9495 26258 9501 26270
rect 9311 26206 9312 26258
rect 9500 26206 9501 26258
rect 9311 26194 9317 26206
rect 9495 26194 9501 26206
rect 9311 26142 9312 26194
rect 9500 26142 9501 26194
rect 9311 26129 9317 26142
rect 9495 26129 9501 26142
rect 9311 26077 9312 26129
rect 9500 26077 9501 26129
rect 9311 26064 9317 26077
rect 9495 26064 9501 26077
rect 9311 26012 9312 26064
rect 9500 26012 9501 26064
rect 9311 25999 9317 26012
rect 9495 25999 9501 26012
rect 9311 25947 9312 25999
rect 9500 25947 9501 25999
rect 9311 25934 9317 25947
rect 9495 25934 9501 25947
rect 9311 25882 9312 25934
rect 9500 25882 9501 25934
rect 9311 25869 9317 25882
rect 9495 25869 9501 25882
rect 9311 25817 9312 25869
rect 9500 25817 9501 25869
rect 9311 25804 9317 25817
rect 9495 25804 9501 25817
rect 9311 25752 9312 25804
rect 9500 25752 9501 25804
rect 9311 25739 9317 25752
rect 9495 25739 9501 25752
rect 9311 25687 9312 25739
rect 9500 25687 9501 25739
rect 9311 25674 9317 25687
rect 9495 25674 9501 25687
rect 9311 25622 9312 25674
rect 9500 25622 9501 25674
rect 9311 25609 9317 25622
rect 9495 25609 9501 25622
rect 9311 25557 9312 25609
rect 9500 25557 9501 25609
rect 9311 25544 9317 25557
rect 9495 25544 9501 25557
rect 9311 25492 9312 25544
rect 9500 25492 9501 25544
rect 9311 25479 9317 25492
rect 9495 25479 9501 25492
rect 9311 25427 9312 25479
rect 9500 25427 9501 25479
rect 9311 25414 9317 25427
rect 9495 25414 9501 25427
rect 9311 25362 9312 25414
rect 9500 25362 9501 25414
rect 9311 23303 9317 25362
rect 9495 23303 9501 25362
rect 9311 22562 9501 23303
rect 9311 22490 9317 22562
rect 9495 22490 9501 22562
rect 9311 22438 9312 22490
rect 9500 22438 9501 22490
rect 9311 22426 9317 22438
rect 9495 22426 9501 22438
rect 9311 22374 9312 22426
rect 9500 22374 9501 22426
rect 9311 22362 9317 22374
rect 9495 22362 9501 22374
rect 9311 22310 9312 22362
rect 9500 22310 9501 22362
rect 9311 22298 9317 22310
rect 9495 22298 9501 22310
rect 9311 22246 9312 22298
rect 9500 22246 9501 22298
rect 9311 22234 9317 22246
rect 9495 22234 9501 22246
rect 9311 22182 9312 22234
rect 9500 22182 9501 22234
rect 9311 22170 9317 22182
rect 9495 22170 9501 22182
rect 9311 22118 9312 22170
rect 9500 22118 9501 22170
rect 9311 22106 9317 22118
rect 9495 22106 9501 22118
rect 9311 22054 9312 22106
rect 9500 22054 9501 22106
rect 9311 22042 9317 22054
rect 9495 22042 9501 22054
rect 9311 21990 9312 22042
rect 9500 21990 9501 22042
rect 9311 21978 9317 21990
rect 9495 21978 9501 21990
rect 9311 21926 9312 21978
rect 9500 21926 9501 21978
rect 9311 21914 9317 21926
rect 9495 21914 9501 21926
rect 9311 21862 9312 21914
rect 9500 21862 9501 21914
rect 9311 21850 9317 21862
rect 9495 21850 9501 21862
rect 9311 21798 9312 21850
rect 9500 21798 9501 21850
rect 9311 21786 9317 21798
rect 9495 21786 9501 21798
rect 9311 21734 9312 21786
rect 9500 21734 9501 21786
rect 9311 21722 9317 21734
rect 9495 21722 9501 21734
rect 9311 21670 9312 21722
rect 9500 21670 9501 21722
rect 9311 21658 9317 21670
rect 9495 21658 9501 21670
rect 9311 21606 9312 21658
rect 9500 21606 9501 21658
rect 9311 21594 9317 21606
rect 9495 21594 9501 21606
rect 9311 21542 9312 21594
rect 9500 21542 9501 21594
rect 9311 21529 9317 21542
rect 9495 21529 9501 21542
rect 9311 21477 9312 21529
rect 9500 21477 9501 21529
rect 9311 21464 9317 21477
rect 9495 21464 9501 21477
rect 9311 21412 9312 21464
rect 9500 21412 9501 21464
rect 9311 21399 9317 21412
rect 9495 21399 9501 21412
rect 9311 21347 9312 21399
rect 9500 21347 9501 21399
rect 9311 21334 9317 21347
rect 9495 21334 9501 21347
rect 9311 21282 9312 21334
rect 9500 21282 9501 21334
rect 9311 21269 9317 21282
rect 9495 21269 9501 21282
rect 9311 21217 9312 21269
rect 9500 21217 9501 21269
rect 9311 21204 9317 21217
rect 9495 21204 9501 21217
rect 9311 21152 9312 21204
rect 9500 21152 9501 21204
rect 9311 21139 9317 21152
rect 9495 21139 9501 21152
rect 9311 21087 9312 21139
rect 9500 21087 9501 21139
rect 9311 21074 9317 21087
rect 9495 21074 9501 21087
rect 9311 21022 9312 21074
rect 9500 21022 9501 21074
rect 9311 21009 9317 21022
rect 9495 21009 9501 21022
rect 9311 20957 9312 21009
rect 9500 20957 9501 21009
rect 9311 20944 9317 20957
rect 9495 20944 9501 20957
rect 9311 20892 9312 20944
rect 9500 20892 9501 20944
rect 9311 20879 9317 20892
rect 9495 20879 9501 20892
rect 9311 20827 9312 20879
rect 9500 20827 9501 20879
rect 9311 20814 9317 20827
rect 9495 20814 9501 20827
rect 9311 20762 9312 20814
rect 9500 20762 9501 20814
rect 9311 19360 9317 20762
rect 9495 19360 9501 20762
rect 9311 19321 9501 19360
rect 9311 19287 9317 19321
rect 9351 19287 9389 19321
rect 9423 19287 9461 19321
rect 9495 19287 9501 19321
rect 9311 19248 9501 19287
rect 9311 19214 9317 19248
rect 9351 19214 9389 19248
rect 9423 19214 9461 19248
rect 9495 19214 9501 19248
rect 9311 19175 9501 19214
rect 9311 19141 9317 19175
rect 9351 19141 9389 19175
rect 9423 19141 9461 19175
rect 9495 19141 9501 19175
rect 9311 19102 9501 19141
rect 9311 19068 9317 19102
rect 9351 19068 9389 19102
rect 9423 19068 9461 19102
rect 9495 19068 9501 19102
rect 9311 19029 9501 19068
rect 9311 18995 9317 19029
rect 9351 18995 9389 19029
rect 9423 18995 9461 19029
rect 9495 18995 9501 19029
rect 9311 18956 9501 18995
rect 9311 18922 9317 18956
rect 9351 18922 9389 18956
rect 9423 18922 9461 18956
rect 9495 18922 9501 18956
rect 9311 18883 9501 18922
rect 9311 18849 9317 18883
rect 9351 18849 9389 18883
rect 9423 18849 9461 18883
rect 9495 18849 9501 18883
rect 9311 18810 9501 18849
rect 9311 18776 9317 18810
rect 9351 18776 9389 18810
rect 9423 18776 9461 18810
rect 9495 18776 9501 18810
rect 9311 18737 9501 18776
rect 9311 18703 9317 18737
rect 9351 18703 9389 18737
rect 9423 18703 9461 18737
rect 9495 18703 9501 18737
rect 9311 17953 9501 18703
rect 9311 17890 9317 17953
rect 9495 17890 9501 17953
rect 9311 17838 9312 17890
rect 9500 17838 9501 17890
rect 9311 17826 9317 17838
rect 9495 17826 9501 17838
rect 9311 17774 9312 17826
rect 9500 17774 9501 17826
rect 9311 17762 9317 17774
rect 9495 17762 9501 17774
rect 9311 17710 9312 17762
rect 9500 17710 9501 17762
rect 9311 17698 9317 17710
rect 9495 17698 9501 17710
rect 9311 17646 9312 17698
rect 9500 17646 9501 17698
rect 9311 17634 9317 17646
rect 9495 17634 9501 17646
rect 9311 17582 9312 17634
rect 9500 17582 9501 17634
rect 9311 17570 9317 17582
rect 9495 17570 9501 17582
rect 9311 17518 9312 17570
rect 9500 17518 9501 17570
rect 9311 17506 9317 17518
rect 9495 17506 9501 17518
rect 9311 17454 9312 17506
rect 9500 17454 9501 17506
rect 9311 17442 9317 17454
rect 9495 17442 9501 17454
rect 9311 17390 9312 17442
rect 9500 17390 9501 17442
rect 9311 17378 9317 17390
rect 9495 17378 9501 17390
rect 9311 17326 9312 17378
rect 9500 17326 9501 17378
rect 9311 17314 9317 17326
rect 9495 17314 9501 17326
rect 9311 17262 9312 17314
rect 9500 17262 9501 17314
rect 9311 17250 9317 17262
rect 9495 17250 9501 17262
rect 9311 17198 9312 17250
rect 9500 17198 9501 17250
rect 9311 17186 9317 17198
rect 9495 17186 9501 17198
rect 9311 17134 9312 17186
rect 9500 17134 9501 17186
rect 9311 17122 9317 17134
rect 9495 17122 9501 17134
rect 9311 17070 9312 17122
rect 9500 17070 9501 17122
rect 9311 17058 9317 17070
rect 9495 17058 9501 17070
rect 9311 17006 9312 17058
rect 9500 17006 9501 17058
rect 9311 16994 9317 17006
rect 9495 16994 9501 17006
rect 9311 16942 9312 16994
rect 9500 16942 9501 16994
rect 9311 16929 9317 16942
rect 9495 16929 9501 16942
rect 9311 16877 9312 16929
rect 9500 16877 9501 16929
rect 9311 16864 9317 16877
rect 9495 16864 9501 16877
rect 9311 16812 9312 16864
rect 9500 16812 9501 16864
rect 9311 16799 9317 16812
rect 9495 16799 9501 16812
rect 9311 16747 9312 16799
rect 9500 16747 9501 16799
rect 9311 16734 9317 16747
rect 9495 16734 9501 16747
rect 9311 16682 9312 16734
rect 9500 16682 9501 16734
rect 9311 16669 9317 16682
rect 9495 16669 9501 16682
rect 9311 16617 9312 16669
rect 9500 16617 9501 16669
rect 9311 16604 9317 16617
rect 9495 16604 9501 16617
rect 9311 16552 9312 16604
rect 9500 16552 9501 16604
rect 9311 16539 9317 16552
rect 9495 16539 9501 16552
rect 9311 16487 9312 16539
rect 9500 16487 9501 16539
rect 9311 16474 9317 16487
rect 9495 16474 9501 16487
rect 9311 16422 9312 16474
rect 9500 16422 9501 16474
rect 9311 16409 9317 16422
rect 9495 16409 9501 16422
rect 9311 16357 9312 16409
rect 9500 16357 9501 16409
rect 9311 16344 9317 16357
rect 9495 16344 9501 16357
rect 9311 16292 9312 16344
rect 9500 16292 9501 16344
rect 9311 16279 9317 16292
rect 9495 16279 9501 16292
rect 9311 16227 9312 16279
rect 9500 16227 9501 16279
rect 9311 16214 9317 16227
rect 9495 16214 9501 16227
rect 9311 16162 9312 16214
rect 9500 16162 9501 16214
rect 9311 14103 9317 16162
rect 9495 14103 9501 16162
rect 9311 13362 9501 14103
rect 9311 13290 9317 13362
rect 9495 13290 9501 13362
rect 9311 13238 9312 13290
rect 9500 13238 9501 13290
rect 9311 13226 9317 13238
rect 9495 13226 9501 13238
rect 9311 13174 9312 13226
rect 9500 13174 9501 13226
rect 9311 13162 9317 13174
rect 9495 13162 9501 13174
rect 9311 13110 9312 13162
rect 9500 13110 9501 13162
rect 9311 13098 9317 13110
rect 9495 13098 9501 13110
rect 9311 13046 9312 13098
rect 9500 13046 9501 13098
rect 9311 13034 9317 13046
rect 9495 13034 9501 13046
rect 9311 12982 9312 13034
rect 9500 12982 9501 13034
rect 9311 12970 9317 12982
rect 9495 12970 9501 12982
rect 9311 12918 9312 12970
rect 9500 12918 9501 12970
rect 9311 12906 9317 12918
rect 9495 12906 9501 12918
rect 9311 12854 9312 12906
rect 9500 12854 9501 12906
rect 9311 12842 9317 12854
rect 9495 12842 9501 12854
rect 9311 12790 9312 12842
rect 9500 12790 9501 12842
rect 9311 12778 9317 12790
rect 9495 12778 9501 12790
rect 9311 12726 9312 12778
rect 9500 12726 9501 12778
rect 9311 12714 9317 12726
rect 9495 12714 9501 12726
rect 9311 12662 9312 12714
rect 9500 12662 9501 12714
rect 9311 12650 9317 12662
rect 9495 12650 9501 12662
rect 9311 12598 9312 12650
rect 9500 12598 9501 12650
rect 9311 12586 9317 12598
rect 9495 12586 9501 12598
rect 9311 12534 9312 12586
rect 9500 12534 9501 12586
rect 9311 12522 9317 12534
rect 9495 12522 9501 12534
rect 9311 12470 9312 12522
rect 9500 12470 9501 12522
rect 9311 12458 9317 12470
rect 9495 12458 9501 12470
rect 9311 12406 9312 12458
rect 9500 12406 9501 12458
rect 9311 12394 9317 12406
rect 9495 12394 9501 12406
rect 9311 12342 9312 12394
rect 9500 12342 9501 12394
rect 9311 12329 9317 12342
rect 9495 12329 9501 12342
rect 9311 12277 9312 12329
rect 9500 12277 9501 12329
rect 9311 12264 9317 12277
rect 9495 12264 9501 12277
rect 9311 12212 9312 12264
rect 9500 12212 9501 12264
rect 9311 12199 9317 12212
rect 9495 12199 9501 12212
rect 9311 12147 9312 12199
rect 9500 12147 9501 12199
rect 9311 12134 9317 12147
rect 9495 12134 9501 12147
rect 9311 12082 9312 12134
rect 9500 12082 9501 12134
rect 9311 12069 9317 12082
rect 9495 12069 9501 12082
rect 9311 12017 9312 12069
rect 9500 12017 9501 12069
rect 9311 12004 9317 12017
rect 9495 12004 9501 12017
rect 9311 11952 9312 12004
rect 9500 11952 9501 12004
rect 9311 11939 9317 11952
rect 9495 11939 9501 11952
rect 9311 11887 9312 11939
rect 9500 11887 9501 11939
rect 9311 11874 9317 11887
rect 9495 11874 9501 11887
rect 9311 11822 9312 11874
rect 9500 11822 9501 11874
rect 9311 11809 9317 11822
rect 9495 11809 9501 11822
rect 9311 11757 9312 11809
rect 9500 11757 9501 11809
rect 9311 11744 9317 11757
rect 9495 11744 9501 11757
rect 9311 11692 9312 11744
rect 9500 11692 9501 11744
rect 9311 11679 9317 11692
rect 9495 11679 9501 11692
rect 9311 11627 9312 11679
rect 9500 11627 9501 11679
rect 9311 11614 9317 11627
rect 9495 11614 9501 11627
rect 9311 11562 9312 11614
rect 9500 11562 9501 11614
rect 9311 10160 9317 11562
rect 9495 10160 9501 11562
rect 9311 10121 9501 10160
rect 9311 10087 9317 10121
rect 9351 10087 9389 10121
rect 9423 10087 9461 10121
rect 9495 10087 9501 10121
rect 9311 10048 9501 10087
rect 9311 10014 9317 10048
rect 9351 10014 9389 10048
rect 9423 10014 9461 10048
rect 9495 10014 9501 10048
rect 9311 9975 9501 10014
rect 9311 9941 9317 9975
rect 9351 9941 9389 9975
rect 9423 9941 9461 9975
rect 9495 9941 9501 9975
rect 9311 9902 9501 9941
rect 9311 9868 9317 9902
rect 9351 9868 9389 9902
rect 9423 9868 9461 9902
rect 9495 9868 9501 9902
rect 9311 9829 9501 9868
rect 9311 9795 9317 9829
rect 9351 9795 9389 9829
rect 9423 9795 9461 9829
rect 9495 9795 9501 9829
rect 9311 9756 9501 9795
rect 9311 9722 9317 9756
rect 9351 9722 9389 9756
rect 9423 9722 9461 9756
rect 9495 9722 9501 9756
rect 9311 9683 9501 9722
rect 9311 9649 9317 9683
rect 9351 9649 9389 9683
rect 9423 9649 9461 9683
rect 9495 9649 9501 9683
rect 9311 9610 9501 9649
rect 9311 9576 9317 9610
rect 9351 9576 9389 9610
rect 9423 9576 9461 9610
rect 9495 9576 9501 9610
rect 9311 9537 9501 9576
rect 9311 9503 9317 9537
rect 9351 9503 9389 9537
rect 9423 9503 9461 9537
rect 9495 9503 9501 9537
rect 9311 9491 9501 9503
rect 9801 37997 9931 38003
rect 9853 37945 9879 37997
rect 9801 37929 9931 37945
rect 9853 37877 9879 37929
rect 9801 37861 9931 37877
rect 9853 37809 9879 37861
rect 9801 37793 9931 37809
rect 9853 37741 9879 37793
rect 9801 37725 9931 37741
rect 9853 37673 9879 37725
rect 9801 37657 9931 37673
rect 9853 37605 9879 37657
rect 9801 37589 9931 37605
rect 9853 37537 9879 37589
rect 9801 37521 9931 37537
rect 9853 37469 9879 37521
rect 9801 37453 9931 37469
rect 9853 37401 9879 37453
rect 9801 37385 9931 37401
rect 9853 37333 9879 37385
rect 9801 37318 9931 37333
rect 9853 37266 9879 37318
rect 9801 37251 9931 37266
rect 9853 37199 9879 37251
rect 9801 37184 9931 37199
rect 9853 37132 9879 37184
rect 9801 37117 9931 37132
rect 9853 37065 9879 37117
rect 9801 34225 9931 37065
rect 9853 34173 9879 34225
rect 9801 34161 9931 34173
rect 9853 34109 9879 34161
rect 9801 34097 9931 34109
rect 9853 34045 9879 34097
rect 9801 34033 9931 34045
rect 9853 33981 9879 34033
rect 9801 33969 9931 33981
rect 9853 33917 9879 33969
rect 9801 33905 9931 33917
rect 9853 33853 9879 33905
rect 9801 33841 9931 33853
rect 9853 33789 9879 33841
rect 9801 33777 9931 33789
rect 9853 33725 9879 33777
rect 9801 33713 9931 33725
rect 9853 33661 9879 33713
rect 9801 33649 9931 33661
rect 9853 33597 9879 33649
rect 9801 33585 9931 33597
rect 9853 33533 9879 33585
rect 9801 33521 9931 33533
rect 9853 33469 9879 33521
rect 9801 33457 9931 33469
rect 9853 33405 9879 33457
rect 9801 33393 9931 33405
rect 9853 33341 9879 33393
rect 9801 33329 9931 33341
rect 9853 33277 9879 33329
rect 9801 33264 9931 33277
rect 9853 33212 9879 33264
rect 9801 33199 9931 33212
rect 9853 33147 9879 33199
rect 9801 33134 9931 33147
rect 9853 33082 9879 33134
rect 9801 33069 9931 33082
rect 9853 33017 9879 33069
rect 9801 33004 9931 33017
rect 9853 32952 9879 33004
rect 9801 32939 9931 32952
rect 9853 32887 9879 32939
rect 9801 32874 9931 32887
rect 9853 32822 9879 32874
rect 9801 32809 9931 32822
rect 9853 32757 9879 32809
rect 9801 32744 9931 32757
rect 9853 32692 9879 32744
rect 9801 32679 9931 32692
rect 9853 32627 9879 32679
rect 9801 32614 9931 32627
rect 9853 32562 9879 32614
rect 9801 32549 9931 32562
rect 9853 32497 9879 32549
rect 9801 29625 9931 32497
rect 9853 29573 9879 29625
rect 9801 29561 9931 29573
rect 9853 29509 9879 29561
rect 9801 29497 9931 29509
rect 9853 29445 9879 29497
rect 9801 29433 9931 29445
rect 9853 29381 9879 29433
rect 9801 29369 9931 29381
rect 9853 29317 9879 29369
rect 9801 29305 9931 29317
rect 9853 29253 9879 29305
rect 9801 29241 9931 29253
rect 9853 29189 9879 29241
rect 9801 29177 9931 29189
rect 9853 29125 9879 29177
rect 9801 29113 9931 29125
rect 9853 29061 9879 29113
rect 9801 29049 9931 29061
rect 9853 28997 9879 29049
rect 9801 28985 9931 28997
rect 9853 28933 9879 28985
rect 9801 28921 9931 28933
rect 9853 28869 9879 28921
rect 9801 28857 9931 28869
rect 9853 28805 9879 28857
rect 9801 28793 9931 28805
rect 9853 28741 9879 28793
rect 9801 28729 9931 28741
rect 9853 28677 9879 28729
rect 9801 28664 9931 28677
rect 9853 28612 9879 28664
rect 9801 28599 9931 28612
rect 9853 28547 9879 28599
rect 9801 28534 9931 28547
rect 9853 28482 9879 28534
rect 9801 28469 9931 28482
rect 9853 28417 9879 28469
rect 9801 28404 9931 28417
rect 9853 28352 9879 28404
rect 9801 28339 9931 28352
rect 9853 28287 9879 28339
rect 9801 28274 9931 28287
rect 9853 28222 9879 28274
rect 9801 28209 9931 28222
rect 9853 28157 9879 28209
rect 9801 28144 9931 28157
rect 9853 28092 9879 28144
rect 9801 28079 9931 28092
rect 9853 28027 9879 28079
rect 9801 28014 9931 28027
rect 9853 27962 9879 28014
rect 9801 27949 9931 27962
rect 9853 27897 9879 27949
rect 9801 25025 9931 27897
rect 9853 24973 9879 25025
rect 9801 24961 9931 24973
rect 9853 24909 9879 24961
rect 9801 24897 9931 24909
rect 9853 24845 9879 24897
rect 9801 24833 9931 24845
rect 9853 24781 9879 24833
rect 9801 24769 9931 24781
rect 9853 24717 9879 24769
rect 9801 24705 9931 24717
rect 9853 24653 9879 24705
rect 9801 24641 9931 24653
rect 9853 24589 9879 24641
rect 9801 24577 9931 24589
rect 9853 24525 9879 24577
rect 9801 24513 9931 24525
rect 9853 24461 9879 24513
rect 9801 24449 9931 24461
rect 9853 24397 9879 24449
rect 9801 24385 9931 24397
rect 9853 24333 9879 24385
rect 9801 24321 9931 24333
rect 9853 24269 9879 24321
rect 9801 24257 9931 24269
rect 9853 24205 9879 24257
rect 9801 24193 9931 24205
rect 9853 24141 9879 24193
rect 9801 24129 9931 24141
rect 9853 24077 9879 24129
rect 9801 24064 9931 24077
rect 9853 24012 9879 24064
rect 9801 23999 9931 24012
rect 9853 23947 9879 23999
rect 9801 23934 9931 23947
rect 9853 23882 9879 23934
rect 9801 23869 9931 23882
rect 9853 23817 9879 23869
rect 9801 23804 9931 23817
rect 9853 23752 9879 23804
rect 9801 23739 9931 23752
rect 9853 23687 9879 23739
rect 9801 23674 9931 23687
rect 9853 23622 9879 23674
rect 9801 23609 9931 23622
rect 9853 23557 9879 23609
rect 9801 23544 9931 23557
rect 9853 23492 9879 23544
rect 9801 23479 9931 23492
rect 9853 23427 9879 23479
rect 9801 23414 9931 23427
rect 9853 23362 9879 23414
rect 9801 23349 9931 23362
rect 9853 23297 9879 23349
rect 9801 20425 9931 23297
rect 9853 20373 9879 20425
rect 9801 20361 9931 20373
rect 9853 20309 9879 20361
rect 9801 20297 9931 20309
rect 9853 20245 9879 20297
rect 9801 20233 9931 20245
rect 9853 20181 9879 20233
rect 9801 20169 9931 20181
rect 9853 20117 9879 20169
rect 9801 20105 9931 20117
rect 9853 20053 9879 20105
rect 9801 20041 9931 20053
rect 9853 19989 9879 20041
rect 9801 19977 9931 19989
rect 9853 19925 9879 19977
rect 9801 19913 9931 19925
rect 9853 19861 9879 19913
rect 9801 19849 9931 19861
rect 9853 19797 9879 19849
rect 9801 19785 9931 19797
rect 9853 19733 9879 19785
rect 9801 19721 9931 19733
rect 9853 19669 9879 19721
rect 9801 19657 9931 19669
rect 9853 19605 9879 19657
rect 9801 19593 9931 19605
rect 9853 19541 9879 19593
rect 9801 19529 9931 19541
rect 9853 19477 9879 19529
rect 9801 19464 9931 19477
rect 9853 19412 9879 19464
rect 9801 19399 9931 19412
rect 9853 19347 9879 19399
rect 9801 19334 9931 19347
rect 9853 19282 9879 19334
rect 9801 19269 9931 19282
rect 9853 19217 9879 19269
rect 9801 19204 9931 19217
rect 9853 19152 9879 19204
rect 9801 19139 9931 19152
rect 9853 19087 9879 19139
rect 9801 19074 9931 19087
rect 9853 19022 9879 19074
rect 9801 19009 9931 19022
rect 9853 18957 9879 19009
rect 9801 18944 9931 18957
rect 9853 18892 9879 18944
rect 9801 18879 9931 18892
rect 9853 18827 9879 18879
rect 9801 18814 9931 18827
rect 9853 18762 9879 18814
rect 9801 18749 9931 18762
rect 9853 18697 9879 18749
rect 9801 15825 9931 18697
rect 9853 15773 9879 15825
rect 9801 15761 9931 15773
rect 9853 15709 9879 15761
rect 9801 15697 9931 15709
rect 9853 15645 9879 15697
rect 9801 15633 9931 15645
rect 9853 15581 9879 15633
rect 9801 15569 9931 15581
rect 9853 15517 9879 15569
rect 9801 15505 9931 15517
rect 9853 15453 9879 15505
rect 9801 15441 9931 15453
rect 9853 15389 9879 15441
rect 9801 15377 9931 15389
rect 9853 15325 9879 15377
rect 9801 15313 9931 15325
rect 9853 15261 9879 15313
rect 9801 15249 9931 15261
rect 9853 15197 9879 15249
rect 9801 15185 9931 15197
rect 9853 15133 9879 15185
rect 9801 15121 9931 15133
rect 9853 15069 9879 15121
rect 9801 15057 9931 15069
rect 9853 15005 9879 15057
rect 9801 14993 9931 15005
rect 9853 14941 9879 14993
rect 9801 14929 9931 14941
rect 9853 14877 9879 14929
rect 9801 14864 9931 14877
rect 9853 14812 9879 14864
rect 9801 14799 9931 14812
rect 9853 14747 9879 14799
rect 9801 14734 9931 14747
rect 9853 14682 9879 14734
rect 9801 14669 9931 14682
rect 9853 14617 9879 14669
rect 9801 14604 9931 14617
rect 9853 14552 9879 14604
rect 9801 14539 9931 14552
rect 9853 14487 9879 14539
rect 9801 14474 9931 14487
rect 9853 14422 9879 14474
rect 9801 14409 9931 14422
rect 9853 14357 9879 14409
rect 9801 14344 9931 14357
rect 9853 14292 9879 14344
rect 9801 14279 9931 14292
rect 9853 14227 9879 14279
rect 9801 14214 9931 14227
rect 9853 14162 9879 14214
rect 9801 14149 9931 14162
rect 9853 14097 9879 14149
rect 9801 11225 9931 14097
rect 9853 11173 9879 11225
rect 9801 11161 9931 11173
rect 9853 11109 9879 11161
rect 9801 11097 9931 11109
rect 9853 11045 9879 11097
rect 9801 11033 9931 11045
rect 9853 10981 9879 11033
rect 9801 10969 9931 10981
rect 9853 10917 9879 10969
rect 9801 10905 9931 10917
rect 9853 10853 9879 10905
rect 9801 10841 9931 10853
rect 9853 10789 9879 10841
rect 9801 10777 9931 10789
rect 9853 10725 9879 10777
rect 9801 10713 9931 10725
rect 9853 10661 9879 10713
rect 9801 10649 9931 10661
rect 9853 10597 9879 10649
rect 9801 10585 9931 10597
rect 9853 10533 9879 10585
rect 9801 10521 9931 10533
rect 9853 10469 9879 10521
rect 9801 10457 9931 10469
rect 9853 10405 9879 10457
rect 9801 10393 9931 10405
rect 9853 10341 9879 10393
rect 9801 10329 9931 10341
rect 9853 10277 9879 10329
rect 9801 10264 9931 10277
rect 9853 10212 9879 10264
rect 9801 10199 9931 10212
rect 9853 10147 9879 10199
rect 9801 10134 9931 10147
rect 9853 10082 9879 10134
rect 9801 10069 9931 10082
rect 9853 10017 9879 10069
rect 9801 10004 9931 10017
rect 9853 9952 9879 10004
rect 9801 9939 9931 9952
rect 9853 9887 9879 9939
rect 9801 9874 9931 9887
rect 9853 9822 9879 9874
rect 9801 9809 9931 9822
rect 9853 9757 9879 9809
rect 9801 9744 9931 9757
rect 9853 9692 9879 9744
rect 9801 9679 9931 9692
rect 9853 9627 9879 9679
rect 9801 9614 9931 9627
rect 9853 9562 9879 9614
rect 9801 9549 9931 9562
rect 9853 9497 9879 9549
rect 9801 9491 9931 9497
rect 10231 37962 10421 38003
rect 10231 37928 10237 37962
rect 10271 37928 10309 37962
rect 10343 37928 10381 37962
rect 10415 37928 10421 37962
rect 10231 37887 10421 37928
rect 10231 37853 10237 37887
rect 10271 37853 10309 37887
rect 10343 37853 10381 37887
rect 10415 37853 10421 37887
rect 10231 37812 10421 37853
rect 10231 37778 10237 37812
rect 10271 37778 10309 37812
rect 10343 37778 10381 37812
rect 10415 37778 10421 37812
rect 10231 37737 10421 37778
rect 10231 37703 10237 37737
rect 10271 37703 10309 37737
rect 10343 37703 10381 37737
rect 10415 37703 10421 37737
rect 10231 37662 10421 37703
rect 10231 37628 10237 37662
rect 10271 37628 10309 37662
rect 10343 37628 10381 37662
rect 10415 37628 10421 37662
rect 10231 37587 10421 37628
rect 10231 37553 10237 37587
rect 10271 37553 10309 37587
rect 10343 37553 10381 37587
rect 10415 37553 10421 37587
rect 10231 37512 10421 37553
rect 10231 37478 10237 37512
rect 10271 37478 10309 37512
rect 10343 37478 10381 37512
rect 10415 37478 10421 37512
rect 10231 37437 10421 37478
rect 10231 37403 10237 37437
rect 10271 37403 10309 37437
rect 10343 37403 10381 37437
rect 10415 37403 10421 37437
rect 10231 37362 10421 37403
rect 10231 37328 10237 37362
rect 10271 37328 10309 37362
rect 10343 37328 10381 37362
rect 10415 37328 10421 37362
rect 10231 37287 10421 37328
rect 10231 37253 10237 37287
rect 10271 37253 10309 37287
rect 10343 37253 10381 37287
rect 10415 37253 10421 37287
rect 10231 37212 10421 37253
rect 10231 37178 10237 37212
rect 10271 37178 10309 37212
rect 10343 37178 10381 37212
rect 10415 37178 10421 37212
rect 10231 37137 10421 37178
rect 10231 37103 10237 37137
rect 10271 37103 10309 37137
rect 10343 37103 10381 37137
rect 10415 37103 10421 37137
rect 10231 36353 10421 37103
rect 10231 36290 10237 36353
rect 10415 36290 10421 36353
rect 10231 36238 10232 36290
rect 10420 36238 10421 36290
rect 10231 36226 10237 36238
rect 10415 36226 10421 36238
rect 10231 36174 10232 36226
rect 10420 36174 10421 36226
rect 10231 36162 10237 36174
rect 10415 36162 10421 36174
rect 10231 36110 10232 36162
rect 10420 36110 10421 36162
rect 10231 36098 10237 36110
rect 10415 36098 10421 36110
rect 10231 36046 10232 36098
rect 10420 36046 10421 36098
rect 10231 36034 10237 36046
rect 10415 36034 10421 36046
rect 10231 35982 10232 36034
rect 10420 35982 10421 36034
rect 10231 35970 10237 35982
rect 10415 35970 10421 35982
rect 10231 35918 10232 35970
rect 10420 35918 10421 35970
rect 10231 35906 10237 35918
rect 10415 35906 10421 35918
rect 10231 35854 10232 35906
rect 10420 35854 10421 35906
rect 10231 35842 10237 35854
rect 10415 35842 10421 35854
rect 10231 35790 10232 35842
rect 10420 35790 10421 35842
rect 10231 35778 10237 35790
rect 10415 35778 10421 35790
rect 10231 35726 10232 35778
rect 10420 35726 10421 35778
rect 10231 35714 10237 35726
rect 10415 35714 10421 35726
rect 10231 35662 10232 35714
rect 10420 35662 10421 35714
rect 10231 35650 10237 35662
rect 10415 35650 10421 35662
rect 10231 35598 10232 35650
rect 10420 35598 10421 35650
rect 10231 35586 10237 35598
rect 10415 35586 10421 35598
rect 10231 35534 10232 35586
rect 10420 35534 10421 35586
rect 10231 35522 10237 35534
rect 10415 35522 10421 35534
rect 10231 35470 10232 35522
rect 10420 35470 10421 35522
rect 10231 35458 10237 35470
rect 10415 35458 10421 35470
rect 10231 35406 10232 35458
rect 10420 35406 10421 35458
rect 10231 35394 10237 35406
rect 10415 35394 10421 35406
rect 10231 35342 10232 35394
rect 10420 35342 10421 35394
rect 10231 35329 10237 35342
rect 10415 35329 10421 35342
rect 10231 35277 10232 35329
rect 10420 35277 10421 35329
rect 10231 35264 10237 35277
rect 10415 35264 10421 35277
rect 10231 35212 10232 35264
rect 10420 35212 10421 35264
rect 10231 35199 10237 35212
rect 10415 35199 10421 35212
rect 10231 35147 10232 35199
rect 10420 35147 10421 35199
rect 10231 35134 10237 35147
rect 10415 35134 10421 35147
rect 10231 35082 10232 35134
rect 10420 35082 10421 35134
rect 10231 35069 10237 35082
rect 10415 35069 10421 35082
rect 10231 35017 10232 35069
rect 10420 35017 10421 35069
rect 10231 35004 10237 35017
rect 10415 35004 10421 35017
rect 10231 34952 10232 35004
rect 10420 34952 10421 35004
rect 10231 34939 10237 34952
rect 10415 34939 10421 34952
rect 10231 34887 10232 34939
rect 10420 34887 10421 34939
rect 10231 34874 10237 34887
rect 10415 34874 10421 34887
rect 10231 34822 10232 34874
rect 10420 34822 10421 34874
rect 10231 34809 10237 34822
rect 10415 34809 10421 34822
rect 10231 34757 10232 34809
rect 10420 34757 10421 34809
rect 10231 34744 10237 34757
rect 10415 34744 10421 34757
rect 10231 34692 10232 34744
rect 10420 34692 10421 34744
rect 10231 34679 10237 34692
rect 10415 34679 10421 34692
rect 10231 34627 10232 34679
rect 10420 34627 10421 34679
rect 10231 34614 10237 34627
rect 10415 34614 10421 34627
rect 10231 34562 10232 34614
rect 10420 34562 10421 34614
rect 10231 32503 10237 34562
rect 10415 32503 10421 34562
rect 10231 31753 10421 32503
rect 10231 31690 10237 31753
rect 10415 31690 10421 31753
rect 10231 31638 10232 31690
rect 10420 31638 10421 31690
rect 10231 31626 10237 31638
rect 10415 31626 10421 31638
rect 10231 31574 10232 31626
rect 10420 31574 10421 31626
rect 10231 31562 10237 31574
rect 10415 31562 10421 31574
rect 10231 31510 10232 31562
rect 10420 31510 10421 31562
rect 10231 31498 10237 31510
rect 10415 31498 10421 31510
rect 10231 31446 10232 31498
rect 10420 31446 10421 31498
rect 10231 31434 10237 31446
rect 10415 31434 10421 31446
rect 10231 31382 10232 31434
rect 10420 31382 10421 31434
rect 10231 31370 10237 31382
rect 10415 31370 10421 31382
rect 10231 31318 10232 31370
rect 10420 31318 10421 31370
rect 10231 31306 10237 31318
rect 10415 31306 10421 31318
rect 10231 31254 10232 31306
rect 10420 31254 10421 31306
rect 10231 31242 10237 31254
rect 10415 31242 10421 31254
rect 10231 31190 10232 31242
rect 10420 31190 10421 31242
rect 10231 31178 10237 31190
rect 10415 31178 10421 31190
rect 10231 31126 10232 31178
rect 10420 31126 10421 31178
rect 10231 31114 10237 31126
rect 10415 31114 10421 31126
rect 10231 31062 10232 31114
rect 10420 31062 10421 31114
rect 10231 31050 10237 31062
rect 10415 31050 10421 31062
rect 10231 30998 10232 31050
rect 10420 30998 10421 31050
rect 10231 30986 10237 30998
rect 10415 30986 10421 30998
rect 10231 30934 10232 30986
rect 10420 30934 10421 30986
rect 10231 30922 10237 30934
rect 10415 30922 10421 30934
rect 10231 30870 10232 30922
rect 10420 30870 10421 30922
rect 10231 30858 10237 30870
rect 10415 30858 10421 30870
rect 10231 30806 10232 30858
rect 10420 30806 10421 30858
rect 10231 30794 10237 30806
rect 10415 30794 10421 30806
rect 10231 30742 10232 30794
rect 10420 30742 10421 30794
rect 10231 30729 10237 30742
rect 10415 30729 10421 30742
rect 10231 30677 10232 30729
rect 10420 30677 10421 30729
rect 10231 30664 10237 30677
rect 10415 30664 10421 30677
rect 10231 30612 10232 30664
rect 10420 30612 10421 30664
rect 10231 30599 10237 30612
rect 10415 30599 10421 30612
rect 10231 30547 10232 30599
rect 10420 30547 10421 30599
rect 10231 30534 10237 30547
rect 10415 30534 10421 30547
rect 10231 30482 10232 30534
rect 10420 30482 10421 30534
rect 10231 30469 10237 30482
rect 10415 30469 10421 30482
rect 10231 30417 10232 30469
rect 10420 30417 10421 30469
rect 10231 30404 10237 30417
rect 10415 30404 10421 30417
rect 10231 30352 10232 30404
rect 10420 30352 10421 30404
rect 10231 30339 10237 30352
rect 10415 30339 10421 30352
rect 10231 30287 10232 30339
rect 10420 30287 10421 30339
rect 10231 30274 10237 30287
rect 10415 30274 10421 30287
rect 10231 30222 10232 30274
rect 10420 30222 10421 30274
rect 10231 30209 10237 30222
rect 10415 30209 10421 30222
rect 10231 30157 10232 30209
rect 10420 30157 10421 30209
rect 10231 30144 10237 30157
rect 10415 30144 10421 30157
rect 10231 30092 10232 30144
rect 10420 30092 10421 30144
rect 10231 30079 10237 30092
rect 10415 30079 10421 30092
rect 10231 30027 10232 30079
rect 10420 30027 10421 30079
rect 10231 30014 10237 30027
rect 10415 30014 10421 30027
rect 10231 29962 10232 30014
rect 10420 29962 10421 30014
rect 10231 27903 10237 29962
rect 10415 27903 10421 29962
rect 10231 27153 10421 27903
rect 10231 27090 10237 27153
rect 10415 27090 10421 27153
rect 10231 27038 10232 27090
rect 10420 27038 10421 27090
rect 10231 27026 10237 27038
rect 10415 27026 10421 27038
rect 10231 26974 10232 27026
rect 10420 26974 10421 27026
rect 10231 26962 10237 26974
rect 10415 26962 10421 26974
rect 10231 26910 10232 26962
rect 10420 26910 10421 26962
rect 10231 26898 10237 26910
rect 10415 26898 10421 26910
rect 10231 26846 10232 26898
rect 10420 26846 10421 26898
rect 10231 26834 10237 26846
rect 10415 26834 10421 26846
rect 10231 26782 10232 26834
rect 10420 26782 10421 26834
rect 10231 26770 10237 26782
rect 10415 26770 10421 26782
rect 10231 26718 10232 26770
rect 10420 26718 10421 26770
rect 10231 26706 10237 26718
rect 10415 26706 10421 26718
rect 10231 26654 10232 26706
rect 10420 26654 10421 26706
rect 10231 26642 10237 26654
rect 10415 26642 10421 26654
rect 10231 26590 10232 26642
rect 10420 26590 10421 26642
rect 10231 26578 10237 26590
rect 10415 26578 10421 26590
rect 10231 26526 10232 26578
rect 10420 26526 10421 26578
rect 10231 26514 10237 26526
rect 10415 26514 10421 26526
rect 10231 26462 10232 26514
rect 10420 26462 10421 26514
rect 10231 26450 10237 26462
rect 10415 26450 10421 26462
rect 10231 26398 10232 26450
rect 10420 26398 10421 26450
rect 10231 26386 10237 26398
rect 10415 26386 10421 26398
rect 10231 26334 10232 26386
rect 10420 26334 10421 26386
rect 10231 26322 10237 26334
rect 10415 26322 10421 26334
rect 10231 26270 10232 26322
rect 10420 26270 10421 26322
rect 10231 26258 10237 26270
rect 10415 26258 10421 26270
rect 10231 26206 10232 26258
rect 10420 26206 10421 26258
rect 10231 26194 10237 26206
rect 10415 26194 10421 26206
rect 10231 26142 10232 26194
rect 10420 26142 10421 26194
rect 10231 26129 10237 26142
rect 10415 26129 10421 26142
rect 10231 26077 10232 26129
rect 10420 26077 10421 26129
rect 10231 26064 10237 26077
rect 10415 26064 10421 26077
rect 10231 26012 10232 26064
rect 10420 26012 10421 26064
rect 10231 25999 10237 26012
rect 10415 25999 10421 26012
rect 10231 25947 10232 25999
rect 10420 25947 10421 25999
rect 10231 25934 10237 25947
rect 10415 25934 10421 25947
rect 10231 25882 10232 25934
rect 10420 25882 10421 25934
rect 10231 25869 10237 25882
rect 10415 25869 10421 25882
rect 10231 25817 10232 25869
rect 10420 25817 10421 25869
rect 10231 25804 10237 25817
rect 10415 25804 10421 25817
rect 10231 25752 10232 25804
rect 10420 25752 10421 25804
rect 10231 25739 10237 25752
rect 10415 25739 10421 25752
rect 10231 25687 10232 25739
rect 10420 25687 10421 25739
rect 10231 25674 10237 25687
rect 10415 25674 10421 25687
rect 10231 25622 10232 25674
rect 10420 25622 10421 25674
rect 10231 25609 10237 25622
rect 10415 25609 10421 25622
rect 10231 25557 10232 25609
rect 10420 25557 10421 25609
rect 10231 25544 10237 25557
rect 10415 25544 10421 25557
rect 10231 25492 10232 25544
rect 10420 25492 10421 25544
rect 10231 25479 10237 25492
rect 10415 25479 10421 25492
rect 10231 25427 10232 25479
rect 10420 25427 10421 25479
rect 10231 25414 10237 25427
rect 10415 25414 10421 25427
rect 10231 25362 10232 25414
rect 10420 25362 10421 25414
rect 10231 23303 10237 25362
rect 10415 23303 10421 25362
rect 10231 22562 10421 23303
rect 10231 22490 10237 22562
rect 10415 22490 10421 22562
rect 10231 22438 10232 22490
rect 10420 22438 10421 22490
rect 10231 22426 10237 22438
rect 10415 22426 10421 22438
rect 10231 22374 10232 22426
rect 10420 22374 10421 22426
rect 10231 22362 10237 22374
rect 10415 22362 10421 22374
rect 10231 22310 10232 22362
rect 10420 22310 10421 22362
rect 10231 22298 10237 22310
rect 10415 22298 10421 22310
rect 10231 22246 10232 22298
rect 10420 22246 10421 22298
rect 10231 22234 10237 22246
rect 10415 22234 10421 22246
rect 10231 22182 10232 22234
rect 10420 22182 10421 22234
rect 10231 22170 10237 22182
rect 10415 22170 10421 22182
rect 10231 22118 10232 22170
rect 10420 22118 10421 22170
rect 10231 22106 10237 22118
rect 10415 22106 10421 22118
rect 10231 22054 10232 22106
rect 10420 22054 10421 22106
rect 10231 22042 10237 22054
rect 10415 22042 10421 22054
rect 10231 21990 10232 22042
rect 10420 21990 10421 22042
rect 10231 21978 10237 21990
rect 10415 21978 10421 21990
rect 10231 21926 10232 21978
rect 10420 21926 10421 21978
rect 10231 21914 10237 21926
rect 10415 21914 10421 21926
rect 10231 21862 10232 21914
rect 10420 21862 10421 21914
rect 10231 21850 10237 21862
rect 10415 21850 10421 21862
rect 10231 21798 10232 21850
rect 10420 21798 10421 21850
rect 10231 21786 10237 21798
rect 10415 21786 10421 21798
rect 10231 21734 10232 21786
rect 10420 21734 10421 21786
rect 10231 21722 10237 21734
rect 10415 21722 10421 21734
rect 10231 21670 10232 21722
rect 10420 21670 10421 21722
rect 10231 21658 10237 21670
rect 10415 21658 10421 21670
rect 10231 21606 10232 21658
rect 10420 21606 10421 21658
rect 10231 21594 10237 21606
rect 10415 21594 10421 21606
rect 10231 21542 10232 21594
rect 10420 21542 10421 21594
rect 10231 21529 10237 21542
rect 10415 21529 10421 21542
rect 10231 21477 10232 21529
rect 10420 21477 10421 21529
rect 10231 21464 10237 21477
rect 10415 21464 10421 21477
rect 10231 21412 10232 21464
rect 10420 21412 10421 21464
rect 10231 21399 10237 21412
rect 10415 21399 10421 21412
rect 10231 21347 10232 21399
rect 10420 21347 10421 21399
rect 10231 21334 10237 21347
rect 10415 21334 10421 21347
rect 10231 21282 10232 21334
rect 10420 21282 10421 21334
rect 10231 21269 10237 21282
rect 10415 21269 10421 21282
rect 10231 21217 10232 21269
rect 10420 21217 10421 21269
rect 10231 21204 10237 21217
rect 10415 21204 10421 21217
rect 10231 21152 10232 21204
rect 10420 21152 10421 21204
rect 10231 21139 10237 21152
rect 10415 21139 10421 21152
rect 10231 21087 10232 21139
rect 10420 21087 10421 21139
rect 10231 21074 10237 21087
rect 10415 21074 10421 21087
rect 10231 21022 10232 21074
rect 10420 21022 10421 21074
rect 10231 21009 10237 21022
rect 10415 21009 10421 21022
rect 10231 20957 10232 21009
rect 10420 20957 10421 21009
rect 10231 20944 10237 20957
rect 10415 20944 10421 20957
rect 10231 20892 10232 20944
rect 10420 20892 10421 20944
rect 10231 20879 10237 20892
rect 10415 20879 10421 20892
rect 10231 20827 10232 20879
rect 10420 20827 10421 20879
rect 10231 20814 10237 20827
rect 10415 20814 10421 20827
rect 10231 20762 10232 20814
rect 10420 20762 10421 20814
rect 10231 19360 10237 20762
rect 10415 19360 10421 20762
rect 10231 19321 10421 19360
rect 10231 19287 10237 19321
rect 10271 19287 10309 19321
rect 10343 19287 10381 19321
rect 10415 19287 10421 19321
rect 10231 19248 10421 19287
rect 10231 19214 10237 19248
rect 10271 19214 10309 19248
rect 10343 19214 10381 19248
rect 10415 19214 10421 19248
rect 10231 19175 10421 19214
rect 10231 19141 10237 19175
rect 10271 19141 10309 19175
rect 10343 19141 10381 19175
rect 10415 19141 10421 19175
rect 10231 19102 10421 19141
rect 10231 19068 10237 19102
rect 10271 19068 10309 19102
rect 10343 19068 10381 19102
rect 10415 19068 10421 19102
rect 10231 19029 10421 19068
rect 10231 18995 10237 19029
rect 10271 18995 10309 19029
rect 10343 18995 10381 19029
rect 10415 18995 10421 19029
rect 10231 18956 10421 18995
rect 10231 18922 10237 18956
rect 10271 18922 10309 18956
rect 10343 18922 10381 18956
rect 10415 18922 10421 18956
rect 10231 18883 10421 18922
rect 10231 18849 10237 18883
rect 10271 18849 10309 18883
rect 10343 18849 10381 18883
rect 10415 18849 10421 18883
rect 10231 18810 10421 18849
rect 10231 18776 10237 18810
rect 10271 18776 10309 18810
rect 10343 18776 10381 18810
rect 10415 18776 10421 18810
rect 10231 18737 10421 18776
rect 10231 18703 10237 18737
rect 10271 18703 10309 18737
rect 10343 18703 10381 18737
rect 10415 18703 10421 18737
rect 10231 17953 10421 18703
rect 10231 17890 10237 17953
rect 10415 17890 10421 17953
rect 10231 17838 10232 17890
rect 10420 17838 10421 17890
rect 10231 17826 10237 17838
rect 10415 17826 10421 17838
rect 10231 17774 10232 17826
rect 10420 17774 10421 17826
rect 10231 17762 10237 17774
rect 10415 17762 10421 17774
rect 10231 17710 10232 17762
rect 10420 17710 10421 17762
rect 10231 17698 10237 17710
rect 10415 17698 10421 17710
rect 10231 17646 10232 17698
rect 10420 17646 10421 17698
rect 10231 17634 10237 17646
rect 10415 17634 10421 17646
rect 10231 17582 10232 17634
rect 10420 17582 10421 17634
rect 10231 17570 10237 17582
rect 10415 17570 10421 17582
rect 10231 17518 10232 17570
rect 10420 17518 10421 17570
rect 10231 17506 10237 17518
rect 10415 17506 10421 17518
rect 10231 17454 10232 17506
rect 10420 17454 10421 17506
rect 10231 17442 10237 17454
rect 10415 17442 10421 17454
rect 10231 17390 10232 17442
rect 10420 17390 10421 17442
rect 10231 17378 10237 17390
rect 10415 17378 10421 17390
rect 10231 17326 10232 17378
rect 10420 17326 10421 17378
rect 10231 17314 10237 17326
rect 10415 17314 10421 17326
rect 10231 17262 10232 17314
rect 10420 17262 10421 17314
rect 10231 17250 10237 17262
rect 10415 17250 10421 17262
rect 10231 17198 10232 17250
rect 10420 17198 10421 17250
rect 10231 17186 10237 17198
rect 10415 17186 10421 17198
rect 10231 17134 10232 17186
rect 10420 17134 10421 17186
rect 10231 17122 10237 17134
rect 10415 17122 10421 17134
rect 10231 17070 10232 17122
rect 10420 17070 10421 17122
rect 10231 17058 10237 17070
rect 10415 17058 10421 17070
rect 10231 17006 10232 17058
rect 10420 17006 10421 17058
rect 10231 16994 10237 17006
rect 10415 16994 10421 17006
rect 10231 16942 10232 16994
rect 10420 16942 10421 16994
rect 10231 16929 10237 16942
rect 10415 16929 10421 16942
rect 10231 16877 10232 16929
rect 10420 16877 10421 16929
rect 10231 16864 10237 16877
rect 10415 16864 10421 16877
rect 10231 16812 10232 16864
rect 10420 16812 10421 16864
rect 10231 16799 10237 16812
rect 10415 16799 10421 16812
rect 10231 16747 10232 16799
rect 10420 16747 10421 16799
rect 10231 16734 10237 16747
rect 10415 16734 10421 16747
rect 10231 16682 10232 16734
rect 10420 16682 10421 16734
rect 10231 16669 10237 16682
rect 10415 16669 10421 16682
rect 10231 16617 10232 16669
rect 10420 16617 10421 16669
rect 10231 16604 10237 16617
rect 10415 16604 10421 16617
rect 10231 16552 10232 16604
rect 10420 16552 10421 16604
rect 10231 16539 10237 16552
rect 10415 16539 10421 16552
rect 10231 16487 10232 16539
rect 10420 16487 10421 16539
rect 10231 16474 10237 16487
rect 10415 16474 10421 16487
rect 10231 16422 10232 16474
rect 10420 16422 10421 16474
rect 10231 16409 10237 16422
rect 10415 16409 10421 16422
rect 10231 16357 10232 16409
rect 10420 16357 10421 16409
rect 10231 16344 10237 16357
rect 10415 16344 10421 16357
rect 10231 16292 10232 16344
rect 10420 16292 10421 16344
rect 10231 16279 10237 16292
rect 10415 16279 10421 16292
rect 10231 16227 10232 16279
rect 10420 16227 10421 16279
rect 10231 16214 10237 16227
rect 10415 16214 10421 16227
rect 10231 16162 10232 16214
rect 10420 16162 10421 16214
rect 10231 14103 10237 16162
rect 10415 14103 10421 16162
rect 10231 13362 10421 14103
rect 10231 13290 10237 13362
rect 10415 13290 10421 13362
rect 10231 13238 10232 13290
rect 10420 13238 10421 13290
rect 10231 13226 10237 13238
rect 10415 13226 10421 13238
rect 10231 13174 10232 13226
rect 10420 13174 10421 13226
rect 10231 13162 10237 13174
rect 10415 13162 10421 13174
rect 10231 13110 10232 13162
rect 10420 13110 10421 13162
rect 10231 13098 10237 13110
rect 10415 13098 10421 13110
rect 10231 13046 10232 13098
rect 10420 13046 10421 13098
rect 10231 13034 10237 13046
rect 10415 13034 10421 13046
rect 10231 12982 10232 13034
rect 10420 12982 10421 13034
rect 10231 12970 10237 12982
rect 10415 12970 10421 12982
rect 10231 12918 10232 12970
rect 10420 12918 10421 12970
rect 10231 12906 10237 12918
rect 10415 12906 10421 12918
rect 10231 12854 10232 12906
rect 10420 12854 10421 12906
rect 10231 12842 10237 12854
rect 10415 12842 10421 12854
rect 10231 12790 10232 12842
rect 10420 12790 10421 12842
rect 10231 12778 10237 12790
rect 10415 12778 10421 12790
rect 10231 12726 10232 12778
rect 10420 12726 10421 12778
rect 10231 12714 10237 12726
rect 10415 12714 10421 12726
rect 10231 12662 10232 12714
rect 10420 12662 10421 12714
rect 10231 12650 10237 12662
rect 10415 12650 10421 12662
rect 10231 12598 10232 12650
rect 10420 12598 10421 12650
rect 10231 12586 10237 12598
rect 10415 12586 10421 12598
rect 10231 12534 10232 12586
rect 10420 12534 10421 12586
rect 10231 12522 10237 12534
rect 10415 12522 10421 12534
rect 10231 12470 10232 12522
rect 10420 12470 10421 12522
rect 10231 12458 10237 12470
rect 10415 12458 10421 12470
rect 10231 12406 10232 12458
rect 10420 12406 10421 12458
rect 10231 12394 10237 12406
rect 10415 12394 10421 12406
rect 10231 12342 10232 12394
rect 10420 12342 10421 12394
rect 10231 12329 10237 12342
rect 10415 12329 10421 12342
rect 10231 12277 10232 12329
rect 10420 12277 10421 12329
rect 10231 12264 10237 12277
rect 10415 12264 10421 12277
rect 10231 12212 10232 12264
rect 10420 12212 10421 12264
rect 10231 12199 10237 12212
rect 10415 12199 10421 12212
rect 10231 12147 10232 12199
rect 10420 12147 10421 12199
rect 10231 12134 10237 12147
rect 10415 12134 10421 12147
rect 10231 12082 10232 12134
rect 10420 12082 10421 12134
rect 10231 12069 10237 12082
rect 10415 12069 10421 12082
rect 10231 12017 10232 12069
rect 10420 12017 10421 12069
rect 10231 12004 10237 12017
rect 10415 12004 10421 12017
rect 10231 11952 10232 12004
rect 10420 11952 10421 12004
rect 10231 11939 10237 11952
rect 10415 11939 10421 11952
rect 10231 11887 10232 11939
rect 10420 11887 10421 11939
rect 10231 11874 10237 11887
rect 10415 11874 10421 11887
rect 10231 11822 10232 11874
rect 10420 11822 10421 11874
rect 10231 11809 10237 11822
rect 10415 11809 10421 11822
rect 10231 11757 10232 11809
rect 10420 11757 10421 11809
rect 10231 11744 10237 11757
rect 10415 11744 10421 11757
rect 10231 11692 10232 11744
rect 10420 11692 10421 11744
rect 10231 11679 10237 11692
rect 10415 11679 10421 11692
rect 10231 11627 10232 11679
rect 10420 11627 10421 11679
rect 10231 11614 10237 11627
rect 10415 11614 10421 11627
rect 10231 11562 10232 11614
rect 10420 11562 10421 11614
rect 10231 10160 10237 11562
rect 10415 10160 10421 11562
rect 10231 10121 10421 10160
rect 10231 10087 10237 10121
rect 10271 10087 10309 10121
rect 10343 10087 10381 10121
rect 10415 10087 10421 10121
rect 10231 10048 10421 10087
rect 10231 10014 10237 10048
rect 10271 10014 10309 10048
rect 10343 10014 10381 10048
rect 10415 10014 10421 10048
rect 10231 9975 10421 10014
rect 10231 9941 10237 9975
rect 10271 9941 10309 9975
rect 10343 9941 10381 9975
rect 10415 9941 10421 9975
rect 10231 9902 10421 9941
rect 10231 9868 10237 9902
rect 10271 9868 10309 9902
rect 10343 9868 10381 9902
rect 10415 9868 10421 9902
rect 10231 9829 10421 9868
rect 10231 9795 10237 9829
rect 10271 9795 10309 9829
rect 10343 9795 10381 9829
rect 10415 9795 10421 9829
rect 10231 9756 10421 9795
rect 10231 9722 10237 9756
rect 10271 9722 10309 9756
rect 10343 9722 10381 9756
rect 10415 9722 10421 9756
rect 10231 9683 10421 9722
rect 10231 9649 10237 9683
rect 10271 9649 10309 9683
rect 10343 9649 10381 9683
rect 10415 9649 10421 9683
rect 10231 9610 10421 9649
rect 10231 9576 10237 9610
rect 10271 9576 10309 9610
rect 10343 9576 10381 9610
rect 10415 9576 10421 9610
rect 10231 9537 10421 9576
rect 10231 9503 10237 9537
rect 10271 9503 10309 9537
rect 10343 9503 10381 9537
rect 10415 9503 10421 9537
rect 10231 9491 10421 9503
rect 10721 37997 10851 38003
rect 10773 37945 10799 37997
rect 10721 37929 10851 37945
rect 10773 37877 10799 37929
rect 10721 37861 10851 37877
rect 10773 37809 10799 37861
rect 10721 37793 10851 37809
rect 10773 37741 10799 37793
rect 10721 37725 10851 37741
rect 10773 37673 10799 37725
rect 10721 37657 10851 37673
rect 10773 37605 10799 37657
rect 10721 37589 10851 37605
rect 10773 37537 10799 37589
rect 10721 37521 10851 37537
rect 10773 37469 10799 37521
rect 10721 37453 10851 37469
rect 10773 37401 10799 37453
rect 10721 37385 10851 37401
rect 10773 37333 10799 37385
rect 10721 37318 10851 37333
rect 10773 37266 10799 37318
rect 10721 37251 10851 37266
rect 10773 37199 10799 37251
rect 10721 37184 10851 37199
rect 10773 37132 10799 37184
rect 10721 37117 10851 37132
rect 10773 37065 10799 37117
rect 10721 34225 10851 37065
rect 10773 34173 10799 34225
rect 10721 34161 10851 34173
rect 10773 34109 10799 34161
rect 10721 34097 10851 34109
rect 10773 34045 10799 34097
rect 10721 34033 10851 34045
rect 10773 33981 10799 34033
rect 10721 33969 10851 33981
rect 10773 33917 10799 33969
rect 10721 33905 10851 33917
rect 10773 33853 10799 33905
rect 10721 33841 10851 33853
rect 10773 33789 10799 33841
rect 10721 33777 10851 33789
rect 10773 33725 10799 33777
rect 10721 33713 10851 33725
rect 10773 33661 10799 33713
rect 10721 33649 10851 33661
rect 10773 33597 10799 33649
rect 10721 33585 10851 33597
rect 10773 33533 10799 33585
rect 10721 33521 10851 33533
rect 10773 33469 10799 33521
rect 10721 33457 10851 33469
rect 10773 33405 10799 33457
rect 10721 33393 10851 33405
rect 10773 33341 10799 33393
rect 10721 33329 10851 33341
rect 10773 33277 10799 33329
rect 10721 33264 10851 33277
rect 10773 33212 10799 33264
rect 10721 33199 10851 33212
rect 10773 33147 10799 33199
rect 10721 33134 10851 33147
rect 10773 33082 10799 33134
rect 10721 33069 10851 33082
rect 10773 33017 10799 33069
rect 10721 33004 10851 33017
rect 10773 32952 10799 33004
rect 10721 32939 10851 32952
rect 10773 32887 10799 32939
rect 10721 32874 10851 32887
rect 10773 32822 10799 32874
rect 10721 32809 10851 32822
rect 10773 32757 10799 32809
rect 10721 32744 10851 32757
rect 10773 32692 10799 32744
rect 10721 32679 10851 32692
rect 10773 32627 10799 32679
rect 10721 32614 10851 32627
rect 10773 32562 10799 32614
rect 10721 32549 10851 32562
rect 10773 32497 10799 32549
rect 10721 29625 10851 32497
rect 10773 29573 10799 29625
rect 10721 29561 10851 29573
rect 10773 29509 10799 29561
rect 10721 29497 10851 29509
rect 10773 29445 10799 29497
rect 10721 29433 10851 29445
rect 10773 29381 10799 29433
rect 10721 29369 10851 29381
rect 10773 29317 10799 29369
rect 10721 29305 10851 29317
rect 10773 29253 10799 29305
rect 10721 29241 10851 29253
rect 10773 29189 10799 29241
rect 10721 29177 10851 29189
rect 10773 29125 10799 29177
rect 10721 29113 10851 29125
rect 10773 29061 10799 29113
rect 10721 29049 10851 29061
rect 10773 28997 10799 29049
rect 10721 28985 10851 28997
rect 10773 28933 10799 28985
rect 10721 28921 10851 28933
rect 10773 28869 10799 28921
rect 10721 28857 10851 28869
rect 10773 28805 10799 28857
rect 10721 28793 10851 28805
rect 10773 28741 10799 28793
rect 10721 28729 10851 28741
rect 10773 28677 10799 28729
rect 10721 28664 10851 28677
rect 10773 28612 10799 28664
rect 10721 28599 10851 28612
rect 10773 28547 10799 28599
rect 10721 28534 10851 28547
rect 10773 28482 10799 28534
rect 10721 28469 10851 28482
rect 10773 28417 10799 28469
rect 10721 28404 10851 28417
rect 10773 28352 10799 28404
rect 10721 28339 10851 28352
rect 10773 28287 10799 28339
rect 10721 28274 10851 28287
rect 10773 28222 10799 28274
rect 10721 28209 10851 28222
rect 10773 28157 10799 28209
rect 10721 28144 10851 28157
rect 10773 28092 10799 28144
rect 10721 28079 10851 28092
rect 10773 28027 10799 28079
rect 10721 28014 10851 28027
rect 10773 27962 10799 28014
rect 10721 27949 10851 27962
rect 10773 27897 10799 27949
rect 10721 25025 10851 27897
rect 10773 24973 10799 25025
rect 10721 24961 10851 24973
rect 10773 24909 10799 24961
rect 10721 24897 10851 24909
rect 10773 24845 10799 24897
rect 10721 24833 10851 24845
rect 10773 24781 10799 24833
rect 10721 24769 10851 24781
rect 10773 24717 10799 24769
rect 10721 24705 10851 24717
rect 10773 24653 10799 24705
rect 10721 24641 10851 24653
rect 10773 24589 10799 24641
rect 10721 24577 10851 24589
rect 10773 24525 10799 24577
rect 10721 24513 10851 24525
rect 10773 24461 10799 24513
rect 10721 24449 10851 24461
rect 10773 24397 10799 24449
rect 10721 24385 10851 24397
rect 10773 24333 10799 24385
rect 10721 24321 10851 24333
rect 10773 24269 10799 24321
rect 10721 24257 10851 24269
rect 10773 24205 10799 24257
rect 10721 24193 10851 24205
rect 10773 24141 10799 24193
rect 10721 24129 10851 24141
rect 10773 24077 10799 24129
rect 10721 24064 10851 24077
rect 10773 24012 10799 24064
rect 10721 23999 10851 24012
rect 10773 23947 10799 23999
rect 10721 23934 10851 23947
rect 10773 23882 10799 23934
rect 10721 23869 10851 23882
rect 10773 23817 10799 23869
rect 10721 23804 10851 23817
rect 10773 23752 10799 23804
rect 10721 23739 10851 23752
rect 10773 23687 10799 23739
rect 10721 23674 10851 23687
rect 10773 23622 10799 23674
rect 10721 23609 10851 23622
rect 10773 23557 10799 23609
rect 10721 23544 10851 23557
rect 10773 23492 10799 23544
rect 10721 23479 10851 23492
rect 10773 23427 10799 23479
rect 10721 23414 10851 23427
rect 10773 23362 10799 23414
rect 10721 23349 10851 23362
rect 10773 23297 10799 23349
rect 10721 20425 10851 23297
rect 10773 20373 10799 20425
rect 10721 20361 10851 20373
rect 10773 20309 10799 20361
rect 10721 20297 10851 20309
rect 10773 20245 10799 20297
rect 10721 20233 10851 20245
rect 10773 20181 10799 20233
rect 10721 20169 10851 20181
rect 10773 20117 10799 20169
rect 10721 20105 10851 20117
rect 10773 20053 10799 20105
rect 10721 20041 10851 20053
rect 10773 19989 10799 20041
rect 10721 19977 10851 19989
rect 10773 19925 10799 19977
rect 10721 19913 10851 19925
rect 10773 19861 10799 19913
rect 10721 19849 10851 19861
rect 10773 19797 10799 19849
rect 10721 19785 10851 19797
rect 10773 19733 10799 19785
rect 10721 19721 10851 19733
rect 10773 19669 10799 19721
rect 10721 19657 10851 19669
rect 10773 19605 10799 19657
rect 10721 19593 10851 19605
rect 10773 19541 10799 19593
rect 10721 19529 10851 19541
rect 10773 19477 10799 19529
rect 10721 19464 10851 19477
rect 10773 19412 10799 19464
rect 10721 19399 10851 19412
rect 10773 19347 10799 19399
rect 10721 19334 10851 19347
rect 10773 19282 10799 19334
rect 10721 19269 10851 19282
rect 10773 19217 10799 19269
rect 10721 19204 10851 19217
rect 10773 19152 10799 19204
rect 10721 19139 10851 19152
rect 10773 19087 10799 19139
rect 10721 19074 10851 19087
rect 10773 19022 10799 19074
rect 10721 19009 10851 19022
rect 10773 18957 10799 19009
rect 10721 18944 10851 18957
rect 10773 18892 10799 18944
rect 10721 18879 10851 18892
rect 10773 18827 10799 18879
rect 10721 18814 10851 18827
rect 10773 18762 10799 18814
rect 10721 18749 10851 18762
rect 10773 18697 10799 18749
rect 10721 15825 10851 18697
rect 10773 15773 10799 15825
rect 10721 15761 10851 15773
rect 10773 15709 10799 15761
rect 10721 15697 10851 15709
rect 10773 15645 10799 15697
rect 10721 15633 10851 15645
rect 10773 15581 10799 15633
rect 10721 15569 10851 15581
rect 10773 15517 10799 15569
rect 10721 15505 10851 15517
rect 10773 15453 10799 15505
rect 10721 15441 10851 15453
rect 10773 15389 10799 15441
rect 10721 15377 10851 15389
rect 10773 15325 10799 15377
rect 10721 15313 10851 15325
rect 10773 15261 10799 15313
rect 10721 15249 10851 15261
rect 10773 15197 10799 15249
rect 10721 15185 10851 15197
rect 10773 15133 10799 15185
rect 10721 15121 10851 15133
rect 10773 15069 10799 15121
rect 10721 15057 10851 15069
rect 10773 15005 10799 15057
rect 10721 14993 10851 15005
rect 10773 14941 10799 14993
rect 10721 14929 10851 14941
rect 10773 14877 10799 14929
rect 10721 14864 10851 14877
rect 10773 14812 10799 14864
rect 10721 14799 10851 14812
rect 10773 14747 10799 14799
rect 10721 14734 10851 14747
rect 10773 14682 10799 14734
rect 10721 14669 10851 14682
rect 10773 14617 10799 14669
rect 10721 14604 10851 14617
rect 10773 14552 10799 14604
rect 10721 14539 10851 14552
rect 10773 14487 10799 14539
rect 10721 14474 10851 14487
rect 10773 14422 10799 14474
rect 10721 14409 10851 14422
rect 10773 14357 10799 14409
rect 10721 14344 10851 14357
rect 10773 14292 10799 14344
rect 10721 14279 10851 14292
rect 10773 14227 10799 14279
rect 10721 14214 10851 14227
rect 10773 14162 10799 14214
rect 10721 14149 10851 14162
rect 10773 14097 10799 14149
rect 10721 11225 10851 14097
rect 10773 11173 10799 11225
rect 10721 11161 10851 11173
rect 10773 11109 10799 11161
rect 10721 11097 10851 11109
rect 10773 11045 10799 11097
rect 10721 11033 10851 11045
rect 10773 10981 10799 11033
rect 10721 10969 10851 10981
rect 10773 10917 10799 10969
rect 10721 10905 10851 10917
rect 10773 10853 10799 10905
rect 10721 10841 10851 10853
rect 10773 10789 10799 10841
rect 10721 10777 10851 10789
rect 10773 10725 10799 10777
rect 10721 10713 10851 10725
rect 10773 10661 10799 10713
rect 10721 10649 10851 10661
rect 10773 10597 10799 10649
rect 10721 10585 10851 10597
rect 10773 10533 10799 10585
rect 10721 10521 10851 10533
rect 10773 10469 10799 10521
rect 10721 10457 10851 10469
rect 10773 10405 10799 10457
rect 10721 10393 10851 10405
rect 10773 10341 10799 10393
rect 10721 10329 10851 10341
rect 10773 10277 10799 10329
rect 10721 10264 10851 10277
rect 10773 10212 10799 10264
rect 10721 10199 10851 10212
rect 10773 10147 10799 10199
rect 10721 10134 10851 10147
rect 10773 10082 10799 10134
rect 10721 10069 10851 10082
rect 10773 10017 10799 10069
rect 10721 10004 10851 10017
rect 10773 9952 10799 10004
rect 10721 9939 10851 9952
rect 10773 9887 10799 9939
rect 10721 9874 10851 9887
rect 10773 9822 10799 9874
rect 10721 9809 10851 9822
rect 10773 9757 10799 9809
rect 10721 9744 10851 9757
rect 10773 9692 10799 9744
rect 10721 9679 10851 9692
rect 10773 9627 10799 9679
rect 10721 9614 10851 9627
rect 10773 9562 10799 9614
rect 10721 9549 10851 9562
rect 10773 9497 10799 9549
rect 10721 9491 10851 9497
rect 11151 37979 11157 38013
rect 11191 37979 11229 38013
rect 11263 37979 11301 38013
rect 11335 37979 11341 38013
rect 12071 39028 12261 39040
rect 12071 39009 12077 39028
rect 12255 39009 12261 39028
rect 12071 38957 12072 39009
rect 12260 38957 12261 39009
rect 12071 38944 12077 38957
rect 12255 38944 12261 38957
rect 12071 38892 12072 38944
rect 12260 38892 12261 38944
rect 12071 38879 12077 38892
rect 12255 38879 12261 38892
rect 12071 38827 12072 38879
rect 12260 38827 12261 38879
rect 12071 38814 12077 38827
rect 12255 38814 12261 38827
rect 12071 38762 12072 38814
rect 12260 38762 12261 38814
rect 12071 38749 12077 38762
rect 12255 38749 12261 38762
rect 12071 38697 12072 38749
rect 12260 38697 12261 38749
rect 12071 38684 12077 38697
rect 12255 38684 12261 38697
rect 12071 38632 12072 38684
rect 12260 38632 12261 38684
rect 12071 38619 12077 38632
rect 12255 38619 12261 38632
rect 12071 38567 12072 38619
rect 12260 38567 12261 38619
rect 12071 38554 12077 38567
rect 12255 38554 12261 38567
rect 12071 38502 12072 38554
rect 12260 38502 12261 38554
rect 12071 38490 12077 38502
rect 12255 38490 12261 38502
rect 12071 38438 12072 38490
rect 12124 38438 12140 38490
rect 12192 38438 12208 38490
rect 12260 38438 12261 38490
rect 12071 38426 12077 38438
rect 12111 38426 12149 38438
rect 12183 38426 12221 38438
rect 12255 38426 12261 38438
rect 12071 38374 12072 38426
rect 12124 38374 12140 38426
rect 12192 38374 12208 38426
rect 12260 38374 12261 38426
rect 12071 38362 12077 38374
rect 12111 38362 12149 38374
rect 12183 38362 12221 38374
rect 12255 38362 12261 38374
rect 12071 38310 12072 38362
rect 12124 38310 12140 38362
rect 12192 38310 12208 38362
rect 12260 38310 12261 38362
rect 12071 38305 12261 38310
rect 12071 38298 12077 38305
rect 12111 38298 12149 38305
rect 12183 38298 12221 38305
rect 12255 38298 12261 38305
rect 12071 38246 12072 38298
rect 12124 38246 12140 38298
rect 12192 38246 12208 38298
rect 12260 38246 12261 38298
rect 12071 38234 12261 38246
rect 12071 38182 12072 38234
rect 12124 38182 12140 38234
rect 12192 38182 12208 38234
rect 12260 38182 12261 38234
rect 12071 38170 12261 38182
rect 12071 38118 12072 38170
rect 12124 38118 12140 38170
rect 12192 38118 12208 38170
rect 12260 38118 12261 38170
rect 12071 38086 12261 38118
rect 12071 38052 12077 38086
rect 12111 38052 12149 38086
rect 12183 38052 12221 38086
rect 12255 38052 12261 38086
rect 12071 38013 12261 38052
rect 11151 37940 11341 37979
rect 11151 37906 11157 37940
rect 11191 37906 11229 37940
rect 11263 37906 11301 37940
rect 11335 37906 11341 37940
rect 11151 37867 11341 37906
rect 11151 37833 11157 37867
rect 11191 37833 11229 37867
rect 11263 37833 11301 37867
rect 11335 37833 11341 37867
rect 11151 37794 11341 37833
rect 11151 37760 11157 37794
rect 11191 37760 11229 37794
rect 11263 37760 11301 37794
rect 11335 37760 11341 37794
rect 11151 37721 11341 37760
rect 11151 37687 11157 37721
rect 11191 37687 11229 37721
rect 11263 37687 11301 37721
rect 11335 37687 11341 37721
rect 11151 37648 11341 37687
rect 11151 37614 11157 37648
rect 11191 37614 11229 37648
rect 11263 37614 11301 37648
rect 11335 37614 11341 37648
rect 11151 37575 11341 37614
rect 11151 37541 11157 37575
rect 11191 37541 11229 37575
rect 11263 37541 11301 37575
rect 11335 37541 11341 37575
rect 11151 37502 11341 37541
rect 11151 37468 11157 37502
rect 11191 37468 11229 37502
rect 11263 37468 11301 37502
rect 11335 37468 11341 37502
rect 11151 37429 11341 37468
rect 11151 37395 11157 37429
rect 11191 37395 11229 37429
rect 11263 37395 11301 37429
rect 11335 37395 11341 37429
rect 11151 37356 11341 37395
rect 11151 37322 11157 37356
rect 11191 37322 11229 37356
rect 11263 37322 11301 37356
rect 11335 37322 11341 37356
rect 11151 37283 11341 37322
rect 11151 37249 11157 37283
rect 11191 37249 11229 37283
rect 11263 37249 11301 37283
rect 11335 37249 11341 37283
rect 11151 37210 11341 37249
rect 11151 37176 11157 37210
rect 11191 37176 11229 37210
rect 11263 37176 11301 37210
rect 11335 37176 11341 37210
rect 11151 37137 11341 37176
rect 11151 37103 11157 37137
rect 11191 37103 11229 37137
rect 11263 37103 11301 37137
rect 11335 37103 11341 37137
rect 11151 36353 11341 37103
rect 11151 36290 11157 36353
rect 11335 36290 11341 36353
rect 11151 36238 11152 36290
rect 11340 36238 11341 36290
rect 11151 36226 11157 36238
rect 11335 36226 11341 36238
rect 11151 36174 11152 36226
rect 11340 36174 11341 36226
rect 11151 36162 11157 36174
rect 11335 36162 11341 36174
rect 11151 36110 11152 36162
rect 11340 36110 11341 36162
rect 11151 36098 11157 36110
rect 11335 36098 11341 36110
rect 11151 36046 11152 36098
rect 11340 36046 11341 36098
rect 11151 36034 11157 36046
rect 11335 36034 11341 36046
rect 11151 35982 11152 36034
rect 11340 35982 11341 36034
rect 11151 35970 11157 35982
rect 11335 35970 11341 35982
rect 11151 35918 11152 35970
rect 11340 35918 11341 35970
rect 11151 35906 11157 35918
rect 11335 35906 11341 35918
rect 11151 35854 11152 35906
rect 11340 35854 11341 35906
rect 11151 35842 11157 35854
rect 11335 35842 11341 35854
rect 11151 35790 11152 35842
rect 11340 35790 11341 35842
rect 11151 35778 11157 35790
rect 11335 35778 11341 35790
rect 11151 35726 11152 35778
rect 11340 35726 11341 35778
rect 11151 35714 11157 35726
rect 11335 35714 11341 35726
rect 11151 35662 11152 35714
rect 11340 35662 11341 35714
rect 11151 35650 11157 35662
rect 11335 35650 11341 35662
rect 11151 35598 11152 35650
rect 11340 35598 11341 35650
rect 11151 35586 11157 35598
rect 11335 35586 11341 35598
rect 11151 35534 11152 35586
rect 11340 35534 11341 35586
rect 11151 35522 11157 35534
rect 11335 35522 11341 35534
rect 11151 35470 11152 35522
rect 11340 35470 11341 35522
rect 11151 35458 11157 35470
rect 11335 35458 11341 35470
rect 11151 35406 11152 35458
rect 11340 35406 11341 35458
rect 11151 35394 11157 35406
rect 11335 35394 11341 35406
rect 11151 35342 11152 35394
rect 11340 35342 11341 35394
rect 11151 35329 11157 35342
rect 11335 35329 11341 35342
rect 11151 35277 11152 35329
rect 11340 35277 11341 35329
rect 11151 35264 11157 35277
rect 11335 35264 11341 35277
rect 11151 35212 11152 35264
rect 11340 35212 11341 35264
rect 11151 35199 11157 35212
rect 11335 35199 11341 35212
rect 11151 35147 11152 35199
rect 11340 35147 11341 35199
rect 11151 35134 11157 35147
rect 11335 35134 11341 35147
rect 11151 35082 11152 35134
rect 11340 35082 11341 35134
rect 11151 35069 11157 35082
rect 11335 35069 11341 35082
rect 11151 35017 11152 35069
rect 11340 35017 11341 35069
rect 11151 35004 11157 35017
rect 11335 35004 11341 35017
rect 11151 34952 11152 35004
rect 11340 34952 11341 35004
rect 11151 34939 11157 34952
rect 11335 34939 11341 34952
rect 11151 34887 11152 34939
rect 11340 34887 11341 34939
rect 11151 34874 11157 34887
rect 11335 34874 11341 34887
rect 11151 34822 11152 34874
rect 11340 34822 11341 34874
rect 11151 34809 11157 34822
rect 11335 34809 11341 34822
rect 11151 34757 11152 34809
rect 11340 34757 11341 34809
rect 11151 34744 11157 34757
rect 11335 34744 11341 34757
rect 11151 34692 11152 34744
rect 11340 34692 11341 34744
rect 11151 34679 11157 34692
rect 11335 34679 11341 34692
rect 11151 34627 11152 34679
rect 11340 34627 11341 34679
rect 11151 34614 11157 34627
rect 11335 34614 11341 34627
rect 11151 34562 11152 34614
rect 11340 34562 11341 34614
rect 11151 32503 11157 34562
rect 11335 32503 11341 34562
rect 11151 31753 11341 32503
rect 11151 31690 11157 31753
rect 11335 31690 11341 31753
rect 11151 31638 11152 31690
rect 11340 31638 11341 31690
rect 11151 31626 11157 31638
rect 11335 31626 11341 31638
rect 11151 31574 11152 31626
rect 11340 31574 11341 31626
rect 11151 31562 11157 31574
rect 11335 31562 11341 31574
rect 11151 31510 11152 31562
rect 11340 31510 11341 31562
rect 11151 31498 11157 31510
rect 11335 31498 11341 31510
rect 11151 31446 11152 31498
rect 11340 31446 11341 31498
rect 11151 31434 11157 31446
rect 11335 31434 11341 31446
rect 11151 31382 11152 31434
rect 11340 31382 11341 31434
rect 11151 31370 11157 31382
rect 11335 31370 11341 31382
rect 11151 31318 11152 31370
rect 11340 31318 11341 31370
rect 11151 31306 11157 31318
rect 11335 31306 11341 31318
rect 11151 31254 11152 31306
rect 11340 31254 11341 31306
rect 11151 31242 11157 31254
rect 11335 31242 11341 31254
rect 11151 31190 11152 31242
rect 11340 31190 11341 31242
rect 11151 31178 11157 31190
rect 11335 31178 11341 31190
rect 11151 31126 11152 31178
rect 11340 31126 11341 31178
rect 11151 31114 11157 31126
rect 11335 31114 11341 31126
rect 11151 31062 11152 31114
rect 11340 31062 11341 31114
rect 11151 31050 11157 31062
rect 11335 31050 11341 31062
rect 11151 30998 11152 31050
rect 11340 30998 11341 31050
rect 11151 30986 11157 30998
rect 11335 30986 11341 30998
rect 11151 30934 11152 30986
rect 11340 30934 11341 30986
rect 11151 30922 11157 30934
rect 11335 30922 11341 30934
rect 11151 30870 11152 30922
rect 11340 30870 11341 30922
rect 11151 30858 11157 30870
rect 11335 30858 11341 30870
rect 11151 30806 11152 30858
rect 11340 30806 11341 30858
rect 11151 30794 11157 30806
rect 11335 30794 11341 30806
rect 11151 30742 11152 30794
rect 11340 30742 11341 30794
rect 11151 30729 11157 30742
rect 11335 30729 11341 30742
rect 11151 30677 11152 30729
rect 11340 30677 11341 30729
rect 11151 30664 11157 30677
rect 11335 30664 11341 30677
rect 11151 30612 11152 30664
rect 11340 30612 11341 30664
rect 11151 30599 11157 30612
rect 11335 30599 11341 30612
rect 11151 30547 11152 30599
rect 11340 30547 11341 30599
rect 11151 30534 11157 30547
rect 11335 30534 11341 30547
rect 11151 30482 11152 30534
rect 11340 30482 11341 30534
rect 11151 30469 11157 30482
rect 11335 30469 11341 30482
rect 11151 30417 11152 30469
rect 11340 30417 11341 30469
rect 11151 30404 11157 30417
rect 11335 30404 11341 30417
rect 11151 30352 11152 30404
rect 11340 30352 11341 30404
rect 11151 30339 11157 30352
rect 11335 30339 11341 30352
rect 11151 30287 11152 30339
rect 11340 30287 11341 30339
rect 11151 30274 11157 30287
rect 11335 30274 11341 30287
rect 11151 30222 11152 30274
rect 11340 30222 11341 30274
rect 11151 30209 11157 30222
rect 11335 30209 11341 30222
rect 11151 30157 11152 30209
rect 11340 30157 11341 30209
rect 11151 30144 11157 30157
rect 11335 30144 11341 30157
rect 11151 30092 11152 30144
rect 11340 30092 11341 30144
rect 11151 30079 11157 30092
rect 11335 30079 11341 30092
rect 11151 30027 11152 30079
rect 11340 30027 11341 30079
rect 11151 30014 11157 30027
rect 11335 30014 11341 30027
rect 11151 29962 11152 30014
rect 11340 29962 11341 30014
rect 11151 27903 11157 29962
rect 11335 27903 11341 29962
rect 11151 27153 11341 27903
rect 11151 27090 11157 27153
rect 11335 27090 11341 27153
rect 11151 27038 11152 27090
rect 11340 27038 11341 27090
rect 11151 27026 11157 27038
rect 11335 27026 11341 27038
rect 11151 26974 11152 27026
rect 11340 26974 11341 27026
rect 11151 26962 11157 26974
rect 11335 26962 11341 26974
rect 11151 26910 11152 26962
rect 11340 26910 11341 26962
rect 11151 26898 11157 26910
rect 11335 26898 11341 26910
rect 11151 26846 11152 26898
rect 11340 26846 11341 26898
rect 11151 26834 11157 26846
rect 11335 26834 11341 26846
rect 11151 26782 11152 26834
rect 11340 26782 11341 26834
rect 11151 26770 11157 26782
rect 11335 26770 11341 26782
rect 11151 26718 11152 26770
rect 11340 26718 11341 26770
rect 11151 26706 11157 26718
rect 11335 26706 11341 26718
rect 11151 26654 11152 26706
rect 11340 26654 11341 26706
rect 11151 26642 11157 26654
rect 11335 26642 11341 26654
rect 11151 26590 11152 26642
rect 11340 26590 11341 26642
rect 11151 26578 11157 26590
rect 11335 26578 11341 26590
rect 11151 26526 11152 26578
rect 11340 26526 11341 26578
rect 11151 26514 11157 26526
rect 11335 26514 11341 26526
rect 11151 26462 11152 26514
rect 11340 26462 11341 26514
rect 11151 26450 11157 26462
rect 11335 26450 11341 26462
rect 11151 26398 11152 26450
rect 11340 26398 11341 26450
rect 11151 26386 11157 26398
rect 11335 26386 11341 26398
rect 11151 26334 11152 26386
rect 11340 26334 11341 26386
rect 11151 26322 11157 26334
rect 11335 26322 11341 26334
rect 11151 26270 11152 26322
rect 11340 26270 11341 26322
rect 11151 26258 11157 26270
rect 11335 26258 11341 26270
rect 11151 26206 11152 26258
rect 11340 26206 11341 26258
rect 11151 26194 11157 26206
rect 11335 26194 11341 26206
rect 11151 26142 11152 26194
rect 11340 26142 11341 26194
rect 11151 26129 11157 26142
rect 11335 26129 11341 26142
rect 11151 26077 11152 26129
rect 11340 26077 11341 26129
rect 11151 26064 11157 26077
rect 11335 26064 11341 26077
rect 11151 26012 11152 26064
rect 11340 26012 11341 26064
rect 11151 25999 11157 26012
rect 11335 25999 11341 26012
rect 11151 25947 11152 25999
rect 11340 25947 11341 25999
rect 11151 25934 11157 25947
rect 11335 25934 11341 25947
rect 11151 25882 11152 25934
rect 11340 25882 11341 25934
rect 11151 25869 11157 25882
rect 11335 25869 11341 25882
rect 11151 25817 11152 25869
rect 11340 25817 11341 25869
rect 11151 25804 11157 25817
rect 11335 25804 11341 25817
rect 11151 25752 11152 25804
rect 11340 25752 11341 25804
rect 11151 25739 11157 25752
rect 11335 25739 11341 25752
rect 11151 25687 11152 25739
rect 11340 25687 11341 25739
rect 11151 25674 11157 25687
rect 11335 25674 11341 25687
rect 11151 25622 11152 25674
rect 11340 25622 11341 25674
rect 11151 25609 11157 25622
rect 11335 25609 11341 25622
rect 11151 25557 11152 25609
rect 11340 25557 11341 25609
rect 11151 25544 11157 25557
rect 11335 25544 11341 25557
rect 11151 25492 11152 25544
rect 11340 25492 11341 25544
rect 11151 25479 11157 25492
rect 11335 25479 11341 25492
rect 11151 25427 11152 25479
rect 11340 25427 11341 25479
rect 11151 25414 11157 25427
rect 11335 25414 11341 25427
rect 11151 25362 11152 25414
rect 11340 25362 11341 25414
rect 11151 23303 11157 25362
rect 11335 23303 11341 25362
rect 11151 22562 11341 23303
rect 11151 22490 11157 22562
rect 11335 22490 11341 22562
rect 11151 22438 11152 22490
rect 11340 22438 11341 22490
rect 11151 22426 11157 22438
rect 11335 22426 11341 22438
rect 11151 22374 11152 22426
rect 11340 22374 11341 22426
rect 11151 22362 11157 22374
rect 11335 22362 11341 22374
rect 11151 22310 11152 22362
rect 11340 22310 11341 22362
rect 11151 22298 11157 22310
rect 11335 22298 11341 22310
rect 11151 22246 11152 22298
rect 11340 22246 11341 22298
rect 11151 22234 11157 22246
rect 11335 22234 11341 22246
rect 11151 22182 11152 22234
rect 11340 22182 11341 22234
rect 11151 22170 11157 22182
rect 11335 22170 11341 22182
rect 11151 22118 11152 22170
rect 11340 22118 11341 22170
rect 11151 22106 11157 22118
rect 11335 22106 11341 22118
rect 11151 22054 11152 22106
rect 11340 22054 11341 22106
rect 11151 22042 11157 22054
rect 11335 22042 11341 22054
rect 11151 21990 11152 22042
rect 11340 21990 11341 22042
rect 11151 21978 11157 21990
rect 11335 21978 11341 21990
rect 11151 21926 11152 21978
rect 11340 21926 11341 21978
rect 11151 21914 11157 21926
rect 11335 21914 11341 21926
rect 11151 21862 11152 21914
rect 11340 21862 11341 21914
rect 11151 21850 11157 21862
rect 11335 21850 11341 21862
rect 11151 21798 11152 21850
rect 11340 21798 11341 21850
rect 11151 21786 11157 21798
rect 11335 21786 11341 21798
rect 11151 21734 11152 21786
rect 11340 21734 11341 21786
rect 11151 21722 11157 21734
rect 11335 21722 11341 21734
rect 11151 21670 11152 21722
rect 11340 21670 11341 21722
rect 11151 21658 11157 21670
rect 11335 21658 11341 21670
rect 11151 21606 11152 21658
rect 11340 21606 11341 21658
rect 11151 21594 11157 21606
rect 11335 21594 11341 21606
rect 11151 21542 11152 21594
rect 11340 21542 11341 21594
rect 11151 21529 11157 21542
rect 11335 21529 11341 21542
rect 11151 21477 11152 21529
rect 11340 21477 11341 21529
rect 11151 21464 11157 21477
rect 11335 21464 11341 21477
rect 11151 21412 11152 21464
rect 11340 21412 11341 21464
rect 11151 21399 11157 21412
rect 11335 21399 11341 21412
rect 11151 21347 11152 21399
rect 11340 21347 11341 21399
rect 11151 21334 11157 21347
rect 11335 21334 11341 21347
rect 11151 21282 11152 21334
rect 11340 21282 11341 21334
rect 11151 21269 11157 21282
rect 11335 21269 11341 21282
rect 11151 21217 11152 21269
rect 11340 21217 11341 21269
rect 11151 21204 11157 21217
rect 11335 21204 11341 21217
rect 11151 21152 11152 21204
rect 11340 21152 11341 21204
rect 11151 21139 11157 21152
rect 11335 21139 11341 21152
rect 11151 21087 11152 21139
rect 11340 21087 11341 21139
rect 11151 21074 11157 21087
rect 11335 21074 11341 21087
rect 11151 21022 11152 21074
rect 11340 21022 11341 21074
rect 11151 21009 11157 21022
rect 11335 21009 11341 21022
rect 11151 20957 11152 21009
rect 11340 20957 11341 21009
rect 11151 20944 11157 20957
rect 11335 20944 11341 20957
rect 11151 20892 11152 20944
rect 11340 20892 11341 20944
rect 11151 20879 11157 20892
rect 11335 20879 11341 20892
rect 11151 20827 11152 20879
rect 11340 20827 11341 20879
rect 11151 20814 11157 20827
rect 11335 20814 11341 20827
rect 11151 20762 11152 20814
rect 11340 20762 11341 20814
rect 11151 19360 11157 20762
rect 11335 19360 11341 20762
rect 11151 19321 11341 19360
rect 11151 19287 11157 19321
rect 11191 19287 11229 19321
rect 11263 19287 11301 19321
rect 11335 19287 11341 19321
rect 11151 19248 11341 19287
rect 11151 19214 11157 19248
rect 11191 19214 11229 19248
rect 11263 19214 11301 19248
rect 11335 19214 11341 19248
rect 11151 19175 11341 19214
rect 11151 19141 11157 19175
rect 11191 19141 11229 19175
rect 11263 19141 11301 19175
rect 11335 19141 11341 19175
rect 11151 19102 11341 19141
rect 11151 19068 11157 19102
rect 11191 19068 11229 19102
rect 11263 19068 11301 19102
rect 11335 19068 11341 19102
rect 11151 19029 11341 19068
rect 11151 18995 11157 19029
rect 11191 18995 11229 19029
rect 11263 18995 11301 19029
rect 11335 18995 11341 19029
rect 11151 18956 11341 18995
rect 11151 18922 11157 18956
rect 11191 18922 11229 18956
rect 11263 18922 11301 18956
rect 11335 18922 11341 18956
rect 11151 18883 11341 18922
rect 11151 18849 11157 18883
rect 11191 18849 11229 18883
rect 11263 18849 11301 18883
rect 11335 18849 11341 18883
rect 11151 18810 11341 18849
rect 11151 18776 11157 18810
rect 11191 18776 11229 18810
rect 11263 18776 11301 18810
rect 11335 18776 11341 18810
rect 11151 18737 11341 18776
rect 11151 18703 11157 18737
rect 11191 18703 11229 18737
rect 11263 18703 11301 18737
rect 11335 18703 11341 18737
rect 11151 17953 11341 18703
rect 11151 17890 11157 17953
rect 11335 17890 11341 17953
rect 11151 17838 11152 17890
rect 11340 17838 11341 17890
rect 11151 17826 11157 17838
rect 11335 17826 11341 17838
rect 11151 17774 11152 17826
rect 11340 17774 11341 17826
rect 11151 17762 11157 17774
rect 11335 17762 11341 17774
rect 11151 17710 11152 17762
rect 11340 17710 11341 17762
rect 11151 17698 11157 17710
rect 11335 17698 11341 17710
rect 11151 17646 11152 17698
rect 11340 17646 11341 17698
rect 11151 17634 11157 17646
rect 11335 17634 11341 17646
rect 11151 17582 11152 17634
rect 11340 17582 11341 17634
rect 11151 17570 11157 17582
rect 11335 17570 11341 17582
rect 11151 17518 11152 17570
rect 11340 17518 11341 17570
rect 11151 17506 11157 17518
rect 11335 17506 11341 17518
rect 11151 17454 11152 17506
rect 11340 17454 11341 17506
rect 11151 17442 11157 17454
rect 11335 17442 11341 17454
rect 11151 17390 11152 17442
rect 11340 17390 11341 17442
rect 11151 17378 11157 17390
rect 11335 17378 11341 17390
rect 11151 17326 11152 17378
rect 11340 17326 11341 17378
rect 11151 17314 11157 17326
rect 11335 17314 11341 17326
rect 11151 17262 11152 17314
rect 11340 17262 11341 17314
rect 11151 17250 11157 17262
rect 11335 17250 11341 17262
rect 11151 17198 11152 17250
rect 11340 17198 11341 17250
rect 11151 17186 11157 17198
rect 11335 17186 11341 17198
rect 11151 17134 11152 17186
rect 11340 17134 11341 17186
rect 11151 17122 11157 17134
rect 11335 17122 11341 17134
rect 11151 17070 11152 17122
rect 11340 17070 11341 17122
rect 11151 17058 11157 17070
rect 11335 17058 11341 17070
rect 11151 17006 11152 17058
rect 11340 17006 11341 17058
rect 11151 16994 11157 17006
rect 11335 16994 11341 17006
rect 11151 16942 11152 16994
rect 11340 16942 11341 16994
rect 11151 16929 11157 16942
rect 11335 16929 11341 16942
rect 11151 16877 11152 16929
rect 11340 16877 11341 16929
rect 11151 16864 11157 16877
rect 11335 16864 11341 16877
rect 11151 16812 11152 16864
rect 11340 16812 11341 16864
rect 11151 16799 11157 16812
rect 11335 16799 11341 16812
rect 11151 16747 11152 16799
rect 11340 16747 11341 16799
rect 11151 16734 11157 16747
rect 11335 16734 11341 16747
rect 11151 16682 11152 16734
rect 11340 16682 11341 16734
rect 11151 16669 11157 16682
rect 11335 16669 11341 16682
rect 11151 16617 11152 16669
rect 11340 16617 11341 16669
rect 11151 16604 11157 16617
rect 11335 16604 11341 16617
rect 11151 16552 11152 16604
rect 11340 16552 11341 16604
rect 11151 16539 11157 16552
rect 11335 16539 11341 16552
rect 11151 16487 11152 16539
rect 11340 16487 11341 16539
rect 11151 16474 11157 16487
rect 11335 16474 11341 16487
rect 11151 16422 11152 16474
rect 11340 16422 11341 16474
rect 11151 16409 11157 16422
rect 11335 16409 11341 16422
rect 11151 16357 11152 16409
rect 11340 16357 11341 16409
rect 11151 16344 11157 16357
rect 11335 16344 11341 16357
rect 11151 16292 11152 16344
rect 11340 16292 11341 16344
rect 11151 16279 11157 16292
rect 11335 16279 11341 16292
rect 11151 16227 11152 16279
rect 11340 16227 11341 16279
rect 11151 16214 11157 16227
rect 11335 16214 11341 16227
rect 11151 16162 11152 16214
rect 11340 16162 11341 16214
rect 11151 14103 11157 16162
rect 11335 14103 11341 16162
rect 11151 13362 11341 14103
rect 11151 13290 11157 13362
rect 11335 13290 11341 13362
rect 11151 13238 11152 13290
rect 11340 13238 11341 13290
rect 11151 13226 11157 13238
rect 11335 13226 11341 13238
rect 11151 13174 11152 13226
rect 11340 13174 11341 13226
rect 11151 13162 11157 13174
rect 11335 13162 11341 13174
rect 11151 13110 11152 13162
rect 11340 13110 11341 13162
rect 11151 13098 11157 13110
rect 11335 13098 11341 13110
rect 11151 13046 11152 13098
rect 11340 13046 11341 13098
rect 11151 13034 11157 13046
rect 11335 13034 11341 13046
rect 11151 12982 11152 13034
rect 11340 12982 11341 13034
rect 11151 12970 11157 12982
rect 11335 12970 11341 12982
rect 11151 12918 11152 12970
rect 11340 12918 11341 12970
rect 11151 12906 11157 12918
rect 11335 12906 11341 12918
rect 11151 12854 11152 12906
rect 11340 12854 11341 12906
rect 11151 12842 11157 12854
rect 11335 12842 11341 12854
rect 11151 12790 11152 12842
rect 11340 12790 11341 12842
rect 11151 12778 11157 12790
rect 11335 12778 11341 12790
rect 11151 12726 11152 12778
rect 11340 12726 11341 12778
rect 11151 12714 11157 12726
rect 11335 12714 11341 12726
rect 11151 12662 11152 12714
rect 11340 12662 11341 12714
rect 11151 12650 11157 12662
rect 11335 12650 11341 12662
rect 11151 12598 11152 12650
rect 11340 12598 11341 12650
rect 11151 12586 11157 12598
rect 11335 12586 11341 12598
rect 11151 12534 11152 12586
rect 11340 12534 11341 12586
rect 11151 12522 11157 12534
rect 11335 12522 11341 12534
rect 11151 12470 11152 12522
rect 11340 12470 11341 12522
rect 11151 12458 11157 12470
rect 11335 12458 11341 12470
rect 11151 12406 11152 12458
rect 11340 12406 11341 12458
rect 11151 12394 11157 12406
rect 11335 12394 11341 12406
rect 11151 12342 11152 12394
rect 11340 12342 11341 12394
rect 11151 12329 11157 12342
rect 11335 12329 11341 12342
rect 11151 12277 11152 12329
rect 11340 12277 11341 12329
rect 11151 12264 11157 12277
rect 11335 12264 11341 12277
rect 11151 12212 11152 12264
rect 11340 12212 11341 12264
rect 11151 12199 11157 12212
rect 11335 12199 11341 12212
rect 11151 12147 11152 12199
rect 11340 12147 11341 12199
rect 11151 12134 11157 12147
rect 11335 12134 11341 12147
rect 11151 12082 11152 12134
rect 11340 12082 11341 12134
rect 11151 12069 11157 12082
rect 11335 12069 11341 12082
rect 11151 12017 11152 12069
rect 11340 12017 11341 12069
rect 11151 12004 11157 12017
rect 11335 12004 11341 12017
rect 11151 11952 11152 12004
rect 11340 11952 11341 12004
rect 11151 11939 11157 11952
rect 11335 11939 11341 11952
rect 11151 11887 11152 11939
rect 11340 11887 11341 11939
rect 11151 11874 11157 11887
rect 11335 11874 11341 11887
rect 11151 11822 11152 11874
rect 11340 11822 11341 11874
rect 11151 11809 11157 11822
rect 11335 11809 11341 11822
rect 11151 11757 11152 11809
rect 11340 11757 11341 11809
rect 11151 11744 11157 11757
rect 11335 11744 11341 11757
rect 11151 11692 11152 11744
rect 11340 11692 11341 11744
rect 11151 11679 11157 11692
rect 11335 11679 11341 11692
rect 11151 11627 11152 11679
rect 11340 11627 11341 11679
rect 11151 11614 11157 11627
rect 11335 11614 11341 11627
rect 11151 11562 11152 11614
rect 11340 11562 11341 11614
rect 11151 10160 11157 11562
rect 11335 10160 11341 11562
rect 11151 10121 11341 10160
rect 11151 10087 11157 10121
rect 11191 10087 11229 10121
rect 11263 10087 11301 10121
rect 11335 10087 11341 10121
rect 11151 10048 11341 10087
rect 11151 10014 11157 10048
rect 11191 10014 11229 10048
rect 11263 10014 11301 10048
rect 11335 10014 11341 10048
rect 11151 9975 11341 10014
rect 11151 9941 11157 9975
rect 11191 9941 11229 9975
rect 11263 9941 11301 9975
rect 11335 9941 11341 9975
rect 11151 9902 11341 9941
rect 11151 9868 11157 9902
rect 11191 9868 11229 9902
rect 11263 9868 11301 9902
rect 11335 9868 11341 9902
rect 11151 9829 11341 9868
rect 11151 9795 11157 9829
rect 11191 9795 11229 9829
rect 11263 9795 11301 9829
rect 11335 9795 11341 9829
rect 11151 9756 11341 9795
rect 11151 9722 11157 9756
rect 11191 9722 11229 9756
rect 11263 9722 11301 9756
rect 11335 9722 11341 9756
rect 11151 9683 11341 9722
rect 11151 9649 11157 9683
rect 11191 9649 11229 9683
rect 11263 9649 11301 9683
rect 11335 9649 11341 9683
rect 11151 9610 11341 9649
rect 11151 9576 11157 9610
rect 11191 9576 11229 9610
rect 11263 9576 11301 9610
rect 11335 9576 11341 9610
rect 11151 9537 11341 9576
rect 11151 9503 11157 9537
rect 11191 9503 11229 9537
rect 11263 9503 11301 9537
rect 11335 9503 11341 9537
rect 11151 9491 11341 9503
rect 11641 37997 11771 38003
rect 11693 37945 11719 37997
rect 11641 37929 11771 37945
rect 11693 37877 11719 37929
rect 11641 37861 11771 37877
rect 11693 37809 11719 37861
rect 11641 37793 11771 37809
rect 11693 37741 11719 37793
rect 11641 37725 11771 37741
rect 11693 37673 11719 37725
rect 11641 37657 11771 37673
rect 11693 37605 11719 37657
rect 11641 37589 11771 37605
rect 11693 37537 11719 37589
rect 11641 37521 11771 37537
rect 11693 37469 11719 37521
rect 11641 37453 11771 37469
rect 11693 37401 11719 37453
rect 11641 37385 11771 37401
rect 11693 37333 11719 37385
rect 11641 37318 11771 37333
rect 11693 37266 11719 37318
rect 11641 37251 11771 37266
rect 11693 37199 11719 37251
rect 11641 37184 11771 37199
rect 11693 37132 11719 37184
rect 11641 37117 11771 37132
rect 11693 37065 11719 37117
rect 11641 34225 11771 37065
rect 11693 34173 11719 34225
rect 11641 34161 11771 34173
rect 11693 34109 11719 34161
rect 11641 34097 11771 34109
rect 11693 34045 11719 34097
rect 11641 34033 11771 34045
rect 11693 33981 11719 34033
rect 11641 33969 11771 33981
rect 11693 33917 11719 33969
rect 11641 33905 11771 33917
rect 11693 33853 11719 33905
rect 11641 33841 11771 33853
rect 11693 33789 11719 33841
rect 11641 33777 11771 33789
rect 11693 33725 11719 33777
rect 11641 33713 11771 33725
rect 11693 33661 11719 33713
rect 11641 33649 11771 33661
rect 11693 33597 11719 33649
rect 11641 33585 11771 33597
rect 11693 33533 11719 33585
rect 11641 33521 11771 33533
rect 11693 33469 11719 33521
rect 11641 33457 11771 33469
rect 11693 33405 11719 33457
rect 11641 33393 11771 33405
rect 11693 33341 11719 33393
rect 11641 33329 11771 33341
rect 11693 33277 11719 33329
rect 11641 33264 11771 33277
rect 11693 33212 11719 33264
rect 11641 33199 11771 33212
rect 11693 33147 11719 33199
rect 11641 33134 11771 33147
rect 11693 33082 11719 33134
rect 11641 33069 11771 33082
rect 11693 33017 11719 33069
rect 11641 33004 11771 33017
rect 11693 32952 11719 33004
rect 11641 32939 11771 32952
rect 11693 32887 11719 32939
rect 11641 32874 11771 32887
rect 11693 32822 11719 32874
rect 11641 32809 11771 32822
rect 11693 32757 11719 32809
rect 11641 32744 11771 32757
rect 11693 32692 11719 32744
rect 11641 32679 11771 32692
rect 11693 32627 11719 32679
rect 11641 32614 11771 32627
rect 11693 32562 11719 32614
rect 11641 32549 11771 32562
rect 11693 32497 11719 32549
rect 11641 29625 11771 32497
rect 11693 29573 11719 29625
rect 11641 29561 11771 29573
rect 11693 29509 11719 29561
rect 11641 29497 11771 29509
rect 11693 29445 11719 29497
rect 11641 29433 11771 29445
rect 11693 29381 11719 29433
rect 11641 29369 11771 29381
rect 11693 29317 11719 29369
rect 11641 29305 11771 29317
rect 11693 29253 11719 29305
rect 11641 29241 11771 29253
rect 11693 29189 11719 29241
rect 11641 29177 11771 29189
rect 11693 29125 11719 29177
rect 11641 29113 11771 29125
rect 11693 29061 11719 29113
rect 11641 29049 11771 29061
rect 11693 28997 11719 29049
rect 11641 28985 11771 28997
rect 11693 28933 11719 28985
rect 11641 28921 11771 28933
rect 11693 28869 11719 28921
rect 11641 28857 11771 28869
rect 11693 28805 11719 28857
rect 11641 28793 11771 28805
rect 11693 28741 11719 28793
rect 11641 28729 11771 28741
rect 11693 28677 11719 28729
rect 11641 28664 11771 28677
rect 11693 28612 11719 28664
rect 11641 28599 11771 28612
rect 11693 28547 11719 28599
rect 11641 28534 11771 28547
rect 11693 28482 11719 28534
rect 11641 28469 11771 28482
rect 11693 28417 11719 28469
rect 11641 28404 11771 28417
rect 11693 28352 11719 28404
rect 11641 28339 11771 28352
rect 11693 28287 11719 28339
rect 11641 28274 11771 28287
rect 11693 28222 11719 28274
rect 11641 28209 11771 28222
rect 11693 28157 11719 28209
rect 11641 28144 11771 28157
rect 11693 28092 11719 28144
rect 11641 28079 11771 28092
rect 11693 28027 11719 28079
rect 11641 28014 11771 28027
rect 11693 27962 11719 28014
rect 11641 27949 11771 27962
rect 11693 27897 11719 27949
rect 11641 25025 11771 27897
rect 11693 24973 11719 25025
rect 11641 24961 11771 24973
rect 11693 24909 11719 24961
rect 11641 24897 11771 24909
rect 11693 24845 11719 24897
rect 11641 24833 11771 24845
rect 11693 24781 11719 24833
rect 11641 24769 11771 24781
rect 11693 24717 11719 24769
rect 11641 24705 11771 24717
rect 11693 24653 11719 24705
rect 11641 24641 11771 24653
rect 11693 24589 11719 24641
rect 11641 24577 11771 24589
rect 11693 24525 11719 24577
rect 11641 24513 11771 24525
rect 11693 24461 11719 24513
rect 11641 24449 11771 24461
rect 11693 24397 11719 24449
rect 11641 24385 11771 24397
rect 11693 24333 11719 24385
rect 11641 24321 11771 24333
rect 11693 24269 11719 24321
rect 11641 24257 11771 24269
rect 11693 24205 11719 24257
rect 11641 24193 11771 24205
rect 11693 24141 11719 24193
rect 11641 24129 11771 24141
rect 11693 24077 11719 24129
rect 11641 24064 11771 24077
rect 11693 24012 11719 24064
rect 11641 23999 11771 24012
rect 11693 23947 11719 23999
rect 11641 23934 11771 23947
rect 11693 23882 11719 23934
rect 11641 23869 11771 23882
rect 11693 23817 11719 23869
rect 11641 23804 11771 23817
rect 11693 23752 11719 23804
rect 11641 23739 11771 23752
rect 11693 23687 11719 23739
rect 11641 23674 11771 23687
rect 11693 23622 11719 23674
rect 11641 23609 11771 23622
rect 11693 23557 11719 23609
rect 11641 23544 11771 23557
rect 11693 23492 11719 23544
rect 11641 23479 11771 23492
rect 11693 23427 11719 23479
rect 11641 23414 11771 23427
rect 11693 23362 11719 23414
rect 11641 23349 11771 23362
rect 11693 23297 11719 23349
rect 11641 20425 11771 23297
rect 11693 20373 11719 20425
rect 11641 20361 11771 20373
rect 11693 20309 11719 20361
rect 11641 20297 11771 20309
rect 11693 20245 11719 20297
rect 11641 20233 11771 20245
rect 11693 20181 11719 20233
rect 11641 20169 11771 20181
rect 11693 20117 11719 20169
rect 11641 20105 11771 20117
rect 11693 20053 11719 20105
rect 11641 20041 11771 20053
rect 11693 19989 11719 20041
rect 11641 19977 11771 19989
rect 11693 19925 11719 19977
rect 11641 19913 11771 19925
rect 11693 19861 11719 19913
rect 11641 19849 11771 19861
rect 11693 19797 11719 19849
rect 11641 19785 11771 19797
rect 11693 19733 11719 19785
rect 11641 19721 11771 19733
rect 11693 19669 11719 19721
rect 11641 19657 11771 19669
rect 11693 19605 11719 19657
rect 11641 19593 11771 19605
rect 11693 19541 11719 19593
rect 11641 19529 11771 19541
rect 11693 19477 11719 19529
rect 11641 19464 11771 19477
rect 11693 19412 11719 19464
rect 11641 19399 11771 19412
rect 11693 19347 11719 19399
rect 11641 19334 11771 19347
rect 11693 19282 11719 19334
rect 11641 19269 11771 19282
rect 11693 19217 11719 19269
rect 11641 19204 11771 19217
rect 11693 19152 11719 19204
rect 11641 19139 11771 19152
rect 11693 19087 11719 19139
rect 11641 19074 11771 19087
rect 11693 19022 11719 19074
rect 11641 19009 11771 19022
rect 11693 18957 11719 19009
rect 11641 18944 11771 18957
rect 11693 18892 11719 18944
rect 11641 18879 11771 18892
rect 11693 18827 11719 18879
rect 11641 18814 11771 18827
rect 11693 18762 11719 18814
rect 11641 18749 11771 18762
rect 11693 18697 11719 18749
rect 11641 15825 11771 18697
rect 11693 15773 11719 15825
rect 11641 15761 11771 15773
rect 11693 15709 11719 15761
rect 11641 15697 11771 15709
rect 11693 15645 11719 15697
rect 11641 15633 11771 15645
rect 11693 15581 11719 15633
rect 11641 15569 11771 15581
rect 11693 15517 11719 15569
rect 11641 15505 11771 15517
rect 11693 15453 11719 15505
rect 11641 15441 11771 15453
rect 11693 15389 11719 15441
rect 11641 15377 11771 15389
rect 11693 15325 11719 15377
rect 11641 15313 11771 15325
rect 11693 15261 11719 15313
rect 11641 15249 11771 15261
rect 11693 15197 11719 15249
rect 11641 15185 11771 15197
rect 11693 15133 11719 15185
rect 11641 15121 11771 15133
rect 11693 15069 11719 15121
rect 11641 15057 11771 15069
rect 11693 15005 11719 15057
rect 11641 14993 11771 15005
rect 11693 14941 11719 14993
rect 11641 14929 11771 14941
rect 11693 14877 11719 14929
rect 11641 14864 11771 14877
rect 11693 14812 11719 14864
rect 11641 14799 11771 14812
rect 11693 14747 11719 14799
rect 11641 14734 11771 14747
rect 11693 14682 11719 14734
rect 11641 14669 11771 14682
rect 11693 14617 11719 14669
rect 11641 14604 11771 14617
rect 11693 14552 11719 14604
rect 11641 14539 11771 14552
rect 11693 14487 11719 14539
rect 11641 14474 11771 14487
rect 11693 14422 11719 14474
rect 11641 14409 11771 14422
rect 11693 14357 11719 14409
rect 11641 14344 11771 14357
rect 11693 14292 11719 14344
rect 11641 14279 11771 14292
rect 11693 14227 11719 14279
rect 11641 14214 11771 14227
rect 11693 14162 11719 14214
rect 11641 14149 11771 14162
rect 11693 14097 11719 14149
rect 11641 11225 11771 14097
rect 11693 11173 11719 11225
rect 11641 11161 11771 11173
rect 11693 11109 11719 11161
rect 11641 11097 11771 11109
rect 11693 11045 11719 11097
rect 11641 11033 11771 11045
rect 11693 10981 11719 11033
rect 11641 10969 11771 10981
rect 11693 10917 11719 10969
rect 11641 10905 11771 10917
rect 11693 10853 11719 10905
rect 11641 10841 11771 10853
rect 11693 10789 11719 10841
rect 11641 10777 11771 10789
rect 11693 10725 11719 10777
rect 11641 10713 11771 10725
rect 11693 10661 11719 10713
rect 11641 10649 11771 10661
rect 11693 10597 11719 10649
rect 11641 10585 11771 10597
rect 11693 10533 11719 10585
rect 11641 10521 11771 10533
rect 11693 10469 11719 10521
rect 11641 10457 11771 10469
rect 11693 10405 11719 10457
rect 11641 10393 11771 10405
rect 11693 10341 11719 10393
rect 11641 10329 11771 10341
rect 11693 10277 11719 10329
rect 11641 10264 11771 10277
rect 11693 10212 11719 10264
rect 11641 10199 11771 10212
rect 11693 10147 11719 10199
rect 11641 10134 11771 10147
rect 11693 10082 11719 10134
rect 11641 10069 11771 10082
rect 11693 10017 11719 10069
rect 11641 10004 11771 10017
rect 11693 9952 11719 10004
rect 11641 9939 11771 9952
rect 11693 9887 11719 9939
rect 11641 9874 11771 9887
rect 11693 9822 11719 9874
rect 11641 9809 11771 9822
rect 11693 9757 11719 9809
rect 11641 9744 11771 9757
rect 11693 9692 11719 9744
rect 11641 9679 11771 9692
rect 11693 9627 11719 9679
rect 11641 9614 11771 9627
rect 11693 9562 11719 9614
rect 11641 9549 11771 9562
rect 11693 9497 11719 9549
rect 11641 9491 11771 9497
rect 12071 37979 12077 38013
rect 12111 37979 12149 38013
rect 12183 37979 12221 38013
rect 12255 37979 12261 38013
rect 12991 39028 13181 39040
rect 12991 39009 12997 39028
rect 13175 39009 13181 39028
rect 12991 38957 12992 39009
rect 13180 38957 13181 39009
rect 12991 38945 12997 38957
rect 13175 38945 13181 38957
rect 12991 38893 12992 38945
rect 13180 38893 13181 38945
rect 12991 38881 12997 38893
rect 13175 38881 13181 38893
rect 12991 38829 12992 38881
rect 13180 38829 13181 38881
rect 12991 38817 12997 38829
rect 13175 38817 13181 38829
rect 12991 38765 12992 38817
rect 13180 38765 13181 38817
rect 12991 38753 12997 38765
rect 13175 38753 13181 38765
rect 12991 38701 12992 38753
rect 13180 38701 13181 38753
rect 12991 38689 12997 38701
rect 13175 38689 13181 38701
rect 12991 38637 12992 38689
rect 13180 38637 13181 38689
rect 12991 38625 12997 38637
rect 13175 38625 13181 38637
rect 12991 38573 12992 38625
rect 13180 38573 13181 38625
rect 12991 38560 12997 38573
rect 13175 38560 13181 38573
rect 12991 38508 12992 38560
rect 13180 38508 13181 38560
rect 12991 38495 12997 38508
rect 13175 38495 13181 38508
rect 12991 38443 12992 38495
rect 13044 38443 13060 38490
rect 13112 38443 13128 38490
rect 13180 38443 13181 38495
rect 12991 38430 12997 38443
rect 13031 38430 13069 38443
rect 13103 38430 13141 38443
rect 13175 38430 13181 38443
rect 12991 38378 12992 38430
rect 13044 38378 13060 38430
rect 13112 38378 13128 38430
rect 13180 38378 13181 38430
rect 12991 38365 12997 38378
rect 13031 38365 13069 38378
rect 13103 38365 13141 38378
rect 13175 38365 13181 38378
rect 12991 38313 12992 38365
rect 13044 38313 13060 38365
rect 13112 38313 13128 38365
rect 13180 38313 13181 38365
rect 12991 38305 13181 38313
rect 12991 38300 12997 38305
rect 13031 38300 13069 38305
rect 13103 38300 13141 38305
rect 13175 38300 13181 38305
rect 12991 38248 12992 38300
rect 13044 38248 13060 38300
rect 13112 38248 13128 38300
rect 13180 38248 13181 38300
rect 12991 38235 13181 38248
rect 12991 38183 12992 38235
rect 13044 38183 13060 38235
rect 13112 38183 13128 38235
rect 13180 38183 13181 38235
rect 12991 38170 13181 38183
rect 12991 38118 12992 38170
rect 13044 38118 13060 38170
rect 13112 38118 13128 38170
rect 13180 38118 13181 38170
rect 12991 38086 13181 38118
rect 12991 38052 12997 38086
rect 13031 38052 13069 38086
rect 13103 38052 13141 38086
rect 13175 38052 13181 38086
rect 12991 38013 13181 38052
rect 12071 37940 12261 37979
rect 12071 37906 12077 37940
rect 12111 37906 12149 37940
rect 12183 37906 12221 37940
rect 12255 37906 12261 37940
rect 12071 37867 12261 37906
rect 12071 37833 12077 37867
rect 12111 37833 12149 37867
rect 12183 37833 12221 37867
rect 12255 37833 12261 37867
rect 12071 37794 12261 37833
rect 12071 37760 12077 37794
rect 12111 37760 12149 37794
rect 12183 37760 12221 37794
rect 12255 37760 12261 37794
rect 12071 37721 12261 37760
rect 12071 37687 12077 37721
rect 12111 37687 12149 37721
rect 12183 37687 12221 37721
rect 12255 37687 12261 37721
rect 12071 37648 12261 37687
rect 12071 37614 12077 37648
rect 12111 37614 12149 37648
rect 12183 37614 12221 37648
rect 12255 37614 12261 37648
rect 12071 37575 12261 37614
rect 12071 37541 12077 37575
rect 12111 37541 12149 37575
rect 12183 37541 12221 37575
rect 12255 37541 12261 37575
rect 12071 37502 12261 37541
rect 12071 37468 12077 37502
rect 12111 37468 12149 37502
rect 12183 37468 12221 37502
rect 12255 37468 12261 37502
rect 12071 37429 12261 37468
rect 12071 37395 12077 37429
rect 12111 37395 12149 37429
rect 12183 37395 12221 37429
rect 12255 37395 12261 37429
rect 12071 37356 12261 37395
rect 12071 37322 12077 37356
rect 12111 37322 12149 37356
rect 12183 37322 12221 37356
rect 12255 37322 12261 37356
rect 12071 37283 12261 37322
rect 12071 37249 12077 37283
rect 12111 37249 12149 37283
rect 12183 37249 12221 37283
rect 12255 37249 12261 37283
rect 12071 37210 12261 37249
rect 12071 37176 12077 37210
rect 12111 37176 12149 37210
rect 12183 37176 12221 37210
rect 12255 37176 12261 37210
rect 12071 37137 12261 37176
rect 12071 37103 12077 37137
rect 12111 37103 12149 37137
rect 12183 37103 12221 37137
rect 12255 37103 12261 37137
rect 12071 36353 12261 37103
rect 12071 32503 12077 36353
rect 12255 32503 12261 36353
rect 12071 31753 12261 32503
rect 12071 27903 12077 31753
rect 12255 27903 12261 31753
rect 12071 27153 12261 27903
rect 12071 23303 12077 27153
rect 12255 23303 12261 27153
rect 12071 22562 12261 23303
rect 12071 19360 12077 22562
rect 12255 19360 12261 22562
rect 12071 19321 12261 19360
rect 12071 19287 12077 19321
rect 12111 19287 12149 19321
rect 12183 19287 12221 19321
rect 12255 19287 12261 19321
rect 12071 19248 12261 19287
rect 12071 19214 12077 19248
rect 12111 19214 12149 19248
rect 12183 19214 12221 19248
rect 12255 19214 12261 19248
rect 12071 19175 12261 19214
rect 12071 19141 12077 19175
rect 12111 19141 12149 19175
rect 12183 19141 12221 19175
rect 12255 19141 12261 19175
rect 12071 19102 12261 19141
rect 12071 19068 12077 19102
rect 12111 19068 12149 19102
rect 12183 19068 12221 19102
rect 12255 19068 12261 19102
rect 12071 19029 12261 19068
rect 12071 18995 12077 19029
rect 12111 18995 12149 19029
rect 12183 18995 12221 19029
rect 12255 18995 12261 19029
rect 12071 18956 12261 18995
rect 12071 18922 12077 18956
rect 12111 18922 12149 18956
rect 12183 18922 12221 18956
rect 12255 18922 12261 18956
rect 12071 18883 12261 18922
rect 12071 18849 12077 18883
rect 12111 18849 12149 18883
rect 12183 18849 12221 18883
rect 12255 18849 12261 18883
rect 12071 18810 12261 18849
rect 12071 18776 12077 18810
rect 12111 18776 12149 18810
rect 12183 18776 12221 18810
rect 12255 18776 12261 18810
rect 12071 18737 12261 18776
rect 12071 18703 12077 18737
rect 12111 18703 12149 18737
rect 12183 18703 12221 18737
rect 12255 18703 12261 18737
rect 12071 17953 12261 18703
rect 12071 14103 12077 17953
rect 12255 14103 12261 17953
rect 12071 13362 12261 14103
rect 12071 10160 12077 13362
rect 12255 10160 12261 13362
rect 12071 10121 12261 10160
rect 12071 10087 12077 10121
rect 12111 10087 12149 10121
rect 12183 10087 12221 10121
rect 12255 10087 12261 10121
rect 12071 10048 12261 10087
rect 12071 10014 12077 10048
rect 12111 10014 12149 10048
rect 12183 10014 12221 10048
rect 12255 10014 12261 10048
rect 12071 9975 12261 10014
rect 12071 9941 12077 9975
rect 12111 9941 12149 9975
rect 12183 9941 12221 9975
rect 12255 9941 12261 9975
rect 12071 9902 12261 9941
rect 12071 9868 12077 9902
rect 12111 9868 12149 9902
rect 12183 9868 12221 9902
rect 12255 9868 12261 9902
rect 12071 9829 12261 9868
rect 12071 9795 12077 9829
rect 12111 9795 12149 9829
rect 12183 9795 12221 9829
rect 12255 9795 12261 9829
rect 12071 9756 12261 9795
rect 12071 9722 12077 9756
rect 12111 9722 12149 9756
rect 12183 9722 12221 9756
rect 12255 9722 12261 9756
rect 12071 9683 12261 9722
rect 12071 9649 12077 9683
rect 12111 9649 12149 9683
rect 12183 9649 12221 9683
rect 12255 9649 12261 9683
rect 12071 9610 12261 9649
rect 12071 9576 12077 9610
rect 12111 9576 12149 9610
rect 12183 9576 12221 9610
rect 12255 9576 12261 9610
rect 12071 9537 12261 9576
rect 12071 9503 12077 9537
rect 12111 9503 12149 9537
rect 12183 9503 12221 9537
rect 12255 9503 12261 9537
rect 12071 9491 12261 9503
rect 12561 37997 12691 38003
rect 12613 37945 12639 37997
rect 12561 37929 12691 37945
rect 12613 37877 12639 37929
rect 12561 37861 12691 37877
rect 12613 37809 12639 37861
rect 12561 37793 12691 37809
rect 12613 37741 12639 37793
rect 12561 37725 12691 37741
rect 12613 37673 12639 37725
rect 12561 37657 12691 37673
rect 12613 37605 12639 37657
rect 12561 37589 12691 37605
rect 12613 37537 12639 37589
rect 12561 37521 12691 37537
rect 12613 37469 12639 37521
rect 12561 37453 12691 37469
rect 12613 37401 12639 37453
rect 12561 37385 12691 37401
rect 12613 37333 12639 37385
rect 12561 37318 12691 37333
rect 12613 37266 12639 37318
rect 12561 37251 12691 37266
rect 12613 37199 12639 37251
rect 12561 37184 12691 37199
rect 12613 37132 12639 37184
rect 12561 37117 12691 37132
rect 12613 37065 12639 37117
rect 12561 34225 12691 37065
rect 12613 34173 12639 34225
rect 12561 34161 12691 34173
rect 12613 34109 12639 34161
rect 12561 34097 12691 34109
rect 12613 34045 12639 34097
rect 12561 34033 12691 34045
rect 12613 33981 12639 34033
rect 12561 33969 12691 33981
rect 12613 33917 12639 33969
rect 12561 33905 12691 33917
rect 12613 33853 12639 33905
rect 12561 33841 12691 33853
rect 12613 33789 12639 33841
rect 12561 33777 12691 33789
rect 12613 33725 12639 33777
rect 12561 33713 12691 33725
rect 12613 33661 12639 33713
rect 12561 33649 12691 33661
rect 12613 33597 12639 33649
rect 12561 33585 12691 33597
rect 12613 33533 12639 33585
rect 12561 33521 12691 33533
rect 12613 33469 12639 33521
rect 12561 33457 12691 33469
rect 12613 33405 12639 33457
rect 12561 33393 12691 33405
rect 12613 33341 12639 33393
rect 12561 33329 12691 33341
rect 12613 33277 12639 33329
rect 12561 33264 12691 33277
rect 12613 33212 12639 33264
rect 12561 33199 12691 33212
rect 12613 33147 12639 33199
rect 12561 33134 12691 33147
rect 12613 33082 12639 33134
rect 12561 33069 12691 33082
rect 12613 33017 12639 33069
rect 12561 33004 12691 33017
rect 12613 32952 12639 33004
rect 12561 32939 12691 32952
rect 12613 32887 12639 32939
rect 12561 32874 12691 32887
rect 12613 32822 12639 32874
rect 12561 32809 12691 32822
rect 12613 32757 12639 32809
rect 12561 32744 12691 32757
rect 12613 32692 12639 32744
rect 12561 32679 12691 32692
rect 12613 32627 12639 32679
rect 12561 32614 12691 32627
rect 12613 32562 12639 32614
rect 12561 32549 12691 32562
rect 12613 32497 12639 32549
rect 12561 29625 12691 32497
rect 12613 29573 12639 29625
rect 12561 29561 12691 29573
rect 12613 29509 12639 29561
rect 12561 29497 12691 29509
rect 12613 29445 12639 29497
rect 12561 29433 12691 29445
rect 12613 29381 12639 29433
rect 12561 29369 12691 29381
rect 12613 29317 12639 29369
rect 12561 29305 12691 29317
rect 12613 29253 12639 29305
rect 12561 29241 12691 29253
rect 12613 29189 12639 29241
rect 12561 29177 12691 29189
rect 12613 29125 12639 29177
rect 12561 29113 12691 29125
rect 12613 29061 12639 29113
rect 12561 29049 12691 29061
rect 12613 28997 12639 29049
rect 12561 28985 12691 28997
rect 12613 28933 12639 28985
rect 12561 28921 12691 28933
rect 12613 28869 12639 28921
rect 12561 28857 12691 28869
rect 12613 28805 12639 28857
rect 12561 28793 12691 28805
rect 12613 28741 12639 28793
rect 12561 28729 12691 28741
rect 12613 28677 12639 28729
rect 12561 28664 12691 28677
rect 12613 28612 12639 28664
rect 12561 28599 12691 28612
rect 12613 28547 12639 28599
rect 12561 28534 12691 28547
rect 12613 28482 12639 28534
rect 12561 28469 12691 28482
rect 12613 28417 12639 28469
rect 12561 28404 12691 28417
rect 12613 28352 12639 28404
rect 12561 28339 12691 28352
rect 12613 28287 12639 28339
rect 12561 28274 12691 28287
rect 12613 28222 12639 28274
rect 12561 28209 12691 28222
rect 12613 28157 12639 28209
rect 12561 28144 12691 28157
rect 12613 28092 12639 28144
rect 12561 28079 12691 28092
rect 12613 28027 12639 28079
rect 12561 28014 12691 28027
rect 12613 27962 12639 28014
rect 12561 27949 12691 27962
rect 12613 27897 12639 27949
rect 12561 25025 12691 27897
rect 12613 24973 12639 25025
rect 12561 24961 12691 24973
rect 12613 24909 12639 24961
rect 12561 24897 12691 24909
rect 12613 24845 12639 24897
rect 12561 24833 12691 24845
rect 12613 24781 12639 24833
rect 12561 24769 12691 24781
rect 12613 24717 12639 24769
rect 12561 24705 12691 24717
rect 12613 24653 12639 24705
rect 12561 24641 12691 24653
rect 12613 24589 12639 24641
rect 12561 24577 12691 24589
rect 12613 24525 12639 24577
rect 12561 24513 12691 24525
rect 12613 24461 12639 24513
rect 12561 24449 12691 24461
rect 12613 24397 12639 24449
rect 12561 24385 12691 24397
rect 12613 24333 12639 24385
rect 12561 24321 12691 24333
rect 12613 24269 12639 24321
rect 12561 24257 12691 24269
rect 12613 24205 12639 24257
rect 12561 24193 12691 24205
rect 12613 24141 12639 24193
rect 12561 24129 12691 24141
rect 12613 24077 12639 24129
rect 12561 24064 12691 24077
rect 12613 24012 12639 24064
rect 12561 23999 12691 24012
rect 12613 23947 12639 23999
rect 12561 23934 12691 23947
rect 12613 23882 12639 23934
rect 12561 23869 12691 23882
rect 12613 23817 12639 23869
rect 12561 23804 12691 23817
rect 12613 23752 12639 23804
rect 12561 23739 12691 23752
rect 12613 23687 12639 23739
rect 12561 23674 12691 23687
rect 12613 23622 12639 23674
rect 12561 23609 12691 23622
rect 12613 23557 12639 23609
rect 12561 23544 12691 23557
rect 12613 23492 12639 23544
rect 12561 23479 12691 23492
rect 12613 23427 12639 23479
rect 12561 23414 12691 23427
rect 12613 23362 12639 23414
rect 12561 23349 12691 23362
rect 12613 23297 12639 23349
rect 12561 20425 12691 23297
rect 12613 20373 12639 20425
rect 12561 20361 12691 20373
rect 12613 20309 12639 20361
rect 12561 20297 12691 20309
rect 12613 20245 12639 20297
rect 12561 20233 12691 20245
rect 12613 20181 12639 20233
rect 12561 20169 12691 20181
rect 12613 20117 12639 20169
rect 12561 20105 12691 20117
rect 12613 20053 12639 20105
rect 12561 20041 12691 20053
rect 12613 19989 12639 20041
rect 12561 19977 12691 19989
rect 12613 19925 12639 19977
rect 12561 19913 12691 19925
rect 12613 19861 12639 19913
rect 12561 19849 12691 19861
rect 12613 19797 12639 19849
rect 12561 19785 12691 19797
rect 12613 19733 12639 19785
rect 12561 19721 12691 19733
rect 12613 19669 12639 19721
rect 12561 19657 12691 19669
rect 12613 19605 12639 19657
rect 12561 19593 12691 19605
rect 12613 19541 12639 19593
rect 12561 19529 12691 19541
rect 12613 19477 12639 19529
rect 12561 19464 12691 19477
rect 12613 19412 12639 19464
rect 12561 19399 12691 19412
rect 12613 19347 12639 19399
rect 12561 19334 12691 19347
rect 12613 19282 12639 19334
rect 12561 19269 12691 19282
rect 12613 19217 12639 19269
rect 12561 19204 12691 19217
rect 12613 19152 12639 19204
rect 12561 19139 12691 19152
rect 12613 19087 12639 19139
rect 12561 19074 12691 19087
rect 12613 19022 12639 19074
rect 12561 19009 12691 19022
rect 12613 18957 12639 19009
rect 12561 18944 12691 18957
rect 12613 18892 12639 18944
rect 12561 18879 12691 18892
rect 12613 18827 12639 18879
rect 12561 18814 12691 18827
rect 12613 18762 12639 18814
rect 12561 18749 12691 18762
rect 12613 18697 12639 18749
rect 12561 15825 12691 18697
rect 12613 15773 12639 15825
rect 12561 15761 12691 15773
rect 12613 15709 12639 15761
rect 12561 15697 12691 15709
rect 12613 15645 12639 15697
rect 12561 15633 12691 15645
rect 12613 15581 12639 15633
rect 12561 15569 12691 15581
rect 12613 15517 12639 15569
rect 12561 15505 12691 15517
rect 12613 15453 12639 15505
rect 12561 15441 12691 15453
rect 12613 15389 12639 15441
rect 12561 15377 12691 15389
rect 12613 15325 12639 15377
rect 12561 15313 12691 15325
rect 12613 15261 12639 15313
rect 12561 15249 12691 15261
rect 12613 15197 12639 15249
rect 12561 15185 12691 15197
rect 12613 15133 12639 15185
rect 12561 15121 12691 15133
rect 12613 15069 12639 15121
rect 12561 15057 12691 15069
rect 12613 15005 12639 15057
rect 12561 14993 12691 15005
rect 12613 14941 12639 14993
rect 12561 14929 12691 14941
rect 12613 14877 12639 14929
rect 12561 14864 12691 14877
rect 12613 14812 12639 14864
rect 12561 14799 12691 14812
rect 12613 14747 12639 14799
rect 12561 14734 12691 14747
rect 12613 14682 12639 14734
rect 12561 14669 12691 14682
rect 12613 14617 12639 14669
rect 12561 14604 12691 14617
rect 12613 14552 12639 14604
rect 12561 14539 12691 14552
rect 12613 14487 12639 14539
rect 12561 14474 12691 14487
rect 12613 14422 12639 14474
rect 12561 14409 12691 14422
rect 12613 14357 12639 14409
rect 12561 14344 12691 14357
rect 12613 14292 12639 14344
rect 12561 14279 12691 14292
rect 12613 14227 12639 14279
rect 12561 14214 12691 14227
rect 12613 14162 12639 14214
rect 12561 14149 12691 14162
rect 12613 14097 12639 14149
rect 12561 11225 12691 14097
rect 12613 11173 12639 11225
rect 12561 11161 12691 11173
rect 12613 11109 12639 11161
rect 12561 11097 12691 11109
rect 12613 11045 12639 11097
rect 12561 11033 12691 11045
rect 12613 10981 12639 11033
rect 12561 10969 12691 10981
rect 12613 10917 12639 10969
rect 12561 10905 12691 10917
rect 12613 10853 12639 10905
rect 12561 10841 12691 10853
rect 12613 10789 12639 10841
rect 12561 10777 12691 10789
rect 12613 10725 12639 10777
rect 12561 10713 12691 10725
rect 12613 10661 12639 10713
rect 12561 10649 12691 10661
rect 12613 10597 12639 10649
rect 12561 10585 12691 10597
rect 12613 10533 12639 10585
rect 12561 10521 12691 10533
rect 12613 10469 12639 10521
rect 12561 10457 12691 10469
rect 12613 10405 12639 10457
rect 12561 10393 12691 10405
rect 12613 10341 12639 10393
rect 12561 10329 12691 10341
rect 12613 10277 12639 10329
rect 12561 10264 12691 10277
rect 12613 10212 12639 10264
rect 12561 10199 12691 10212
rect 12613 10147 12639 10199
rect 12561 10134 12691 10147
rect 12613 10082 12639 10134
rect 12561 10069 12691 10082
rect 12613 10017 12639 10069
rect 12561 10004 12691 10017
rect 12613 9952 12639 10004
rect 12561 9939 12691 9952
rect 12613 9887 12639 9939
rect 12561 9874 12691 9887
rect 12613 9822 12639 9874
rect 12561 9809 12691 9822
rect 12613 9757 12639 9809
rect 12561 9744 12691 9757
rect 12613 9692 12639 9744
rect 12561 9679 12691 9692
rect 12613 9627 12639 9679
rect 12561 9614 12691 9627
rect 12613 9562 12639 9614
rect 12561 9549 12691 9562
rect 12613 9497 12639 9549
rect 12561 9491 12691 9497
rect 12991 37979 12997 38013
rect 13031 37979 13069 38013
rect 13103 37979 13141 38013
rect 13175 37979 13181 38013
rect 12991 37940 13181 37979
rect 12991 37906 12997 37940
rect 13031 37906 13069 37940
rect 13103 37906 13141 37940
rect 13175 37906 13181 37940
rect 12991 37867 13181 37906
rect 12991 37833 12997 37867
rect 13031 37833 13069 37867
rect 13103 37833 13141 37867
rect 13175 37833 13181 37867
rect 12991 37794 13181 37833
rect 12991 37760 12997 37794
rect 13031 37760 13069 37794
rect 13103 37760 13141 37794
rect 13175 37760 13181 37794
rect 12991 37721 13181 37760
rect 12991 37687 12997 37721
rect 13031 37687 13069 37721
rect 13103 37687 13141 37721
rect 13175 37687 13181 37721
rect 12991 37648 13181 37687
rect 12991 37614 12997 37648
rect 13031 37614 13069 37648
rect 13103 37614 13141 37648
rect 13175 37614 13181 37648
rect 12991 37575 13181 37614
rect 12991 37541 12997 37575
rect 13031 37541 13069 37575
rect 13103 37541 13141 37575
rect 13175 37541 13181 37575
rect 12991 37502 13181 37541
rect 12991 37468 12997 37502
rect 13031 37468 13069 37502
rect 13103 37468 13141 37502
rect 13175 37468 13181 37502
rect 12991 37429 13181 37468
rect 12991 37395 12997 37429
rect 13031 37395 13069 37429
rect 13103 37395 13141 37429
rect 13175 37395 13181 37429
rect 12991 37356 13181 37395
rect 12991 37322 12997 37356
rect 13031 37322 13069 37356
rect 13103 37322 13141 37356
rect 13175 37322 13181 37356
rect 12991 37283 13181 37322
rect 12991 37249 12997 37283
rect 13031 37249 13069 37283
rect 13103 37249 13141 37283
rect 13175 37249 13181 37283
rect 12991 37210 13181 37249
rect 12991 37176 12997 37210
rect 13031 37176 13069 37210
rect 13103 37176 13141 37210
rect 13175 37176 13181 37210
rect 12991 37137 13181 37176
rect 12991 37103 12997 37137
rect 13031 37103 13069 37137
rect 13103 37103 13141 37137
rect 13175 37103 13181 37137
rect 12991 36353 13181 37103
rect 12991 32503 12997 36353
rect 13175 32503 13181 36353
rect 13447 39036 13637 39074
rect 13447 39002 13453 39036
rect 13487 39035 13637 39036
rect 13487 39002 13525 39035
rect 13447 39001 13525 39002
rect 13559 39001 13597 39035
rect 13631 39001 13637 39035
rect 13447 38963 13637 39001
rect 13447 38929 13453 38963
rect 13487 38962 13637 38963
rect 13487 38929 13525 38962
rect 13447 38928 13525 38929
rect 13559 38928 13597 38962
rect 13631 38928 13637 38962
rect 13447 38890 13637 38928
rect 13447 38856 13453 38890
rect 13487 38889 13637 38890
rect 13487 38856 13525 38889
rect 13447 38855 13525 38856
rect 13559 38855 13597 38889
rect 13631 38855 13637 38889
rect 13447 38817 13637 38855
rect 13447 38783 13453 38817
rect 13487 38816 13637 38817
rect 13487 38783 13525 38816
rect 13447 38782 13525 38783
rect 13559 38782 13597 38816
rect 13631 38782 13637 38816
rect 13447 38744 13637 38782
rect 13447 38710 13453 38744
rect 13487 38743 13637 38744
rect 13487 38710 13525 38743
rect 13447 38709 13525 38710
rect 13559 38709 13597 38743
rect 13631 38709 13637 38743
rect 13447 38671 13637 38709
rect 13447 38637 13453 38671
rect 13487 38670 13637 38671
rect 13487 38637 13525 38670
rect 13447 38636 13525 38637
rect 13559 38636 13597 38670
rect 13631 38636 13637 38670
rect 13447 38598 13637 38636
rect 13447 38564 13453 38598
rect 13487 38597 13637 38598
rect 13487 38564 13525 38597
rect 13447 38563 13525 38564
rect 13559 38563 13597 38597
rect 13631 38563 13637 38597
rect 13447 38525 13637 38563
rect 13447 38491 13453 38525
rect 13487 38524 13637 38525
rect 13487 38491 13525 38524
rect 13447 38490 13525 38491
rect 13559 38490 13597 38524
rect 13631 38490 13637 38524
rect 13447 38452 13637 38490
rect 13447 38418 13453 38452
rect 13487 38451 13637 38452
rect 13487 38418 13525 38451
rect 13447 38417 13525 38418
rect 13559 38417 13597 38451
rect 13631 38417 13637 38451
rect 13447 38379 13637 38417
rect 13447 38345 13453 38379
rect 13487 38378 13637 38379
rect 13487 38345 13525 38378
rect 13447 38344 13525 38345
rect 13559 38344 13597 38378
rect 13631 38344 13637 38378
rect 13447 38306 13637 38344
rect 13447 38272 13453 38306
rect 13487 38305 13637 38306
rect 13487 38272 13525 38305
rect 13447 38271 13525 38272
rect 13559 38271 13597 38305
rect 13631 38271 13637 38305
rect 13447 38233 13637 38271
rect 13447 38199 13453 38233
rect 13487 38232 13637 38233
rect 13487 38199 13525 38232
rect 13447 38198 13525 38199
rect 13559 38198 13597 38232
rect 13631 38198 13637 38232
rect 13447 38160 13637 38198
rect 13447 38126 13453 38160
rect 13487 38159 13637 38160
rect 13487 38126 13525 38159
rect 13447 38125 13525 38126
rect 13559 38125 13597 38159
rect 13631 38125 13637 38159
rect 13447 38087 13637 38125
rect 13447 38053 13453 38087
rect 13487 38086 13637 38087
rect 13487 38053 13525 38086
rect 13447 38052 13525 38053
rect 13559 38052 13597 38086
rect 13631 38052 13637 38086
rect 13447 38014 13637 38052
rect 13447 37980 13453 38014
rect 13487 38013 13637 38014
rect 13487 37980 13525 38013
rect 13447 37979 13525 37980
rect 13559 37979 13597 38013
rect 13631 37979 13637 38013
rect 13447 37941 13637 37979
rect 13447 37907 13453 37941
rect 13487 37940 13637 37941
rect 13487 37907 13525 37940
rect 13447 37906 13525 37907
rect 13559 37906 13597 37940
rect 13631 37906 13637 37940
rect 13447 37868 13637 37906
rect 13447 37834 13453 37868
rect 13487 37867 13637 37868
rect 13487 37834 13525 37867
rect 13447 37833 13525 37834
rect 13559 37833 13597 37867
rect 13631 37833 13637 37867
rect 13447 37795 13637 37833
rect 13447 37761 13453 37795
rect 13487 37794 13637 37795
rect 13487 37761 13525 37794
rect 13447 37760 13525 37761
rect 13559 37760 13597 37794
rect 13631 37760 13637 37794
rect 13447 37722 13637 37760
rect 13447 37688 13453 37722
rect 13487 37721 13637 37722
rect 13487 37688 13525 37721
rect 13447 37687 13525 37688
rect 13559 37687 13597 37721
rect 13631 37687 13637 37721
rect 13447 37649 13637 37687
rect 13447 37615 13453 37649
rect 13487 37648 13637 37649
rect 13487 37615 13525 37648
rect 13447 37614 13525 37615
rect 13559 37614 13597 37648
rect 13631 37614 13637 37648
rect 13447 37576 13637 37614
rect 13447 37542 13453 37576
rect 13487 37575 13637 37576
rect 13487 37542 13525 37575
rect 13447 37541 13525 37542
rect 13559 37541 13597 37575
rect 13631 37541 13637 37575
rect 13447 37503 13637 37541
rect 13447 37469 13453 37503
rect 13487 37502 13637 37503
rect 13487 37469 13525 37502
rect 13447 37468 13525 37469
rect 13559 37468 13597 37502
rect 13631 37468 13637 37502
rect 13447 37430 13637 37468
rect 13447 37396 13453 37430
rect 13487 37429 13637 37430
rect 13487 37396 13525 37429
rect 13447 37395 13525 37396
rect 13559 37395 13597 37429
rect 13631 37395 13637 37429
rect 13447 37357 13637 37395
rect 13447 37323 13453 37357
rect 13487 37356 13637 37357
rect 13487 37323 13525 37356
rect 13447 37322 13525 37323
rect 13559 37322 13597 37356
rect 13631 37322 13637 37356
rect 13447 37284 13637 37322
rect 13447 37250 13453 37284
rect 13487 37283 13637 37284
rect 13487 37250 13525 37283
rect 13447 37249 13525 37250
rect 13559 37249 13597 37283
rect 13631 37249 13637 37283
rect 13447 37211 13637 37249
rect 13447 37177 13453 37211
rect 13487 37210 13637 37211
rect 13487 37177 13525 37210
rect 13447 37176 13525 37177
rect 13559 37176 13597 37210
rect 13631 37176 13637 37210
rect 13447 37138 13637 37176
rect 13447 37104 13453 37138
rect 13487 37137 13637 37138
rect 13487 37104 13525 37137
rect 13447 37103 13525 37104
rect 13559 37103 13597 37137
rect 13631 37103 13637 37137
rect 13447 37065 13637 37103
rect 13447 37031 13453 37065
rect 13487 37064 13637 37065
rect 13487 37031 13525 37064
rect 13447 37030 13525 37031
rect 13559 37030 13597 37064
rect 13631 37030 13637 37064
rect 13447 36992 13637 37030
rect 13447 36958 13453 36992
rect 13487 36991 13637 36992
rect 13487 36958 13525 36991
rect 13447 36957 13525 36958
rect 13559 36957 13597 36991
rect 13631 36957 13637 36991
rect 13447 36919 13637 36957
rect 13447 36885 13453 36919
rect 13487 36918 13637 36919
rect 13487 36885 13525 36918
rect 13447 36884 13525 36885
rect 13559 36884 13597 36918
rect 13631 36884 13637 36918
rect 13447 36846 13637 36884
rect 13447 36812 13453 36846
rect 13487 36845 13637 36846
rect 13487 36812 13525 36845
rect 13447 36811 13525 36812
rect 13559 36811 13597 36845
rect 13631 36811 13637 36845
rect 13447 36773 13637 36811
rect 13447 36739 13453 36773
rect 13487 36772 13637 36773
rect 13487 36739 13525 36772
rect 13447 36738 13525 36739
rect 13559 36738 13597 36772
rect 13631 36738 13637 36772
rect 13447 36700 13637 36738
rect 13447 36666 13453 36700
rect 13487 36699 13637 36700
rect 13487 36666 13525 36699
rect 13447 36665 13525 36666
rect 13559 36665 13597 36699
rect 13631 36665 13637 36699
rect 13447 36627 13637 36665
rect 13447 36593 13453 36627
rect 13487 36626 13637 36627
rect 13487 36593 13525 36626
rect 13447 36592 13525 36593
rect 13559 36592 13597 36626
rect 13631 36592 13637 36626
rect 13447 36554 13637 36592
rect 13447 36520 13453 36554
rect 13487 36553 13637 36554
rect 13487 36520 13525 36553
rect 13447 36519 13525 36520
rect 13559 36519 13597 36553
rect 13631 36519 13637 36553
rect 13447 36481 13637 36519
rect 13447 36447 13453 36481
rect 13487 36480 13637 36481
rect 13487 36447 13525 36480
rect 13447 36446 13525 36447
rect 13559 36446 13597 36480
rect 13631 36446 13637 36480
rect 13447 36408 13637 36446
rect 13447 36374 13453 36408
rect 13487 36407 13637 36408
rect 13487 36374 13525 36407
rect 13447 36373 13525 36374
rect 13559 36373 13597 36407
rect 13631 36373 13637 36407
rect 13447 36335 13637 36373
rect 13447 36301 13453 36335
rect 13487 36334 13637 36335
rect 13487 36301 13525 36334
rect 13447 36300 13525 36301
rect 13559 36300 13597 36334
rect 13631 36300 13637 36334
rect 13447 36262 13637 36300
rect 13447 36228 13453 36262
rect 13487 36261 13637 36262
rect 13487 36228 13525 36261
rect 13447 36227 13525 36228
rect 13559 36227 13597 36261
rect 13631 36227 13637 36261
rect 13447 36189 13637 36227
rect 13447 36155 13453 36189
rect 13487 36188 13637 36189
rect 13487 36155 13525 36188
rect 13447 36154 13525 36155
rect 13559 36154 13597 36188
rect 13631 36154 13637 36188
rect 13447 36116 13637 36154
rect 13447 36082 13453 36116
rect 13487 36115 13637 36116
rect 13487 36082 13525 36115
rect 13447 36081 13525 36082
rect 13559 36081 13597 36115
rect 13631 36081 13637 36115
rect 13447 36043 13637 36081
rect 13447 36009 13453 36043
rect 13487 36042 13637 36043
rect 13487 36009 13525 36042
rect 13447 36008 13525 36009
rect 13559 36008 13597 36042
rect 13631 36008 13637 36042
rect 13447 35970 13637 36008
rect 13447 35936 13453 35970
rect 13487 35969 13637 35970
rect 13487 35936 13525 35969
rect 13447 35935 13525 35936
rect 13559 35935 13597 35969
rect 13631 35935 13637 35969
rect 13447 35897 13637 35935
rect 13447 35863 13453 35897
rect 13487 35896 13637 35897
rect 13487 35863 13525 35896
rect 13447 35824 13525 35863
rect 13447 33198 13453 35824
rect 13631 33198 13637 35896
rect 13447 33186 13637 33198
tri 13447 33132 13501 33186 ne
rect 12991 31753 13181 32503
rect 12991 27903 12997 31753
rect 13175 27903 13181 31753
rect 12991 27153 13181 27903
rect 12991 23303 12997 27153
rect 13175 23303 13181 27153
rect 12991 22562 13181 23303
rect 12991 19360 12997 22562
rect 13175 19360 13181 22562
rect 13501 33118 13637 33186
rect 13501 33084 13507 33118
rect 13541 33084 13597 33118
rect 13631 33084 13637 33118
rect 13501 33046 13637 33084
rect 13501 33012 13507 33046
rect 13541 33012 13597 33046
rect 13631 33012 13637 33046
rect 13501 32974 13637 33012
rect 13501 32940 13507 32974
rect 13541 32940 13597 32974
rect 13631 32940 13637 32974
rect 13501 32902 13637 32940
rect 13501 32868 13507 32902
rect 13541 32868 13597 32902
rect 13631 32868 13637 32902
rect 13501 32830 13637 32868
rect 13501 32796 13507 32830
rect 13541 32796 13597 32830
rect 13631 32796 13637 32830
rect 13501 32758 13637 32796
rect 13501 32724 13507 32758
rect 13541 32724 13597 32758
rect 13631 32724 13637 32758
rect 13501 32686 13637 32724
rect 13501 32652 13507 32686
rect 13541 32652 13597 32686
rect 13631 32652 13637 32686
rect 13501 32614 13637 32652
rect 13501 32580 13507 32614
rect 13541 32580 13597 32614
rect 13631 32580 13637 32614
rect 13501 32542 13637 32580
rect 13501 32508 13507 32542
rect 13541 32508 13597 32542
rect 13631 32508 13637 32542
rect 13501 32470 13637 32508
rect 13501 32436 13507 32470
rect 13541 32436 13597 32470
rect 13631 32436 13637 32470
rect 13501 32398 13637 32436
rect 13501 32364 13507 32398
rect 13541 32364 13597 32398
rect 13631 32364 13637 32398
rect 13501 32326 13637 32364
rect 13501 32292 13507 32326
rect 13541 32292 13597 32326
rect 13631 32292 13637 32326
rect 13501 32254 13637 32292
rect 13501 32220 13507 32254
rect 13541 32220 13597 32254
rect 13631 32220 13637 32254
rect 13501 32182 13637 32220
rect 13501 32148 13507 32182
rect 13541 32148 13597 32182
rect 13631 32148 13637 32182
rect 13501 32110 13637 32148
rect 13501 32076 13507 32110
rect 13541 32076 13597 32110
rect 13631 32076 13637 32110
rect 13501 32038 13637 32076
rect 13501 32004 13507 32038
rect 13541 32004 13597 32038
rect 13631 32004 13637 32038
rect 13501 31966 13637 32004
rect 13501 31932 13507 31966
rect 13541 31932 13597 31966
rect 13631 31932 13637 31966
rect 13501 31894 13637 31932
rect 13501 31860 13507 31894
rect 13541 31860 13597 31894
rect 13631 31860 13637 31894
rect 13501 31822 13637 31860
rect 13501 31788 13507 31822
rect 13541 31788 13597 31822
rect 13631 31788 13637 31822
rect 13501 31750 13637 31788
rect 13501 31716 13507 31750
rect 13541 31716 13597 31750
rect 13631 31716 13637 31750
rect 13501 31678 13637 31716
rect 13501 31644 13507 31678
rect 13541 31644 13597 31678
rect 13631 31644 13637 31678
rect 13501 31606 13637 31644
rect 13501 31572 13507 31606
rect 13541 31572 13597 31606
rect 13631 31572 13637 31606
rect 13501 31534 13637 31572
rect 13501 31500 13507 31534
rect 13541 31500 13597 31534
rect 13631 31500 13637 31534
rect 13501 31462 13637 31500
rect 13501 31428 13507 31462
rect 13541 31428 13597 31462
rect 13631 31428 13637 31462
rect 13501 31390 13637 31428
rect 13501 31356 13507 31390
rect 13541 31356 13597 31390
rect 13631 31356 13637 31390
rect 13501 31318 13637 31356
rect 13501 31284 13507 31318
rect 13541 31284 13597 31318
rect 13631 31284 13637 31318
rect 13501 31246 13637 31284
rect 13501 31212 13507 31246
rect 13541 31212 13597 31246
rect 13631 31212 13637 31246
rect 13501 31174 13637 31212
rect 13501 31140 13507 31174
rect 13541 31140 13597 31174
rect 13631 31140 13637 31174
rect 13501 31102 13637 31140
rect 13501 31068 13507 31102
rect 13541 31068 13597 31102
rect 13631 31068 13637 31102
rect 13501 31030 13637 31068
rect 13501 30996 13507 31030
rect 13541 30996 13597 31030
rect 13631 30996 13637 31030
rect 13501 30958 13637 30996
rect 13501 30924 13507 30958
rect 13541 30924 13597 30958
rect 13631 30924 13637 30958
rect 13501 30886 13637 30924
rect 13501 30852 13507 30886
rect 13541 30852 13597 30886
rect 13631 30852 13637 30886
rect 13501 30814 13637 30852
rect 13501 30780 13507 30814
rect 13541 30780 13597 30814
rect 13631 30780 13637 30814
rect 13501 30742 13637 30780
rect 13501 30708 13507 30742
rect 13541 30708 13597 30742
rect 13631 30708 13637 30742
rect 13501 30670 13637 30708
rect 13501 30636 13507 30670
rect 13541 30636 13597 30670
rect 13631 30636 13637 30670
rect 13501 30598 13637 30636
rect 13501 30564 13507 30598
rect 13541 30564 13597 30598
rect 13631 30564 13637 30598
rect 13501 30526 13637 30564
rect 13501 30492 13507 30526
rect 13541 30492 13597 30526
rect 13631 30492 13637 30526
rect 13501 30454 13637 30492
rect 13501 30420 13507 30454
rect 13541 30420 13597 30454
rect 13631 30420 13637 30454
rect 13501 30382 13637 30420
rect 13501 30348 13507 30382
rect 13541 30348 13597 30382
rect 13631 30348 13637 30382
rect 13501 30310 13637 30348
rect 13501 30276 13507 30310
rect 13541 30276 13597 30310
rect 13631 30276 13637 30310
rect 13501 30238 13637 30276
rect 13501 30204 13507 30238
rect 13541 30204 13597 30238
rect 13631 30204 13637 30238
rect 13501 30166 13637 30204
rect 13501 30132 13507 30166
rect 13541 30132 13597 30166
rect 13631 30132 13637 30166
rect 13501 30094 13637 30132
rect 13501 30060 13507 30094
rect 13541 30060 13597 30094
rect 13631 30060 13637 30094
rect 13501 30022 13637 30060
rect 13501 29988 13507 30022
rect 13541 29988 13597 30022
rect 13631 29988 13637 30022
rect 13501 29950 13637 29988
rect 13501 29916 13507 29950
rect 13541 29916 13597 29950
rect 13631 29916 13637 29950
rect 13501 29878 13637 29916
rect 13501 29844 13507 29878
rect 13541 29844 13597 29878
rect 13631 29844 13637 29878
rect 13501 29806 13637 29844
rect 13501 29772 13507 29806
rect 13541 29772 13597 29806
rect 13631 29772 13637 29806
rect 13501 29734 13637 29772
rect 13501 29700 13507 29734
rect 13541 29700 13597 29734
rect 13631 29700 13637 29734
rect 13501 29662 13637 29700
rect 13501 29628 13507 29662
rect 13541 29628 13597 29662
rect 13631 29628 13637 29662
rect 13501 29590 13637 29628
rect 13501 29556 13507 29590
rect 13541 29556 13597 29590
rect 13631 29556 13637 29590
rect 13501 29518 13637 29556
rect 13501 29484 13507 29518
rect 13541 29484 13597 29518
rect 13631 29484 13637 29518
rect 13501 29446 13637 29484
rect 13501 29412 13507 29446
rect 13541 29412 13597 29446
rect 13631 29412 13637 29446
rect 13501 29374 13637 29412
rect 13501 29340 13507 29374
rect 13541 29340 13597 29374
rect 13631 29340 13637 29374
rect 13501 29302 13637 29340
rect 13501 29268 13507 29302
rect 13541 29268 13597 29302
rect 13631 29268 13637 29302
rect 13501 29230 13637 29268
rect 13501 29196 13507 29230
rect 13541 29196 13597 29230
rect 13631 29196 13637 29230
rect 13501 29158 13637 29196
rect 13501 29124 13507 29158
rect 13541 29124 13597 29158
rect 13631 29124 13637 29158
rect 13501 29086 13637 29124
rect 13501 29052 13507 29086
rect 13541 29052 13597 29086
rect 13631 29052 13637 29086
rect 13501 29014 13637 29052
rect 13501 28980 13507 29014
rect 13541 28980 13597 29014
rect 13631 28980 13637 29014
rect 13501 28942 13637 28980
rect 13501 28908 13507 28942
rect 13541 28908 13597 28942
rect 13631 28908 13637 28942
rect 13501 28870 13637 28908
rect 13501 28836 13507 28870
rect 13541 28836 13597 28870
rect 13631 28836 13637 28870
rect 13501 28798 13637 28836
rect 13501 28764 13507 28798
rect 13541 28764 13597 28798
rect 13631 28764 13637 28798
rect 13501 28726 13637 28764
rect 13501 28692 13507 28726
rect 13541 28692 13597 28726
rect 13631 28692 13637 28726
rect 13501 28654 13637 28692
rect 13501 28620 13507 28654
rect 13541 28620 13597 28654
rect 13631 28620 13637 28654
rect 13501 28582 13637 28620
rect 13501 28548 13507 28582
rect 13541 28548 13597 28582
rect 13631 28548 13637 28582
rect 13501 28510 13637 28548
rect 13501 28476 13507 28510
rect 13541 28476 13597 28510
rect 13631 28476 13637 28510
rect 13501 28438 13637 28476
rect 13501 28404 13507 28438
rect 13541 28404 13597 28438
rect 13631 28404 13637 28438
rect 13501 28366 13637 28404
rect 13501 28332 13507 28366
rect 13541 28332 13597 28366
rect 13631 28332 13637 28366
rect 13501 28294 13637 28332
rect 13501 28260 13507 28294
rect 13541 28260 13597 28294
rect 13631 28260 13637 28294
rect 13501 28222 13637 28260
rect 13501 28188 13507 28222
rect 13541 28188 13597 28222
rect 13631 28188 13637 28222
rect 13501 28150 13637 28188
rect 13501 28116 13507 28150
rect 13541 28116 13597 28150
rect 13631 28116 13637 28150
rect 13501 28078 13637 28116
rect 13501 28044 13507 28078
rect 13541 28044 13597 28078
rect 13631 28044 13637 28078
rect 13501 28006 13637 28044
rect 13501 27972 13507 28006
rect 13541 27972 13597 28006
rect 13631 27972 13637 28006
rect 13501 27934 13637 27972
rect 13501 27900 13507 27934
rect 13541 27900 13597 27934
rect 13631 27900 13637 27934
rect 13501 27862 13637 27900
rect 13501 27828 13507 27862
rect 13541 27828 13597 27862
rect 13631 27828 13637 27862
rect 13501 27790 13637 27828
rect 13501 27756 13507 27790
rect 13541 27756 13597 27790
rect 13631 27756 13637 27790
rect 13501 27718 13637 27756
rect 13501 27684 13507 27718
rect 13541 27684 13597 27718
rect 13631 27684 13637 27718
rect 13501 27646 13637 27684
rect 13501 27612 13507 27646
rect 13541 27612 13597 27646
rect 13631 27612 13637 27646
rect 13501 27574 13637 27612
rect 13501 27540 13507 27574
rect 13541 27540 13597 27574
rect 13631 27540 13637 27574
rect 13501 27502 13637 27540
rect 13501 27468 13507 27502
rect 13541 27468 13597 27502
rect 13631 27468 13637 27502
rect 13501 27430 13637 27468
rect 13501 27396 13507 27430
rect 13541 27396 13597 27430
rect 13631 27396 13637 27430
rect 13501 27358 13637 27396
rect 13501 27324 13507 27358
rect 13541 27324 13597 27358
rect 13631 27324 13637 27358
rect 13501 27286 13637 27324
rect 13501 27252 13507 27286
rect 13541 27252 13597 27286
rect 13631 27252 13637 27286
rect 13501 27214 13637 27252
rect 13501 27180 13507 27214
rect 13541 27180 13597 27214
rect 13631 27180 13637 27214
rect 13501 27142 13637 27180
rect 13501 27108 13507 27142
rect 13541 27108 13597 27142
rect 13631 27108 13637 27142
rect 13501 27070 13637 27108
rect 13501 27036 13507 27070
rect 13541 27036 13597 27070
rect 13631 27036 13637 27070
rect 13501 26998 13637 27036
rect 13501 26964 13507 26998
rect 13541 26964 13597 26998
rect 13631 26964 13637 26998
rect 13501 26926 13637 26964
rect 13501 26892 13507 26926
rect 13541 26892 13597 26926
rect 13631 26892 13637 26926
rect 13501 26854 13637 26892
rect 13501 26820 13507 26854
rect 13541 26820 13597 26854
rect 13631 26820 13637 26854
rect 13501 26782 13637 26820
rect 13501 26748 13507 26782
rect 13541 26748 13597 26782
rect 13631 26748 13637 26782
rect 13501 26710 13637 26748
rect 13501 26676 13507 26710
rect 13541 26676 13597 26710
rect 13631 26676 13637 26710
rect 13501 26638 13637 26676
rect 13501 26604 13507 26638
rect 13541 26604 13597 26638
rect 13631 26604 13637 26638
rect 13501 26566 13637 26604
rect 13501 26532 13507 26566
rect 13541 26532 13597 26566
rect 13631 26532 13637 26566
rect 13501 26494 13637 26532
rect 13501 26460 13507 26494
rect 13541 26460 13597 26494
rect 13631 26460 13637 26494
rect 13501 26422 13637 26460
rect 13501 26388 13507 26422
rect 13541 26388 13597 26422
rect 13631 26388 13637 26422
rect 13501 26350 13637 26388
rect 13501 26316 13507 26350
rect 13541 26316 13597 26350
rect 13631 26316 13637 26350
rect 13501 26278 13637 26316
rect 13501 26244 13507 26278
rect 13541 26244 13597 26278
rect 13631 26244 13637 26278
rect 13501 26206 13637 26244
rect 13501 26172 13507 26206
rect 13541 26172 13597 26206
rect 13631 26172 13637 26206
rect 13501 26134 13637 26172
rect 13501 26100 13507 26134
rect 13541 26100 13597 26134
rect 13631 26100 13637 26134
rect 13501 26062 13637 26100
rect 13501 26028 13507 26062
rect 13541 26028 13597 26062
rect 13631 26028 13637 26062
rect 13501 25990 13637 26028
rect 13501 25956 13507 25990
rect 13541 25956 13597 25990
rect 13631 25956 13637 25990
rect 13501 25918 13637 25956
rect 13501 25884 13507 25918
rect 13541 25884 13597 25918
rect 13631 25884 13637 25918
rect 13501 25846 13637 25884
rect 13501 25812 13507 25846
rect 13541 25812 13597 25846
rect 13631 25812 13637 25846
rect 13501 25774 13637 25812
rect 13501 25740 13507 25774
rect 13541 25740 13597 25774
rect 13631 25740 13637 25774
rect 13501 25702 13637 25740
rect 13501 25668 13507 25702
rect 13541 25668 13597 25702
rect 13631 25668 13637 25702
rect 13501 25630 13637 25668
rect 13501 25596 13507 25630
rect 13541 25596 13597 25630
rect 13631 25596 13637 25630
rect 13501 25558 13637 25596
rect 13501 25524 13507 25558
rect 13541 25524 13597 25558
rect 13631 25524 13637 25558
rect 13501 25486 13637 25524
rect 13501 25452 13507 25486
rect 13541 25452 13597 25486
rect 13631 25452 13637 25486
rect 13501 25413 13637 25452
rect 13501 25379 13507 25413
rect 13541 25379 13597 25413
rect 13631 25379 13637 25413
rect 13501 25340 13637 25379
rect 13501 25306 13507 25340
rect 13541 25306 13597 25340
rect 13631 25306 13637 25340
rect 13501 25267 13637 25306
rect 13501 25233 13507 25267
rect 13541 25233 13597 25267
rect 13631 25233 13637 25267
rect 13501 25194 13637 25233
rect 13501 25160 13507 25194
rect 13541 25160 13597 25194
rect 13631 25160 13637 25194
rect 13501 25121 13637 25160
rect 13501 25087 13507 25121
rect 13541 25087 13597 25121
rect 13631 25087 13637 25121
rect 13501 25048 13637 25087
rect 13501 25014 13507 25048
rect 13541 25014 13597 25048
rect 13631 25014 13637 25048
rect 13501 24975 13637 25014
rect 13501 24941 13507 24975
rect 13541 24941 13597 24975
rect 13631 24941 13637 24975
rect 13501 24902 13637 24941
rect 13501 24868 13507 24902
rect 13541 24868 13597 24902
rect 13631 24868 13637 24902
rect 13501 24829 13637 24868
rect 13501 24795 13507 24829
rect 13541 24795 13597 24829
rect 13631 24795 13637 24829
rect 13501 24756 13637 24795
rect 13501 24722 13507 24756
rect 13541 24722 13597 24756
rect 13631 24722 13637 24756
rect 13501 24683 13637 24722
rect 13501 24649 13507 24683
rect 13541 24649 13597 24683
rect 13631 24649 13637 24683
rect 13501 24610 13637 24649
rect 13501 24576 13507 24610
rect 13541 24576 13597 24610
rect 13631 24576 13637 24610
rect 13501 24537 13637 24576
rect 13501 24503 13507 24537
rect 13541 24503 13597 24537
rect 13631 24503 13637 24537
rect 13501 24464 13637 24503
rect 13501 24430 13507 24464
rect 13541 24430 13597 24464
rect 13631 24430 13637 24464
rect 13501 24391 13637 24430
rect 13501 24357 13507 24391
rect 13541 24357 13597 24391
rect 13631 24357 13637 24391
rect 13501 24318 13637 24357
rect 13501 24284 13507 24318
rect 13541 24284 13597 24318
rect 13631 24284 13637 24318
rect 13501 24245 13637 24284
rect 13501 24211 13507 24245
rect 13541 24211 13597 24245
rect 13631 24211 13637 24245
rect 13501 24172 13637 24211
rect 13501 24138 13507 24172
rect 13541 24138 13597 24172
rect 13631 24138 13637 24172
rect 13501 24099 13637 24138
rect 13501 24065 13507 24099
rect 13541 24065 13597 24099
rect 13631 24065 13637 24099
rect 13501 24026 13637 24065
rect 13501 23992 13507 24026
rect 13541 23992 13597 24026
rect 13631 23992 13637 24026
rect 13501 23953 13637 23992
rect 13501 23919 13507 23953
rect 13541 23919 13597 23953
rect 13631 23919 13637 23953
rect 13501 23880 13637 23919
rect 13501 23846 13507 23880
rect 13541 23846 13597 23880
rect 13631 23846 13637 23880
rect 13501 23807 13637 23846
rect 13501 23773 13507 23807
rect 13541 23773 13597 23807
rect 13631 23773 13637 23807
rect 13501 23734 13637 23773
rect 13501 23700 13507 23734
rect 13541 23700 13597 23734
rect 13631 23700 13637 23734
rect 13501 23661 13637 23700
rect 13501 23627 13507 23661
rect 13541 23627 13597 23661
rect 13631 23627 13637 23661
rect 13501 23588 13637 23627
rect 13501 23554 13507 23588
rect 13541 23554 13597 23588
rect 13631 23554 13637 23588
rect 13501 23515 13637 23554
rect 13501 23481 13507 23515
rect 13541 23481 13597 23515
rect 13631 23481 13637 23515
rect 13501 23442 13637 23481
rect 13501 23408 13507 23442
rect 13541 23408 13597 23442
rect 13631 23408 13637 23442
rect 13501 23369 13637 23408
rect 13501 23335 13507 23369
rect 13541 23335 13597 23369
rect 13631 23335 13637 23369
rect 13501 23296 13637 23335
rect 13501 23262 13507 23296
rect 13541 23262 13597 23296
rect 13631 23262 13637 23296
rect 13501 23223 13637 23262
rect 13501 23189 13507 23223
rect 13541 23189 13597 23223
rect 13631 23189 13637 23223
rect 13501 23150 13637 23189
rect 13501 23116 13507 23150
rect 13541 23116 13597 23150
rect 13631 23116 13637 23150
rect 13501 23077 13637 23116
rect 13501 23043 13507 23077
rect 13541 23043 13597 23077
rect 13631 23043 13637 23077
rect 13501 23004 13637 23043
rect 13501 22970 13507 23004
rect 13541 22970 13597 23004
rect 13631 22970 13637 23004
rect 13501 22931 13637 22970
rect 13501 22897 13507 22931
rect 13541 22897 13597 22931
rect 13631 22897 13637 22931
rect 13501 22858 13637 22897
rect 13501 22824 13507 22858
rect 13541 22824 13597 22858
rect 13631 22824 13637 22858
rect 13501 22785 13637 22824
rect 13501 22751 13507 22785
rect 13541 22751 13597 22785
rect 13631 22751 13637 22785
rect 13501 22712 13637 22751
rect 13501 22678 13507 22712
rect 13541 22678 13597 22712
rect 13631 22678 13637 22712
rect 13501 22639 13637 22678
rect 13501 22605 13507 22639
rect 13541 22605 13597 22639
rect 13631 22605 13637 22639
rect 13501 22566 13637 22605
rect 13501 22532 13507 22566
rect 13541 22532 13597 22566
rect 13631 22532 13637 22566
rect 13501 22493 13637 22532
rect 13501 22459 13507 22493
rect 13541 22459 13597 22493
rect 13631 22459 13637 22493
rect 13501 22420 13637 22459
rect 13501 22386 13507 22420
rect 13541 22386 13597 22420
rect 13631 22386 13637 22420
rect 13501 22347 13637 22386
rect 13501 22313 13507 22347
rect 13541 22313 13597 22347
rect 13631 22313 13637 22347
rect 13501 22274 13637 22313
rect 13501 22240 13507 22274
rect 13541 22240 13597 22274
rect 13631 22240 13637 22274
rect 13501 22201 13637 22240
rect 13501 22167 13507 22201
rect 13541 22167 13597 22201
rect 13631 22167 13637 22201
rect 13501 22128 13637 22167
rect 13501 22094 13507 22128
rect 13541 22094 13597 22128
rect 13631 22094 13637 22128
rect 13501 22055 13637 22094
rect 13501 22021 13507 22055
rect 13541 22021 13597 22055
rect 13631 22021 13637 22055
rect 13501 21982 13637 22021
rect 13501 21948 13507 21982
rect 13541 21948 13597 21982
rect 13631 21948 13637 21982
rect 13501 21909 13637 21948
rect 13501 21875 13507 21909
rect 13541 21875 13597 21909
rect 13631 21875 13637 21909
rect 13501 21836 13637 21875
rect 13501 21802 13507 21836
rect 13541 21802 13597 21836
rect 13631 21802 13637 21836
rect 13501 21763 13637 21802
rect 13501 21729 13507 21763
rect 13541 21729 13597 21763
rect 13631 21729 13637 21763
rect 13501 21690 13637 21729
rect 13501 21656 13507 21690
rect 13541 21656 13597 21690
rect 13631 21656 13637 21690
rect 13501 21617 13637 21656
rect 13501 21583 13507 21617
rect 13541 21583 13597 21617
rect 13631 21583 13637 21617
rect 13501 21544 13637 21583
rect 13501 21510 13507 21544
rect 13541 21510 13597 21544
rect 13631 21510 13637 21544
rect 13501 21471 13637 21510
rect 13501 21437 13507 21471
rect 13541 21437 13597 21471
rect 13631 21437 13637 21471
rect 13501 21398 13637 21437
rect 13501 21364 13507 21398
rect 13541 21364 13597 21398
rect 13631 21364 13637 21398
rect 13501 21325 13637 21364
rect 13501 21291 13507 21325
rect 13541 21291 13597 21325
rect 13631 21291 13637 21325
rect 13501 21252 13637 21291
rect 13501 21218 13507 21252
rect 13541 21218 13597 21252
rect 13631 21218 13637 21252
rect 13501 21179 13637 21218
rect 13501 21145 13507 21179
rect 13541 21145 13597 21179
rect 13631 21145 13637 21179
rect 13501 21106 13637 21145
rect 13501 21072 13507 21106
rect 13541 21072 13597 21106
rect 13631 21072 13637 21106
rect 13501 21033 13637 21072
rect 13501 20999 13507 21033
rect 13541 20999 13597 21033
rect 13631 20999 13637 21033
rect 13501 20960 13637 20999
rect 13501 20926 13507 20960
rect 13541 20926 13597 20960
rect 13631 20926 13637 20960
rect 13501 20887 13637 20926
rect 13501 20853 13507 20887
rect 13541 20853 13597 20887
rect 13631 20853 13637 20887
rect 13501 20814 13637 20853
rect 13501 20780 13507 20814
rect 13541 20780 13597 20814
rect 13631 20780 13637 20814
rect 13501 20741 13637 20780
rect 13501 20707 13507 20741
rect 13541 20707 13597 20741
rect 13631 20707 13637 20741
rect 13501 20668 13637 20707
rect 13501 20634 13507 20668
rect 13541 20634 13597 20668
rect 13631 20634 13637 20668
rect 13501 20595 13637 20634
rect 13501 20561 13507 20595
rect 13541 20561 13597 20595
rect 13631 20561 13637 20595
rect 13501 20522 13637 20561
rect 13501 20488 13507 20522
rect 13541 20488 13597 20522
rect 13631 20488 13637 20522
rect 13501 20449 13637 20488
rect 13501 20415 13507 20449
rect 13541 20415 13597 20449
rect 13631 20415 13637 20449
rect 13501 20376 13637 20415
rect 13501 20342 13507 20376
rect 13541 20342 13597 20376
rect 13631 20342 13637 20376
rect 12991 19321 13181 19360
rect 12991 19287 12997 19321
rect 13031 19287 13069 19321
rect 13103 19287 13141 19321
rect 13175 19287 13181 19321
rect 12991 19248 13181 19287
rect 12991 19214 12997 19248
rect 13031 19214 13069 19248
rect 13103 19214 13141 19248
rect 13175 19214 13181 19248
rect 12991 19175 13181 19214
rect 12991 19141 12997 19175
rect 13031 19141 13069 19175
rect 13103 19141 13141 19175
rect 13175 19141 13181 19175
rect 12991 19102 13181 19141
rect 12991 19068 12997 19102
rect 13031 19068 13069 19102
rect 13103 19068 13141 19102
rect 13175 19068 13181 19102
rect 12991 19029 13181 19068
rect 12991 18995 12997 19029
rect 13031 18995 13069 19029
rect 13103 18995 13141 19029
rect 13175 18995 13181 19029
rect 12991 18956 13181 18995
rect 12991 18922 12997 18956
rect 13031 18922 13069 18956
rect 13103 18922 13141 18956
rect 13175 18922 13181 18956
rect 12991 18883 13181 18922
rect 12991 18849 12997 18883
rect 13031 18849 13069 18883
rect 13103 18849 13141 18883
rect 13175 18849 13181 18883
rect 12991 18810 13181 18849
rect 12991 18776 12997 18810
rect 13031 18776 13069 18810
rect 13103 18776 13141 18810
rect 13175 18776 13181 18810
rect 12991 18737 13181 18776
rect 12991 18703 12997 18737
rect 13031 18703 13069 18737
rect 13103 18703 13141 18737
rect 13175 18703 13181 18737
rect 12991 17953 13181 18703
rect 12991 14103 12997 17953
rect 13175 14103 13181 17953
rect 12991 13362 13181 14103
rect 12991 10160 12997 13362
rect 13175 10160 13181 13362
rect 12991 10121 13181 10160
rect 12991 10087 12997 10121
rect 13031 10087 13069 10121
rect 13103 10087 13141 10121
rect 13175 10087 13181 10121
rect 12991 10048 13181 10087
rect 12991 10014 12997 10048
rect 13031 10014 13069 10048
rect 13103 10014 13141 10048
rect 13175 10014 13181 10048
rect 12991 9975 13181 10014
rect 12991 9941 12997 9975
rect 13031 9941 13069 9975
rect 13103 9941 13141 9975
rect 13175 9941 13181 9975
rect 12991 9902 13181 9941
rect 12991 9868 12997 9902
rect 13031 9868 13069 9902
rect 13103 9868 13141 9902
rect 13175 9868 13181 9902
rect 12991 9829 13181 9868
rect 12991 9795 12997 9829
rect 13031 9795 13069 9829
rect 13103 9795 13141 9829
rect 13175 9795 13181 9829
rect 12991 9756 13181 9795
rect 12991 9722 12997 9756
rect 13031 9722 13069 9756
rect 13103 9722 13141 9756
rect 13175 9722 13181 9756
rect 12991 9683 13181 9722
rect 12991 9649 12997 9683
rect 13031 9649 13069 9683
rect 13103 9649 13141 9683
rect 13175 9649 13181 9683
rect 12991 9610 13181 9649
rect 12991 9576 12997 9610
rect 13031 9576 13069 9610
rect 13103 9576 13141 9610
rect 13175 9576 13181 9610
rect 12991 9537 13181 9576
rect 12991 9503 12997 9537
rect 13031 9503 13069 9537
rect 13103 9503 13141 9537
rect 13175 9503 13181 9537
rect 12991 9491 13181 9503
tri 13447 20275 13501 20329 se
rect 13501 20275 13637 20342
rect 13447 20263 13637 20275
rect 13447 20229 13453 20263
rect 13487 20229 13525 20263
rect 13559 20229 13597 20263
rect 13631 20229 13637 20263
rect 13447 20190 13637 20229
rect 13447 20156 13453 20190
rect 13487 20156 13525 20190
rect 13559 20156 13597 20190
rect 13631 20156 13637 20190
rect 13447 20117 13637 20156
rect 13447 20083 13453 20117
rect 13487 20083 13525 20117
rect 13559 20083 13597 20117
rect 13631 20083 13637 20117
rect 13447 20044 13637 20083
rect 13447 20010 13453 20044
rect 13487 20010 13525 20044
rect 13559 20010 13597 20044
rect 13631 20010 13637 20044
rect 13447 19971 13637 20010
rect 13447 19937 13453 19971
rect 13487 19937 13525 19971
rect 13559 19937 13597 19971
rect 13631 19937 13637 19971
rect 13447 19898 13637 19937
rect 13447 19864 13453 19898
rect 13487 19864 13525 19898
rect 13559 19864 13597 19898
rect 13631 19864 13637 19898
rect 13447 19825 13637 19864
rect 13447 19791 13453 19825
rect 13487 19791 13525 19825
rect 13559 19791 13597 19825
rect 13631 19791 13637 19825
rect 13447 19752 13637 19791
rect 13447 19718 13453 19752
rect 13487 19718 13525 19752
rect 13559 19718 13597 19752
rect 13631 19718 13637 19752
rect 13447 19679 13637 19718
rect 13447 19645 13453 19679
rect 13487 19645 13525 19679
rect 13559 19645 13597 19679
rect 13631 19645 13637 19679
rect 13447 19606 13637 19645
rect 13447 19572 13453 19606
rect 13487 19572 13525 19606
rect 13559 19572 13597 19606
rect 13631 19572 13637 19606
rect 13447 19533 13637 19572
rect 13447 19499 13453 19533
rect 13487 19499 13525 19533
rect 13559 19499 13597 19533
rect 13631 19499 13637 19533
rect 13447 19460 13637 19499
rect 13447 19426 13453 19460
rect 13487 19426 13525 19460
rect 13559 19426 13597 19460
rect 13631 19426 13637 19460
rect 13447 19387 13637 19426
rect 13447 19353 13453 19387
rect 13487 19353 13525 19387
rect 13559 19353 13597 19387
rect 13631 19353 13637 19387
rect 13447 19314 13637 19353
rect 13447 19280 13453 19314
rect 13487 19280 13525 19314
rect 13559 19280 13597 19314
rect 13631 19280 13637 19314
rect 13447 19241 13637 19280
rect 13447 19207 13453 19241
rect 13487 19207 13525 19241
rect 13559 19207 13597 19241
rect 13631 19207 13637 19241
rect 13447 19168 13637 19207
rect 13447 19134 13453 19168
rect 13487 19134 13525 19168
rect 13559 19134 13597 19168
rect 13631 19134 13637 19168
rect 13447 19095 13637 19134
rect 13447 19061 13453 19095
rect 13487 19061 13525 19095
rect 13559 19061 13597 19095
rect 13631 19061 13637 19095
rect 13447 19022 13637 19061
rect 13447 18988 13453 19022
rect 13487 18988 13525 19022
rect 13559 18988 13597 19022
rect 13631 18988 13637 19022
rect 13447 18949 13637 18988
rect 13447 18915 13453 18949
rect 13487 18915 13525 18949
rect 13559 18915 13597 18949
rect 13631 18915 13637 18949
rect 13447 18876 13637 18915
rect 13447 18842 13453 18876
rect 13487 18842 13525 18876
rect 13559 18842 13597 18876
rect 13631 18842 13637 18876
rect 13447 18803 13637 18842
rect 13447 18769 13453 18803
rect 13487 18769 13525 18803
rect 13559 18769 13597 18803
rect 13631 18769 13637 18803
rect 13447 18730 13637 18769
rect 13447 18696 13453 18730
rect 13487 18696 13525 18730
rect 13559 18696 13597 18730
rect 13631 18696 13637 18730
rect 13447 18657 13637 18696
rect 13447 18623 13453 18657
rect 13487 18623 13525 18657
rect 13559 18623 13597 18657
rect 13631 18623 13637 18657
rect 13447 18584 13637 18623
rect 13447 18550 13453 18584
rect 13487 18550 13525 18584
rect 13559 18550 13597 18584
rect 13631 18550 13637 18584
rect 13447 18511 13637 18550
rect 13447 18477 13453 18511
rect 13487 18477 13525 18511
rect 13559 18477 13597 18511
rect 13631 18477 13637 18511
rect 13447 18438 13637 18477
rect 13447 18404 13453 18438
rect 13487 18404 13525 18438
rect 13559 18404 13597 18438
rect 13631 18404 13637 18438
rect 13447 18365 13637 18404
rect 13447 18331 13453 18365
rect 13487 18331 13525 18365
rect 13559 18331 13597 18365
rect 13631 18331 13637 18365
rect 13447 18292 13637 18331
rect 13447 18258 13453 18292
rect 13487 18258 13525 18292
rect 13559 18258 13597 18292
rect 13631 18258 13637 18292
rect 13447 18219 13637 18258
rect 13447 18185 13453 18219
rect 13487 18185 13525 18219
rect 13559 18185 13597 18219
rect 13631 18185 13637 18219
rect 13447 18146 13637 18185
rect 13447 18112 13453 18146
rect 13487 18112 13525 18146
rect 13559 18112 13597 18146
rect 13631 18112 13637 18146
rect 13447 18073 13637 18112
rect 13447 18039 13453 18073
rect 13487 18039 13525 18073
rect 13559 18039 13597 18073
rect 13631 18039 13637 18073
rect 13447 18000 13637 18039
rect 13447 17966 13453 18000
rect 13487 17966 13525 18000
rect 13559 17966 13597 18000
rect 13631 17966 13637 18000
rect 13447 17927 13637 17966
rect 13447 17893 13453 17927
rect 13487 17893 13525 17927
rect 13559 17893 13597 17927
rect 13631 17893 13637 17927
rect 13447 17854 13637 17893
rect 13447 17820 13453 17854
rect 13487 17820 13525 17854
rect 13559 17820 13597 17854
rect 13631 17820 13637 17854
rect 13447 17781 13637 17820
rect 13447 17747 13453 17781
rect 13487 17747 13525 17781
rect 13559 17747 13597 17781
rect 13631 17747 13637 17781
rect 13447 17708 13637 17747
rect 13447 17674 13453 17708
rect 13487 17674 13525 17708
rect 13559 17674 13597 17708
rect 13631 17674 13637 17708
rect 13447 17635 13637 17674
rect 13447 17601 13453 17635
rect 13487 17601 13525 17635
rect 13559 17601 13597 17635
rect 13631 17601 13637 17635
rect 13447 17562 13637 17601
rect 13447 17528 13453 17562
rect 13487 17528 13525 17562
rect 13559 17528 13597 17562
rect 13631 17528 13637 17562
rect 13447 17489 13637 17528
rect 13447 17455 13453 17489
rect 13487 17455 13525 17489
rect 13559 17455 13597 17489
rect 13631 17455 13637 17489
rect 13447 17416 13637 17455
rect 13447 17382 13453 17416
rect 13487 17382 13525 17416
rect 13559 17382 13597 17416
rect 13631 17382 13637 17416
rect 13447 17343 13637 17382
rect 13447 17309 13453 17343
rect 13487 17309 13525 17343
rect 13559 17309 13597 17343
rect 13631 17309 13637 17343
rect 13447 17270 13637 17309
rect 13447 17236 13453 17270
rect 13487 17236 13525 17270
rect 13559 17236 13597 17270
rect 13631 17236 13637 17270
rect 13447 17197 13637 17236
rect 13447 17163 13453 17197
rect 13487 17163 13525 17197
rect 13559 17163 13597 17197
rect 13631 17163 13637 17197
rect 13447 17124 13637 17163
rect 13447 17090 13453 17124
rect 13487 17090 13525 17124
rect 13559 17090 13597 17124
rect 13631 17090 13637 17124
rect 13447 17051 13637 17090
rect 13447 17017 13453 17051
rect 13487 17017 13525 17051
rect 13559 17017 13597 17051
rect 13631 17017 13637 17051
rect 13447 16978 13637 17017
rect 13447 16944 13453 16978
rect 13487 16944 13525 16978
rect 13559 16944 13597 16978
rect 13631 16944 13637 16978
rect 13447 16905 13637 16944
rect 13447 16871 13453 16905
rect 13487 16871 13525 16905
rect 13559 16871 13597 16905
rect 13631 16871 13637 16905
rect 13447 16832 13637 16871
rect 13447 16798 13453 16832
rect 13487 16798 13525 16832
rect 13559 16798 13597 16832
rect 13631 16798 13637 16832
rect 13447 16759 13637 16798
rect 13447 16725 13453 16759
rect 13487 16725 13525 16759
rect 13559 16725 13597 16759
rect 13631 16725 13637 16759
rect 13447 16686 13637 16725
rect 2611 9436 2617 9470
rect 2651 9436 2657 9470
rect 2611 9397 2657 9436
tri 2657 9397 2716 9456 sw
rect 2611 9363 2617 9397
rect 2651 9391 12899 9397
rect 2651 9363 2697 9391
rect 2611 9357 2697 9363
rect 2731 9357 2770 9391
rect 2804 9357 2843 9391
rect 2877 9357 2916 9391
rect 2950 9357 2989 9391
rect 3023 9357 3061 9391
rect 3095 9357 3133 9391
rect 3167 9357 3205 9391
rect 3239 9357 3277 9391
rect 3311 9357 3349 9391
rect 3383 9357 3421 9391
rect 3455 9357 3493 9391
rect 3527 9357 3565 9391
rect 3599 9357 3637 9391
rect 3671 9357 3709 9391
rect 3743 9357 3781 9391
rect 3815 9357 3853 9391
rect 3887 9357 3925 9391
rect 3959 9357 3997 9391
rect 4031 9357 4069 9391
rect 4103 9357 4141 9391
rect 4175 9357 4213 9391
rect 4247 9357 4285 9391
rect 4319 9357 4357 9391
rect 4391 9357 4429 9391
rect 4463 9357 4501 9391
rect 4535 9357 4573 9391
rect 4607 9357 4645 9391
rect 4679 9357 4717 9391
rect 4751 9357 4789 9391
rect 4823 9357 4861 9391
rect 4895 9357 4933 9391
rect 4967 9357 5005 9391
rect 5039 9357 5077 9391
rect 5111 9357 5149 9391
rect 5183 9357 5221 9391
rect 5255 9357 5293 9391
rect 5327 9357 5365 9391
rect 5399 9357 5437 9391
rect 5471 9357 5509 9391
rect 5543 9357 5581 9391
rect 5615 9357 5653 9391
rect 5687 9357 5725 9391
rect 5759 9357 5797 9391
rect 5831 9357 5869 9391
rect 5903 9357 5941 9391
rect 5975 9357 6013 9391
rect 6047 9357 6085 9391
rect 6119 9357 6157 9391
rect 6191 9357 6229 9391
rect 6263 9357 6301 9391
rect 6335 9357 6373 9391
rect 6407 9357 6445 9391
rect 6479 9357 6517 9391
rect 6551 9357 6589 9391
rect 6623 9357 6661 9391
rect 6695 9357 6733 9391
rect 6767 9357 6805 9391
rect 6839 9357 6877 9391
rect 6911 9357 6949 9391
rect 6983 9357 7021 9391
rect 7055 9357 7093 9391
rect 7127 9357 7165 9391
rect 7199 9357 7237 9391
rect 7271 9357 7309 9391
rect 7343 9357 7381 9391
rect 7415 9357 7453 9391
rect 7487 9357 7525 9391
rect 7559 9357 7597 9391
rect 7631 9357 7669 9391
rect 7703 9357 7741 9391
rect 7775 9357 7813 9391
rect 7847 9357 7885 9391
rect 7919 9357 7957 9391
rect 7991 9357 8029 9391
rect 8063 9357 8101 9391
rect 8135 9357 8173 9391
rect 8207 9357 8245 9391
rect 8279 9357 8317 9391
rect 8351 9357 8389 9391
rect 8423 9357 8461 9391
rect 8495 9357 8533 9391
rect 8567 9357 8605 9391
rect 8639 9357 8677 9391
rect 8711 9357 8749 9391
rect 8783 9357 8821 9391
rect 8855 9357 8893 9391
rect 8927 9357 8965 9391
rect 8999 9357 9037 9391
rect 9071 9357 9109 9391
rect 9143 9357 9181 9391
rect 9215 9357 9253 9391
rect 9287 9357 9325 9391
rect 9359 9357 9397 9391
rect 9431 9357 9469 9391
rect 9503 9357 9541 9391
rect 9575 9357 9613 9391
rect 9647 9357 9685 9391
rect 9719 9357 9757 9391
rect 9791 9357 9829 9391
rect 9863 9357 9901 9391
rect 9935 9357 9973 9391
rect 10007 9357 10045 9391
rect 10079 9357 10117 9391
rect 10151 9357 10189 9391
rect 10223 9357 10261 9391
rect 10295 9357 10333 9391
rect 10367 9357 10405 9391
rect 10439 9357 10477 9391
rect 10511 9357 10549 9391
rect 10583 9357 10621 9391
rect 10655 9357 10693 9391
rect 10727 9357 10765 9391
rect 10799 9357 10837 9391
rect 10871 9357 10909 9391
rect 10943 9357 10981 9391
rect 11015 9357 11053 9391
rect 11087 9357 11125 9391
rect 11159 9357 11197 9391
rect 11231 9357 11269 9391
rect 11303 9357 11341 9391
rect 11375 9357 11413 9391
rect 11447 9357 11485 9391
rect 11519 9357 11557 9391
rect 11591 9357 11629 9391
rect 11663 9357 11701 9391
rect 11735 9357 11773 9391
rect 11807 9357 11845 9391
rect 11879 9357 11917 9391
rect 11951 9357 11989 9391
rect 12023 9357 12061 9391
rect 12095 9357 12133 9391
rect 12167 9357 12205 9391
rect 12239 9357 12277 9391
rect 12311 9357 12349 9391
rect 12383 9357 12421 9391
rect 12455 9357 12493 9391
rect 12527 9357 12565 9391
rect 12599 9357 12637 9391
rect 12671 9357 12709 9391
rect 12743 9357 12781 9391
rect 12815 9357 12853 9391
rect 12887 9357 12899 9391
rect 2215 9344 2233 9352
rect 2285 9344 2335 9352
rect 2215 9310 2221 9344
rect 2285 9310 2293 9344
rect 2327 9310 2335 9344
rect 2387 9351 2405 9352
tri 2405 9351 2408 9354 sw
rect 2611 9351 12899 9357
rect 2387 9343 2408 9351
rect 2215 9300 2233 9310
rect 2285 9300 2335 9310
rect 2399 9309 2408 9343
rect 2387 9300 2408 9309
rect 2215 9287 2408 9300
rect 2215 9271 2233 9287
rect 2285 9271 2335 9287
rect 2215 9237 2221 9271
rect 2285 9237 2293 9271
rect 2327 9237 2335 9271
rect 2387 9276 2408 9287
tri 2408 9276 2483 9351 sw
tri 13379 9276 13447 9344 se
rect 13447 9276 13453 16686
rect 2387 9270 13453 9276
rect 2215 9235 2233 9237
rect 2285 9235 2335 9237
rect 2215 9222 2365 9235
rect 2215 9198 2233 9222
rect 2285 9198 2335 9222
rect 2215 9164 2221 9198
rect 2285 9170 2293 9198
rect 2255 9164 2293 9170
rect 13631 9164 13637 16686
rect 2215 9157 2293 9164
rect 1821 9065 1827 9099
rect 1861 9065 1899 9099
rect 1933 9098 2083 9099
rect 1933 9065 1971 9098
rect 1821 9064 1971 9065
rect 2005 9097 2083 9098
rect 2005 9064 2043 9097
rect 1821 9063 2043 9064
rect 2077 9092 2083 9097
tri 2083 9092 2122 9131 sw
rect 2215 9105 2233 9157
rect 2285 9105 2293 9157
rect 2215 9092 2293 9105
rect 13559 9092 13637 9164
rect 13769 39504 14031 39541
rect 13769 39470 13775 39504
rect 13809 39503 14031 39504
rect 13809 39470 13847 39503
rect 13769 39469 13847 39470
rect 13881 39502 14031 39503
rect 13881 39469 13919 39502
rect 13769 39468 13919 39469
rect 13953 39468 13991 39502
rect 14025 39468 14031 39502
rect 13769 39431 14031 39468
rect 13769 39397 13775 39431
rect 13809 39430 14031 39431
rect 13809 39397 13847 39430
rect 13769 39396 13847 39397
rect 13881 39429 14031 39430
rect 13881 39396 13919 39429
rect 13769 39395 13919 39396
rect 13953 39395 13991 39429
rect 14025 39395 14031 39429
rect 13769 39358 14031 39395
rect 13769 39324 13775 39358
rect 13809 39357 14031 39358
rect 13809 39324 13847 39357
rect 13769 39323 13847 39324
rect 13881 39356 14031 39357
rect 13881 39323 13919 39356
rect 13769 39322 13919 39323
rect 13953 39322 13991 39356
rect 14025 39322 14031 39356
rect 13769 39285 14031 39322
rect 13769 39251 13775 39285
rect 13809 39284 14031 39285
rect 13809 39251 13847 39284
rect 13769 39250 13847 39251
rect 13881 39283 14031 39284
rect 13881 39250 13919 39283
rect 13769 39249 13919 39250
rect 13953 39249 13991 39283
rect 14025 39249 14031 39283
rect 13769 39212 14031 39249
rect 13769 39178 13775 39212
rect 13809 39211 14031 39212
rect 13809 39178 13847 39211
rect 13769 39177 13847 39178
rect 13881 39210 14031 39211
rect 13881 39177 13919 39210
rect 13769 39176 13919 39177
rect 13953 39176 13991 39210
rect 14025 39176 14031 39210
rect 13769 39139 14031 39176
rect 13769 39105 13775 39139
rect 13809 39138 14031 39139
rect 13809 39105 13847 39138
rect 13769 39104 13847 39105
rect 13881 39137 14031 39138
rect 13881 39104 13919 39137
rect 13769 39103 13919 39104
rect 13953 39103 13991 39137
rect 14025 39103 14031 39137
rect 13769 39066 14031 39103
rect 13769 39032 13775 39066
rect 13809 39065 14031 39066
rect 13809 39032 13847 39065
rect 13769 39031 13847 39032
rect 13881 39064 14031 39065
rect 13881 39031 13919 39064
rect 13769 39030 13919 39031
rect 13953 39030 13991 39064
rect 14025 39030 14031 39064
rect 13769 38993 14031 39030
rect 13769 38959 13775 38993
rect 13809 38992 14031 38993
rect 13809 38959 13847 38992
rect 13769 38958 13847 38959
rect 13881 38991 14031 38992
rect 13881 38958 13919 38991
rect 13769 38957 13919 38958
rect 13953 38957 13991 38991
rect 14025 38957 14031 38991
rect 13769 38920 14031 38957
rect 13769 38886 13775 38920
rect 13809 38919 14031 38920
rect 13809 38886 13847 38919
rect 13769 38885 13847 38886
rect 13881 38918 14031 38919
rect 13881 38885 13919 38918
rect 13769 38884 13919 38885
rect 13953 38884 13991 38918
rect 14025 38884 14031 38918
rect 13769 38847 14031 38884
rect 13769 38813 13775 38847
rect 13809 38846 14031 38847
rect 13809 38813 13847 38846
rect 13769 38812 13847 38813
rect 13881 38845 14031 38846
rect 13881 38812 13919 38845
rect 13769 38811 13919 38812
rect 13953 38811 13991 38845
rect 14025 38811 14031 38845
rect 13769 38774 14031 38811
rect 13769 38740 13775 38774
rect 13809 38773 14031 38774
rect 13809 38740 13847 38773
rect 13769 38739 13847 38740
rect 13881 38772 14031 38773
rect 13881 38739 13919 38772
rect 13769 38738 13919 38739
rect 13953 38738 13991 38772
rect 14025 38738 14031 38772
rect 13769 38701 14031 38738
rect 13769 38667 13775 38701
rect 13809 38700 14031 38701
rect 13809 38667 13847 38700
rect 13769 38666 13847 38667
rect 13881 38699 14031 38700
rect 13881 38666 13919 38699
rect 13769 38665 13919 38666
rect 13953 38665 13991 38699
rect 14025 38665 14031 38699
rect 13769 38628 14031 38665
rect 13769 38594 13775 38628
rect 13809 38627 14031 38628
rect 13809 38594 13847 38627
rect 13769 38593 13847 38594
rect 13881 38626 14031 38627
rect 13881 38593 13919 38626
rect 13769 38592 13919 38593
rect 13953 38592 13991 38626
rect 14025 38592 14031 38626
rect 13769 38555 14031 38592
rect 13769 38521 13775 38555
rect 13809 38554 14031 38555
rect 13809 38521 13847 38554
rect 13769 38520 13847 38521
rect 13881 38553 14031 38554
rect 13881 38520 13919 38553
rect 13769 38519 13919 38520
rect 13953 38519 13991 38553
rect 14025 38519 14031 38553
rect 13769 38482 14031 38519
rect 13769 38448 13775 38482
rect 13809 38481 14031 38482
rect 13809 38448 13847 38481
rect 13769 38447 13847 38448
rect 13881 38480 14031 38481
rect 13881 38447 13919 38480
rect 13769 38446 13919 38447
rect 13953 38446 13991 38480
rect 14025 38446 14031 38480
rect 13769 38409 14031 38446
rect 13769 38375 13775 38409
rect 13809 38408 14031 38409
rect 13809 38375 13847 38408
rect 13769 38374 13847 38375
rect 13881 38407 14031 38408
rect 13881 38374 13919 38407
rect 13769 38373 13919 38374
rect 13953 38373 13991 38407
rect 14025 38373 14031 38407
rect 13769 38336 14031 38373
rect 13769 38302 13775 38336
rect 13809 38335 14031 38336
rect 13809 38302 13847 38335
rect 13769 38301 13847 38302
rect 13881 38334 14031 38335
rect 13881 38301 13919 38334
rect 13769 38300 13919 38301
rect 13953 38300 13991 38334
rect 14025 38300 14031 38334
rect 13769 38263 14031 38300
rect 13769 38229 13775 38263
rect 13809 38262 14031 38263
rect 13809 38229 13847 38262
rect 13769 38228 13847 38229
rect 13881 38261 14031 38262
rect 13881 38228 13919 38261
rect 13769 38227 13919 38228
rect 13953 38227 13991 38261
rect 14025 38227 14031 38261
rect 13769 38190 14031 38227
rect 13769 38156 13775 38190
rect 13809 38189 14031 38190
rect 13809 38156 13847 38189
rect 13769 38155 13847 38156
rect 13881 38188 14031 38189
rect 13881 38155 13919 38188
rect 13769 38154 13919 38155
rect 13953 38154 13991 38188
rect 14025 38154 14031 38188
rect 13769 38117 14031 38154
rect 13769 38083 13775 38117
rect 13809 38116 14031 38117
rect 13809 38083 13847 38116
rect 13769 38082 13847 38083
rect 13881 38115 14031 38116
rect 13881 38082 13919 38115
rect 13769 38081 13919 38082
rect 13953 38081 13991 38115
rect 14025 38081 14031 38115
rect 13769 38044 14031 38081
rect 13769 38010 13775 38044
rect 13809 38043 14031 38044
rect 13809 38010 13847 38043
rect 13769 38009 13847 38010
rect 13881 38042 14031 38043
rect 13881 38009 13919 38042
rect 13769 38008 13919 38009
rect 13953 38008 13991 38042
rect 14025 38008 14031 38042
rect 13769 37971 14031 38008
rect 13769 37937 13775 37971
rect 13809 37970 14031 37971
rect 13809 37937 13847 37970
rect 13769 37936 13847 37937
rect 13881 37969 14031 37970
rect 13881 37936 13919 37969
rect 13769 37935 13919 37936
rect 13953 37935 13991 37969
rect 14025 37935 14031 37969
rect 13769 37898 14031 37935
rect 13769 37864 13775 37898
rect 13809 37897 14031 37898
rect 13809 37864 13847 37897
rect 13769 37863 13847 37864
rect 13881 37896 14031 37897
rect 13881 37863 13919 37896
rect 13769 37862 13919 37863
rect 13953 37862 13991 37896
rect 14025 37862 14031 37896
rect 13769 37825 14031 37862
rect 13769 37791 13775 37825
rect 13809 37824 14031 37825
rect 13809 37791 13847 37824
rect 13769 37790 13847 37791
rect 13881 37823 14031 37824
rect 13881 37790 13919 37823
rect 13769 37789 13919 37790
rect 13953 37789 13991 37823
rect 14025 37789 14031 37823
rect 13769 37752 14031 37789
rect 13769 37718 13775 37752
rect 13809 37751 14031 37752
rect 13809 37718 13847 37751
rect 13769 37717 13847 37718
rect 13881 37750 14031 37751
rect 13881 37717 13919 37750
rect 13769 37716 13919 37717
rect 13953 37716 13991 37750
rect 14025 37716 14031 37750
rect 13769 37679 14031 37716
rect 13769 37645 13775 37679
rect 13809 37678 14031 37679
rect 13809 37645 13847 37678
rect 13769 37644 13847 37645
rect 13881 37677 14031 37678
rect 13881 37644 13919 37677
rect 13769 37643 13919 37644
rect 13953 37643 13991 37677
rect 14025 37643 14031 37677
rect 13769 37606 14031 37643
rect 13769 37572 13775 37606
rect 13809 37605 14031 37606
rect 13809 37572 13847 37605
rect 13769 37571 13847 37572
rect 13881 37604 14031 37605
rect 13881 37571 13919 37604
rect 13769 37570 13919 37571
rect 13953 37570 13991 37604
rect 14025 37570 14031 37604
rect 13769 37533 14031 37570
rect 13769 37499 13775 37533
rect 13809 37532 14031 37533
rect 13809 37499 13847 37532
rect 13769 37498 13847 37499
rect 13881 37531 14031 37532
rect 13881 37498 13919 37531
rect 13769 37497 13919 37498
rect 13953 37497 13991 37531
rect 14025 37497 14031 37531
rect 13769 37460 14031 37497
rect 13769 37426 13775 37460
rect 13809 37459 14031 37460
rect 13809 37426 13847 37459
rect 13769 37425 13847 37426
rect 13881 37458 14031 37459
rect 13881 37425 13919 37458
rect 13769 37424 13919 37425
rect 13953 37424 13991 37458
rect 14025 37424 14031 37458
rect 13769 37387 14031 37424
rect 13769 37353 13775 37387
rect 13809 37386 14031 37387
rect 13809 37353 13847 37386
rect 13769 37352 13847 37353
rect 13881 37385 14031 37386
rect 13881 37352 13919 37385
rect 13769 37351 13919 37352
rect 13953 37351 13991 37385
rect 14025 37351 14031 37385
rect 13769 37314 14031 37351
rect 13769 37280 13775 37314
rect 13809 37313 14031 37314
rect 13809 37280 13847 37313
rect 13769 37279 13847 37280
rect 13881 37312 14031 37313
rect 13881 37279 13919 37312
rect 13769 37278 13919 37279
rect 13953 37278 13991 37312
rect 14025 37278 14031 37312
rect 13769 37241 14031 37278
rect 13769 37207 13775 37241
rect 13809 37240 14031 37241
rect 13809 37207 13847 37240
rect 13769 37206 13847 37207
rect 13881 37239 14031 37240
rect 13881 37206 13919 37239
rect 13769 37205 13919 37206
rect 13953 37205 13991 37239
rect 14025 37205 14031 37239
rect 13769 37168 14031 37205
rect 13769 37134 13775 37168
rect 13809 37167 14031 37168
rect 13809 37134 13847 37167
rect 13769 37133 13847 37134
rect 13881 37166 14031 37167
rect 13881 37133 13919 37166
rect 13769 37132 13919 37133
rect 13953 37132 13991 37166
rect 14025 37132 14031 37166
rect 13769 37095 14031 37132
rect 13769 37061 13775 37095
rect 13809 37094 14031 37095
rect 13809 37061 13847 37094
rect 13769 37060 13847 37061
rect 13881 37093 14031 37094
rect 13881 37060 13919 37093
rect 13769 37059 13919 37060
rect 13953 37059 13991 37093
rect 14025 37059 14031 37093
rect 13769 37022 14031 37059
rect 13769 36988 13775 37022
rect 13809 37021 14031 37022
rect 13809 36988 13847 37021
rect 13769 36987 13847 36988
rect 13881 37020 14031 37021
rect 13881 36987 13919 37020
rect 13769 36986 13919 36987
rect 13953 36986 13991 37020
rect 14025 36986 14031 37020
rect 13769 36949 14031 36986
rect 13769 36915 13775 36949
rect 13809 36948 14031 36949
rect 13809 36915 13847 36948
rect 13769 36914 13847 36915
rect 13881 36947 14031 36948
rect 13881 36914 13919 36947
rect 13769 36913 13919 36914
rect 13953 36913 13991 36947
rect 14025 36913 14031 36947
rect 13769 36876 14031 36913
rect 13769 36842 13775 36876
rect 13809 36875 14031 36876
rect 13809 36842 13847 36875
rect 13769 36841 13847 36842
rect 13881 36874 14031 36875
rect 13881 36841 13919 36874
rect 13769 36840 13919 36841
rect 13953 36840 13991 36874
rect 14025 36840 14031 36874
rect 13769 36803 14031 36840
rect 13769 36769 13775 36803
rect 13809 36802 14031 36803
rect 13809 36769 13847 36802
rect 13769 36768 13847 36769
rect 13881 36801 14031 36802
rect 13881 36768 13919 36801
rect 13769 36767 13919 36768
rect 13953 36767 13991 36801
rect 14025 36767 14031 36801
rect 13769 36730 14031 36767
rect 13769 36696 13775 36730
rect 13809 36729 14031 36730
rect 13809 36696 13847 36729
rect 13769 36695 13847 36696
rect 13881 36728 14031 36729
rect 13881 36695 13919 36728
rect 13769 36694 13919 36695
rect 13953 36694 13991 36728
rect 14025 36694 14031 36728
rect 13769 36657 14031 36694
rect 13769 36623 13775 36657
rect 13809 36656 14031 36657
rect 13809 36623 13847 36656
rect 13769 36622 13847 36623
rect 13881 36655 14031 36656
rect 13881 36622 13919 36655
rect 13769 36621 13919 36622
rect 13953 36621 13991 36655
rect 14025 36621 14031 36655
rect 13769 36584 14031 36621
rect 13769 36550 13775 36584
rect 13809 36583 14031 36584
rect 13809 36550 13847 36583
rect 13769 36549 13847 36550
rect 13881 36582 14031 36583
rect 13881 36549 13919 36582
rect 13769 36548 13919 36549
rect 13953 36548 13991 36582
rect 14025 36548 14031 36582
rect 13769 36511 14031 36548
rect 13769 36477 13775 36511
rect 13809 36510 14031 36511
rect 13809 36477 13847 36510
rect 13769 36476 13847 36477
rect 13881 36509 14031 36510
rect 13881 36476 13919 36509
rect 13769 36475 13919 36476
rect 13953 36475 13991 36509
rect 14025 36475 14031 36509
rect 13769 36438 14031 36475
rect 13769 36404 13775 36438
rect 13809 36437 14031 36438
rect 13809 36404 13847 36437
rect 13769 36403 13847 36404
rect 13881 36436 14031 36437
rect 13881 36403 13919 36436
rect 13769 36402 13919 36403
rect 13953 36402 13991 36436
rect 14025 36402 14031 36436
rect 13769 36365 14031 36402
rect 13769 36331 13775 36365
rect 13809 36364 14031 36365
rect 13809 36331 13847 36364
rect 13769 36330 13847 36331
rect 13881 36363 14031 36364
rect 13881 36330 13919 36363
rect 13769 36329 13919 36330
rect 13953 36329 13991 36363
rect 14025 36329 14031 36363
rect 13769 36292 14031 36329
rect 13769 36258 13775 36292
rect 13809 36291 14031 36292
rect 13809 36258 13847 36291
rect 13769 36257 13847 36258
rect 13881 36290 14031 36291
rect 13881 36257 13919 36290
rect 13769 36256 13919 36257
rect 13953 36256 13991 36290
rect 14025 36256 14031 36290
rect 13769 36219 14031 36256
rect 13769 36185 13775 36219
rect 13809 36218 14031 36219
rect 13809 36185 13847 36218
rect 13769 36184 13847 36185
rect 13881 36217 14031 36218
rect 13881 36184 13919 36217
rect 13769 36183 13919 36184
rect 13953 36183 13991 36217
rect 14025 36183 14031 36217
rect 13769 36146 14031 36183
rect 13769 36112 13775 36146
rect 13809 36145 14031 36146
rect 13809 36112 13847 36145
rect 13769 36111 13847 36112
rect 13881 36144 14031 36145
rect 13881 36111 13919 36144
rect 13769 36110 13919 36111
rect 13953 36110 13991 36144
rect 14025 36110 14031 36144
rect 13769 36073 14031 36110
rect 13769 36039 13775 36073
rect 13809 36072 14031 36073
rect 13809 36039 13847 36072
rect 13769 36038 13847 36039
rect 13881 36071 14031 36072
rect 13881 36038 13919 36071
rect 13769 36037 13919 36038
rect 13953 36037 13991 36071
rect 14025 36037 14031 36071
rect 13769 36000 14031 36037
rect 13769 35966 13775 36000
rect 13809 35999 14031 36000
rect 13809 35966 13847 35999
rect 13769 35965 13847 35966
rect 13881 35998 14031 35999
rect 13881 35965 13919 35998
rect 13769 35964 13919 35965
rect 13953 35964 13991 35998
rect 14025 35964 14031 35998
rect 13769 35927 14031 35964
rect 13769 35893 13775 35927
rect 13809 35926 14031 35927
rect 13809 35893 13847 35926
rect 13769 35892 13847 35893
rect 13881 35925 14031 35926
rect 13881 35892 13919 35925
rect 13769 35891 13919 35892
rect 13953 35891 13991 35925
rect 14025 35891 14031 35925
rect 13769 35854 14031 35891
rect 13769 35820 13775 35854
rect 13809 35853 14031 35854
rect 13809 35820 13847 35853
rect 13769 35819 13847 35820
rect 13881 35852 14031 35853
rect 13881 35819 13919 35852
rect 13769 35818 13919 35819
rect 13953 35818 13991 35852
rect 14025 35818 14031 35852
rect 13769 35781 14031 35818
rect 13769 35747 13775 35781
rect 13809 35780 14031 35781
rect 13809 35747 13847 35780
rect 13769 35746 13847 35747
rect 13881 35779 14031 35780
rect 13881 35746 13919 35779
rect 13769 35745 13919 35746
rect 13953 35745 13991 35779
rect 14025 35745 14031 35779
rect 13769 35708 14031 35745
rect 13769 35674 13775 35708
rect 13809 35707 14031 35708
rect 13809 35674 13847 35707
rect 13769 35673 13847 35674
rect 13881 35706 14031 35707
rect 13881 35673 13919 35706
rect 13769 35672 13919 35673
rect 13953 35672 13991 35706
rect 14025 35672 14031 35706
rect 13769 35635 14031 35672
rect 13769 35601 13775 35635
rect 13809 35634 14031 35635
rect 13809 35601 13847 35634
rect 13769 35600 13847 35601
rect 13881 35633 14031 35634
rect 13881 35600 13919 35633
rect 13769 35599 13919 35600
rect 13953 35599 13991 35633
rect 14025 35599 14031 35633
rect 13769 35562 14031 35599
rect 13769 35528 13775 35562
rect 13809 35561 14031 35562
rect 13809 35528 13847 35561
rect 13769 35527 13847 35528
rect 13881 35560 14031 35561
rect 13881 35527 13919 35560
rect 13769 35526 13919 35527
rect 13953 35526 13991 35560
rect 14025 35526 14031 35560
rect 13769 35489 14031 35526
rect 13769 35455 13775 35489
rect 13809 35488 14031 35489
rect 13809 35455 13847 35488
rect 13769 35454 13847 35455
rect 13881 35487 14031 35488
rect 13881 35454 13919 35487
rect 13769 35453 13919 35454
rect 13953 35453 13991 35487
rect 14025 35453 14031 35487
rect 13769 35416 14031 35453
rect 13769 35382 13775 35416
rect 13809 35415 14031 35416
rect 13809 35382 13847 35415
rect 13769 35381 13847 35382
rect 13881 35414 14031 35415
rect 13881 35381 13919 35414
rect 13769 35380 13919 35381
rect 13953 35380 13991 35414
rect 14025 35380 14031 35414
rect 13769 35343 14031 35380
rect 13769 35309 13775 35343
rect 13809 35342 14031 35343
rect 13809 35309 13847 35342
rect 13769 35308 13847 35309
rect 13881 35341 14031 35342
rect 13881 35308 13919 35341
rect 13769 35307 13919 35308
rect 13953 35307 13991 35341
rect 14025 35307 14031 35341
rect 13769 35270 14031 35307
rect 13769 35236 13775 35270
rect 13809 35269 14031 35270
rect 13809 35236 13847 35269
rect 13769 35235 13847 35236
rect 13881 35268 14031 35269
rect 13881 35235 13919 35268
rect 13769 35234 13919 35235
rect 13953 35234 13991 35268
rect 14025 35234 14031 35268
rect 13769 35197 14031 35234
rect 13769 35163 13775 35197
rect 13809 35196 14031 35197
rect 13809 35163 13847 35196
rect 13769 35162 13847 35163
rect 13881 35195 14031 35196
rect 13881 35162 13919 35195
rect 13769 35161 13919 35162
rect 13953 35161 13991 35195
rect 14025 35161 14031 35195
rect 13769 35124 14031 35161
rect 13769 35090 13775 35124
rect 13809 35123 14031 35124
rect 13809 35090 13847 35123
rect 13769 35089 13847 35090
rect 13881 35122 14031 35123
rect 13881 35089 13919 35122
rect 13769 35051 13919 35089
rect 13769 35017 13775 35051
rect 13809 35050 13919 35051
rect 13809 35017 13847 35050
rect 13769 34978 13847 35017
rect 13769 32712 13775 34978
rect 14025 32712 14031 35122
rect 13769 32657 14031 32712
rect 13769 32623 13775 32657
rect 13809 32623 13847 32657
rect 13881 32623 13919 32657
rect 13953 32623 13991 32657
rect 14025 32623 14031 32657
rect 13769 32584 14031 32623
rect 13769 32550 13775 32584
rect 13809 32550 13847 32584
rect 13881 32550 13919 32584
rect 13953 32550 13991 32584
rect 14025 32550 14031 32584
rect 13769 32511 14031 32550
rect 13769 32477 13775 32511
rect 13809 32477 13847 32511
rect 13881 32477 13919 32511
rect 13953 32477 13991 32511
rect 14025 32477 14031 32511
rect 13769 32438 14031 32477
rect 13769 32404 13775 32438
rect 13809 32404 13847 32438
rect 13881 32404 13919 32438
rect 13953 32404 13991 32438
rect 14025 32404 14031 32438
rect 13769 32365 14031 32404
rect 13769 32331 13775 32365
rect 13809 32331 13847 32365
rect 13881 32331 13919 32365
rect 13953 32331 13991 32365
rect 14025 32331 14031 32365
rect 13769 32292 14031 32331
rect 13769 32258 13775 32292
rect 13809 32258 13847 32292
rect 13881 32258 13919 32292
rect 13953 32258 13991 32292
rect 14025 32258 14031 32292
rect 13769 32219 14031 32258
rect 13769 32185 13775 32219
rect 13809 32185 13847 32219
rect 13881 32185 13919 32219
rect 13953 32185 13991 32219
rect 14025 32185 14031 32219
rect 13769 32146 14031 32185
rect 13769 32112 13775 32146
rect 13809 32112 13847 32146
rect 13881 32112 13919 32146
rect 13953 32112 13991 32146
rect 14025 32112 14031 32146
rect 13769 32073 14031 32112
rect 13769 32039 13775 32073
rect 13809 32039 13847 32073
rect 13881 32039 13919 32073
rect 13953 32039 13991 32073
rect 14025 32039 14031 32073
rect 13769 32000 14031 32039
rect 13769 31966 13775 32000
rect 13809 31966 13847 32000
rect 13881 31966 13919 32000
rect 13953 31966 13991 32000
rect 14025 31966 14031 32000
rect 13769 31927 14031 31966
rect 13769 31893 13775 31927
rect 13809 31893 13847 31927
rect 13881 31893 13919 31927
rect 13953 31893 13991 31927
rect 14025 31893 14031 31927
rect 13769 31854 14031 31893
rect 13769 31820 13775 31854
rect 13809 31820 13847 31854
rect 13881 31820 13919 31854
rect 13953 31820 13991 31854
rect 14025 31820 14031 31854
rect 13769 31781 14031 31820
rect 13769 31747 13775 31781
rect 13809 31747 13847 31781
rect 13881 31747 13919 31781
rect 13953 31747 13991 31781
rect 14025 31747 14031 31781
rect 13769 31708 14031 31747
rect 13769 31674 13775 31708
rect 13809 31674 13847 31708
rect 13881 31674 13919 31708
rect 13953 31674 13991 31708
rect 14025 31674 14031 31708
rect 13769 31635 14031 31674
rect 13769 31601 13775 31635
rect 13809 31601 13847 31635
rect 13881 31601 13919 31635
rect 13953 31601 13991 31635
rect 14025 31601 14031 31635
rect 13769 31562 14031 31601
rect 13769 31528 13775 31562
rect 13809 31528 13847 31562
rect 13881 31528 13919 31562
rect 13953 31528 13991 31562
rect 14025 31528 14031 31562
rect 13769 31489 14031 31528
rect 13769 31455 13775 31489
rect 13809 31455 13847 31489
rect 13881 31455 13919 31489
rect 13953 31455 13991 31489
rect 14025 31455 14031 31489
rect 13769 31416 14031 31455
rect 13769 31382 13775 31416
rect 13809 31382 13847 31416
rect 13881 31382 13919 31416
rect 13953 31382 13991 31416
rect 14025 31382 14031 31416
rect 13769 31343 14031 31382
rect 13769 31309 13775 31343
rect 13809 31309 13847 31343
rect 13881 31309 13919 31343
rect 13953 31309 13991 31343
rect 14025 31309 14031 31343
rect 13769 31270 14031 31309
rect 13769 31236 13775 31270
rect 13809 31236 13847 31270
rect 13881 31236 13919 31270
rect 13953 31236 13991 31270
rect 14025 31236 14031 31270
rect 13769 31197 14031 31236
rect 13769 31163 13775 31197
rect 13809 31163 13847 31197
rect 13881 31163 13919 31197
rect 13953 31163 13991 31197
rect 14025 31163 14031 31197
rect 13769 31124 14031 31163
rect 13769 31090 13775 31124
rect 13809 31090 13847 31124
rect 13881 31090 13919 31124
rect 13953 31090 13991 31124
rect 14025 31090 14031 31124
rect 13769 31051 14031 31090
rect 13769 31017 13775 31051
rect 13809 31017 13847 31051
rect 13881 31017 13919 31051
rect 13953 31017 13991 31051
rect 14025 31017 14031 31051
rect 13769 30978 14031 31017
rect 13769 30944 13775 30978
rect 13809 30944 13847 30978
rect 13881 30944 13919 30978
rect 13953 30944 13991 30978
rect 14025 30944 14031 30978
rect 13769 30905 14031 30944
rect 13769 30871 13775 30905
rect 13809 30871 13847 30905
rect 13881 30871 13919 30905
rect 13953 30871 13991 30905
rect 14025 30871 14031 30905
rect 13769 30832 14031 30871
rect 13769 30798 13775 30832
rect 13809 30798 13847 30832
rect 13881 30798 13919 30832
rect 13953 30798 13991 30832
rect 14025 30798 14031 30832
rect 13769 30759 14031 30798
rect 13769 30725 13775 30759
rect 13809 30725 13847 30759
rect 13881 30725 13919 30759
rect 13953 30725 13991 30759
rect 14025 30725 14031 30759
rect 13769 30686 14031 30725
rect 13769 30652 13775 30686
rect 13809 30652 13847 30686
rect 13881 30652 13919 30686
rect 13953 30652 13991 30686
rect 14025 30652 14031 30686
rect 13769 30613 14031 30652
rect 13769 30579 13775 30613
rect 13809 30579 13847 30613
rect 13881 30579 13919 30613
rect 13953 30579 13991 30613
rect 14025 30579 14031 30613
rect 13769 30540 14031 30579
rect 13769 30506 13775 30540
rect 13809 30506 13847 30540
rect 13881 30506 13919 30540
rect 13953 30506 13991 30540
rect 14025 30506 14031 30540
rect 13769 30467 14031 30506
rect 13769 30433 13775 30467
rect 13809 30433 13847 30467
rect 13881 30433 13919 30467
rect 13953 30433 13991 30467
rect 14025 30433 14031 30467
rect 13769 30394 14031 30433
rect 13769 30360 13775 30394
rect 13809 30360 13847 30394
rect 13881 30360 13919 30394
rect 13953 30360 13991 30394
rect 14025 30360 14031 30394
rect 13769 30321 14031 30360
rect 13769 30287 13775 30321
rect 13809 30287 13847 30321
rect 13881 30287 13919 30321
rect 13953 30287 13991 30321
rect 14025 30287 14031 30321
rect 13769 30248 14031 30287
rect 13769 30214 13775 30248
rect 13809 30214 13847 30248
rect 13881 30214 13919 30248
rect 13953 30214 13991 30248
rect 14025 30214 14031 30248
rect 13769 30175 14031 30214
rect 13769 30141 13775 30175
rect 13809 30141 13847 30175
rect 13881 30141 13919 30175
rect 13953 30141 13991 30175
rect 14025 30141 14031 30175
rect 13769 30102 14031 30141
rect 13769 30068 13775 30102
rect 13809 30068 13847 30102
rect 13881 30068 13919 30102
rect 13953 30068 13991 30102
rect 14025 30068 14031 30102
rect 13769 30029 14031 30068
rect 13769 29995 13775 30029
rect 13809 29995 13847 30029
rect 13881 29995 13919 30029
rect 13953 29995 13991 30029
rect 14025 29995 14031 30029
rect 13769 29956 14031 29995
rect 13769 29922 13775 29956
rect 13809 29922 13847 29956
rect 13881 29922 13919 29956
rect 13953 29922 13991 29956
rect 14025 29922 14031 29956
rect 13769 29883 14031 29922
rect 13769 29849 13775 29883
rect 13809 29849 13847 29883
rect 13881 29849 13919 29883
rect 13953 29849 13991 29883
rect 14025 29849 14031 29883
rect 13769 29810 14031 29849
rect 13769 29776 13775 29810
rect 13809 29776 13847 29810
rect 13881 29776 13919 29810
rect 13953 29776 13991 29810
rect 14025 29776 14031 29810
rect 13769 29737 14031 29776
rect 13769 29703 13775 29737
rect 13809 29703 13847 29737
rect 13881 29703 13919 29737
rect 13953 29703 13991 29737
rect 14025 29703 14031 29737
rect 13769 29664 14031 29703
rect 13769 29630 13775 29664
rect 13809 29630 13847 29664
rect 13881 29630 13919 29664
rect 13953 29630 13991 29664
rect 14025 29630 14031 29664
rect 13769 29591 14031 29630
rect 13769 29557 13775 29591
rect 13809 29557 13847 29591
rect 13881 29557 13919 29591
rect 13953 29557 13991 29591
rect 14025 29557 14031 29591
rect 13769 29518 14031 29557
rect 13769 29484 13775 29518
rect 13809 29484 13847 29518
rect 13881 29484 13919 29518
rect 13953 29484 13991 29518
rect 14025 29484 14031 29518
rect 13769 29445 14031 29484
rect 13769 29411 13775 29445
rect 13809 29411 13847 29445
rect 13881 29411 13919 29445
rect 13953 29411 13991 29445
rect 14025 29411 14031 29445
rect 13769 29372 14031 29411
rect 13769 29338 13775 29372
rect 13809 29338 13847 29372
rect 13881 29338 13919 29372
rect 13953 29338 13991 29372
rect 14025 29338 14031 29372
rect 13769 29299 14031 29338
rect 13769 29265 13775 29299
rect 13809 29265 13847 29299
rect 13881 29265 13919 29299
rect 13953 29265 13991 29299
rect 14025 29265 14031 29299
rect 13769 29226 14031 29265
rect 13769 29192 13775 29226
rect 13809 29192 13847 29226
rect 13881 29192 13919 29226
rect 13953 29192 13991 29226
rect 14025 29192 14031 29226
rect 13769 29153 14031 29192
rect 13769 29119 13775 29153
rect 13809 29119 13847 29153
rect 13881 29119 13919 29153
rect 13953 29119 13991 29153
rect 14025 29119 14031 29153
rect 13769 29080 14031 29119
rect 13769 29046 13775 29080
rect 13809 29046 13847 29080
rect 13881 29046 13919 29080
rect 13953 29046 13991 29080
rect 14025 29046 14031 29080
rect 13769 29007 14031 29046
rect 13769 28973 13775 29007
rect 13809 28973 13847 29007
rect 13881 28973 13919 29007
rect 13953 28973 13991 29007
rect 14025 28973 14031 29007
rect 13769 28934 14031 28973
rect 13769 28900 13775 28934
rect 13809 28900 13847 28934
rect 13881 28900 13919 28934
rect 13953 28900 13991 28934
rect 14025 28900 14031 28934
rect 13769 28861 14031 28900
rect 13769 28827 13775 28861
rect 13809 28827 13847 28861
rect 13881 28827 13919 28861
rect 13953 28827 13991 28861
rect 14025 28827 14031 28861
rect 13769 28788 14031 28827
rect 13769 28754 13775 28788
rect 13809 28754 13847 28788
rect 13881 28754 13919 28788
rect 13953 28754 13991 28788
rect 14025 28754 14031 28788
rect 13769 28715 14031 28754
rect 13769 28681 13775 28715
rect 13809 28681 13847 28715
rect 13881 28681 13919 28715
rect 13953 28681 13991 28715
rect 14025 28681 14031 28715
rect 13769 28642 14031 28681
rect 13769 28608 13775 28642
rect 13809 28608 13847 28642
rect 13881 28608 13919 28642
rect 13953 28608 13991 28642
rect 14025 28608 14031 28642
rect 13769 28569 14031 28608
rect 13769 28535 13775 28569
rect 13809 28535 13847 28569
rect 13881 28535 13919 28569
rect 13953 28535 13991 28569
rect 14025 28535 14031 28569
rect 13769 28496 14031 28535
rect 13769 28462 13775 28496
rect 13809 28462 13847 28496
rect 13881 28462 13919 28496
rect 13953 28462 13991 28496
rect 14025 28462 14031 28496
rect 13769 28423 14031 28462
rect 13769 9165 13775 28423
rect 14025 9165 14031 28423
rect 13769 9121 14031 9165
rect 13769 9119 13919 9121
rect 13769 9116 13847 9119
rect 2077 9086 2122 9092
tri 2122 9086 2128 9092 sw
rect 2215 9086 13637 9092
tri 13750 9086 13769 9105 se
rect 13769 9086 13775 9116
rect 2077 9082 2128 9086
tri 2128 9082 2132 9086 sw
tri 13746 9082 13750 9086 se
rect 13750 9082 13775 9086
rect 13809 9085 13847 9116
rect 13881 9087 13919 9119
rect 13953 9087 13991 9121
rect 14025 9087 14031 9121
rect 13881 9085 14031 9087
rect 13809 9082 14031 9085
rect 2077 9063 2132 9082
rect 1821 9043 2132 9063
tri 2132 9043 2171 9082 sw
tri 13707 9043 13746 9082 se
rect 13746 9043 14031 9082
rect 1821 9039 2171 9043
tri 2171 9039 2175 9043 sw
tri 13703 9039 13707 9043 se
rect 13707 9039 13919 9043
rect 1821 9033 2175 9039
tri 2175 9033 2181 9039 sw
tri 13697 9033 13703 9039 se
rect 13703 9033 13847 9039
rect 1821 9026 2181 9033
rect 1821 8992 1827 9026
rect 1861 8992 1899 9026
rect 1933 9025 2181 9026
rect 1933 8992 1971 9025
rect 1821 8991 1971 8992
rect 2005 9024 2181 9025
rect 2005 8991 2043 9024
rect 1821 8990 2043 8991
rect 2077 8999 2181 9024
tri 2181 8999 2215 9033 sw
tri 13663 8999 13697 9033 se
rect 13697 8999 13775 9033
rect 13809 9005 13847 9033
rect 13881 9009 13919 9039
rect 13953 9009 13991 9043
rect 14025 9009 14031 9043
rect 13881 9005 14031 9009
rect 13809 8999 14031 9005
rect 2077 8990 2215 8999
rect 1821 8966 2215 8990
tri 2215 8966 2248 8999 sw
tri 13630 8966 13663 8999 se
rect 13663 8966 14031 8999
rect 1821 8959 2248 8966
tri 2248 8959 2255 8966 sw
tri 13623 8959 13630 8966 se
rect 13630 8959 13919 8966
rect 1821 8957 2255 8959
tri 2255 8957 2257 8959 sw
tri 13621 8957 13623 8959 se
rect 13623 8957 13847 8959
rect 1821 8953 13847 8957
rect 1821 8919 1827 8953
rect 1861 8919 1899 8953
rect 1933 8952 13847 8953
rect 1933 8919 1971 8952
rect 1821 8918 1971 8919
rect 2005 8951 13847 8952
rect 2005 8918 2043 8951
rect 1821 8880 2043 8918
rect 1821 8846 1827 8880
rect 1861 8846 1899 8880
rect 1933 8879 2043 8880
rect 8845 8917 8884 8951
rect 8918 8917 8957 8951
rect 8991 8917 9030 8951
rect 9064 8917 9103 8951
rect 9137 8917 9176 8951
rect 9210 8917 9249 8951
rect 9283 8917 9322 8951
rect 9356 8917 9395 8951
rect 9429 8917 9468 8951
rect 9502 8917 9541 8951
rect 9575 8917 9614 8951
rect 9648 8917 9687 8951
rect 9721 8917 9760 8951
rect 9794 8917 9833 8951
rect 9867 8917 9906 8951
rect 9940 8917 9979 8951
rect 10013 8917 10052 8951
rect 10086 8917 10125 8951
rect 10159 8917 10198 8951
rect 10232 8917 10271 8951
rect 10305 8917 10344 8951
rect 10378 8917 10417 8951
rect 10451 8917 10490 8951
rect 10524 8917 10563 8951
rect 10597 8917 10636 8951
rect 10670 8917 10709 8951
rect 10743 8917 10782 8951
rect 10816 8917 10855 8951
rect 10889 8917 10928 8951
rect 10962 8917 11001 8951
rect 11035 8917 11074 8951
rect 11108 8917 11147 8951
rect 11181 8917 11220 8951
rect 11254 8917 11293 8951
rect 11327 8917 11366 8951
rect 11400 8917 11439 8951
rect 11473 8917 11512 8951
rect 11546 8917 11585 8951
rect 11619 8917 11658 8951
rect 11692 8917 11731 8951
rect 11765 8917 11804 8951
rect 11838 8917 11877 8951
rect 11911 8917 11950 8951
rect 11984 8917 12023 8951
rect 12057 8917 12096 8951
rect 12130 8917 12169 8951
rect 12203 8917 12242 8951
rect 12276 8917 12315 8951
rect 12349 8917 12388 8951
rect 12422 8917 12461 8951
rect 12495 8917 12534 8951
rect 12568 8917 12607 8951
rect 12641 8917 12680 8951
rect 12714 8917 12753 8951
rect 12787 8917 12826 8951
rect 12860 8917 12899 8951
rect 12933 8917 12972 8951
rect 13006 8917 13045 8951
rect 13079 8917 13118 8951
rect 13152 8917 13191 8951
rect 13225 8917 13264 8951
rect 13298 8917 13337 8951
rect 13371 8917 13410 8951
rect 13444 8917 13483 8951
rect 13517 8917 13556 8951
rect 13590 8917 13629 8951
rect 13663 8917 13702 8951
rect 13736 8917 13775 8951
rect 13809 8925 13847 8951
rect 13881 8932 13919 8959
rect 13953 8932 13991 8966
rect 14025 8932 14031 8966
rect 13881 8925 14031 8932
rect 13809 8917 14031 8925
rect 8845 8889 14031 8917
rect 8845 8881 13919 8889
rect 8845 8879 11204 8881
rect 1933 8846 1971 8879
rect 1821 8807 1971 8846
rect 8917 8845 8956 8879
rect 8990 8845 9029 8879
rect 9063 8845 9102 8879
rect 9136 8845 9175 8879
rect 9209 8845 9248 8879
rect 9282 8845 9321 8879
rect 9355 8845 9394 8879
rect 9428 8845 9467 8879
rect 9501 8845 9540 8879
rect 9574 8845 9613 8879
rect 9647 8845 9686 8879
rect 9720 8845 9759 8879
rect 9793 8845 9832 8879
rect 9866 8845 9905 8879
rect 9939 8845 9978 8879
rect 10012 8845 10051 8879
rect 10085 8845 10124 8879
rect 10158 8845 10197 8879
rect 10231 8845 10270 8879
rect 10304 8845 10343 8879
rect 10377 8845 10416 8879
rect 10450 8845 10489 8879
rect 10523 8845 10562 8879
rect 10596 8845 10635 8879
rect 10669 8845 10708 8879
rect 10742 8845 10781 8879
rect 10815 8845 10854 8879
rect 10888 8845 10927 8879
rect 10961 8845 11000 8879
rect 11034 8845 11073 8879
rect 11107 8845 11146 8879
rect 11180 8845 11204 8879
rect 8917 8829 11204 8845
rect 11256 8829 11274 8881
rect 11326 8829 11344 8881
rect 11396 8879 11414 8881
rect 11466 8879 11483 8881
rect 11535 8879 11552 8881
rect 11604 8879 11621 8881
rect 11673 8879 11690 8881
rect 11742 8879 11759 8881
rect 11811 8879 11828 8881
rect 11880 8879 11897 8881
rect 11949 8879 13919 8881
rect 11399 8845 11414 8879
rect 11472 8845 11483 8879
rect 11545 8845 11552 8879
rect 11618 8845 11621 8879
rect 11983 8845 12022 8879
rect 12056 8845 12095 8879
rect 12129 8845 12168 8879
rect 12202 8845 12241 8879
rect 12275 8845 12314 8879
rect 12348 8845 12387 8879
rect 12421 8845 12460 8879
rect 12494 8845 12533 8879
rect 12567 8845 12606 8879
rect 12640 8845 12679 8879
rect 12713 8845 12752 8879
rect 12786 8845 12825 8879
rect 12859 8845 12898 8879
rect 12932 8845 12971 8879
rect 13005 8845 13044 8879
rect 13078 8845 13117 8879
rect 13151 8845 13190 8879
rect 13224 8845 13263 8879
rect 13297 8845 13336 8879
rect 13370 8845 13409 8879
rect 13443 8845 13482 8879
rect 13516 8845 13555 8879
rect 13589 8845 13628 8879
rect 13662 8845 13701 8879
rect 13735 8845 13774 8879
rect 13808 8845 13847 8879
rect 13881 8855 13919 8879
rect 13953 8855 13991 8889
rect 14025 8855 14031 8889
rect 13881 8845 14031 8855
rect 11396 8829 11414 8845
rect 11466 8829 11483 8845
rect 11535 8829 11552 8845
rect 11604 8829 11621 8845
rect 11673 8829 11690 8845
rect 11742 8829 11759 8845
rect 11811 8829 11828 8845
rect 11880 8829 11897 8845
rect 11949 8829 14031 8845
rect 8917 8812 14031 8829
rect 8917 8807 13991 8812
rect 357 8773 470 8779
tri 470 8773 476 8779 nw
rect 1821 8773 1827 8807
rect 1861 8773 1899 8807
rect 357 5403 437 8773
tri 437 8740 470 8773 nw
rect 1821 8701 1899 8773
rect 8989 8773 9028 8807
rect 9062 8773 9101 8807
rect 9135 8773 9174 8807
rect 9208 8773 9247 8807
rect 9281 8773 9320 8807
rect 9354 8773 9393 8807
rect 9427 8773 9466 8807
rect 9500 8773 9539 8807
rect 9573 8773 9612 8807
rect 9646 8773 9685 8807
rect 9719 8773 9758 8807
rect 9792 8773 9831 8807
rect 9865 8773 9904 8807
rect 9938 8773 9977 8807
rect 10011 8773 10050 8807
rect 10084 8773 10123 8807
rect 10157 8773 10196 8807
rect 10230 8773 10269 8807
rect 10303 8773 10342 8807
rect 10376 8773 10415 8807
rect 10449 8773 10488 8807
rect 10522 8773 10561 8807
rect 10595 8773 10634 8807
rect 10668 8773 10707 8807
rect 10741 8773 10780 8807
rect 10814 8773 10853 8807
rect 10887 8773 10926 8807
rect 10960 8773 10999 8807
rect 11033 8773 11072 8807
rect 11106 8773 11145 8807
rect 11179 8773 11218 8807
rect 11252 8773 11291 8807
rect 11325 8773 11364 8807
rect 11398 8773 11437 8807
rect 11471 8773 11510 8807
rect 11544 8773 11583 8807
rect 11617 8773 11656 8807
rect 11690 8773 11729 8807
rect 11763 8773 11802 8807
rect 11836 8773 11875 8807
rect 11909 8773 11948 8807
rect 11982 8773 12021 8807
rect 12055 8773 12094 8807
rect 12128 8773 12167 8807
rect 12201 8773 12240 8807
rect 12274 8773 12313 8807
rect 12347 8773 12386 8807
rect 12420 8773 12459 8807
rect 12493 8773 12532 8807
rect 12566 8773 12605 8807
rect 12639 8773 12678 8807
rect 12712 8773 12751 8807
rect 12785 8773 12824 8807
rect 12858 8773 12897 8807
rect 12931 8773 12970 8807
rect 13004 8773 13043 8807
rect 13077 8773 13116 8807
rect 13150 8773 13189 8807
rect 13223 8773 13262 8807
rect 13296 8773 13335 8807
rect 13369 8773 13408 8807
rect 13442 8773 13481 8807
rect 13515 8773 13554 8807
rect 13588 8773 13627 8807
rect 13661 8773 13700 8807
rect 13734 8773 13773 8807
rect 13807 8773 13846 8807
rect 13880 8773 13919 8807
rect 13953 8778 13991 8807
rect 14025 8778 14031 8812
rect 13953 8773 14031 8778
rect 8989 8759 14031 8773
rect 8989 8735 11204 8759
rect 8989 8701 9028 8735
rect 9062 8701 9101 8735
rect 9135 8701 9174 8735
rect 9208 8701 9247 8735
rect 9281 8701 9320 8735
rect 9354 8701 9393 8735
rect 9427 8701 9466 8735
rect 9500 8701 9539 8735
rect 9573 8701 9612 8735
rect 9646 8701 9685 8735
rect 9719 8701 9758 8735
rect 9792 8701 9831 8735
rect 9865 8701 9904 8735
rect 9938 8701 9977 8735
rect 10011 8701 10050 8735
rect 10084 8701 10123 8735
rect 10157 8701 10196 8735
rect 10230 8701 10269 8735
rect 10303 8701 10342 8735
rect 10376 8701 10415 8735
rect 10449 8701 10488 8735
rect 10522 8701 10561 8735
rect 10595 8701 10634 8735
rect 10668 8701 10707 8735
rect 10741 8701 10780 8735
rect 10814 8701 10853 8735
rect 10887 8701 10926 8735
rect 10960 8701 10999 8735
rect 11033 8701 11072 8735
rect 11106 8701 11145 8735
rect 11179 8707 11204 8735
rect 11256 8707 11274 8759
rect 11326 8707 11344 8759
rect 11396 8735 11414 8759
rect 11466 8735 11483 8759
rect 11535 8735 11552 8759
rect 11604 8735 11621 8759
rect 11673 8735 11690 8759
rect 11742 8735 11759 8759
rect 11811 8735 11828 8759
rect 11880 8735 11897 8759
rect 11949 8735 14031 8759
rect 11398 8707 11414 8735
rect 11471 8707 11483 8735
rect 11544 8707 11552 8735
rect 11617 8707 11621 8735
rect 11179 8701 11218 8707
rect 11252 8701 11291 8707
rect 11325 8701 11364 8707
rect 11398 8701 11437 8707
rect 11471 8701 11510 8707
rect 11544 8701 11583 8707
rect 11617 8701 11656 8707
rect 11690 8701 11729 8707
rect 11763 8701 11802 8707
rect 11836 8701 11875 8707
rect 11909 8701 11948 8707
rect 11982 8701 12021 8735
rect 12055 8701 12094 8735
rect 12128 8701 12167 8735
rect 12201 8701 12240 8735
rect 12274 8701 12313 8735
rect 12347 8701 12386 8735
rect 12420 8701 12459 8735
rect 12493 8701 12532 8735
rect 12566 8701 12605 8735
rect 12639 8701 12678 8735
rect 12712 8701 12751 8735
rect 12785 8701 12824 8735
rect 12858 8701 12897 8735
rect 12931 8701 12970 8735
rect 13004 8701 13043 8735
rect 13077 8701 13116 8735
rect 13150 8701 13189 8735
rect 13223 8701 13262 8735
rect 13296 8701 13335 8735
rect 13369 8701 13408 8735
rect 13442 8701 13481 8735
rect 13515 8701 13554 8735
rect 13588 8701 13627 8735
rect 13661 8701 13700 8735
rect 13734 8701 13773 8735
rect 13807 8701 13846 8735
rect 13880 8701 13919 8735
rect 13953 8701 14031 8735
rect 1821 8695 14031 8701
rect 1598 8688 1728 8694
rect 1598 8654 1610 8688
rect 1644 8654 1682 8688
rect 1716 8654 1728 8688
rect 1598 8648 1728 8654
tri 1632 8600 1680 8648 ne
rect 1680 8605 1728 8648
tri 1728 8605 1762 8639 sw
rect 1680 8598 14212 8605
rect 1680 8564 14094 8598
rect 14128 8564 14166 8598
rect 14200 8564 14212 8598
rect 1680 8557 14212 8564
rect 14476 8596 14524 39836
tri 14524 39802 14558 39836 nw
tri 14524 8596 14576 8648 sw
rect 14476 8548 14724 8596
tri 14598 8505 14641 8548 ne
rect 14641 8505 14724 8548
rect 10458 8499 13779 8505
rect 10458 8465 10536 8499
rect 10570 8465 10609 8499
rect 10643 8465 10682 8499
rect 10716 8465 10755 8499
rect 10789 8465 10828 8499
rect 10862 8465 10901 8499
rect 10935 8465 10974 8499
rect 11008 8465 11047 8499
rect 11081 8465 11120 8499
rect 11154 8465 11193 8499
rect 11227 8495 11266 8499
rect 11300 8495 11339 8499
rect 11373 8495 11412 8499
rect 11446 8495 11485 8499
rect 11519 8495 11558 8499
rect 11592 8495 11631 8499
rect 11665 8495 11704 8499
rect 11738 8495 11777 8499
rect 11811 8495 11850 8499
rect 11884 8495 11923 8499
rect 11256 8465 11266 8495
rect 11326 8465 11339 8495
rect 11396 8465 11412 8495
rect 10458 8443 11204 8465
rect 11256 8443 11274 8465
rect 11326 8443 11344 8465
rect 11396 8443 11414 8465
rect 11466 8443 11483 8495
rect 11535 8443 11552 8495
rect 11604 8443 11621 8495
rect 11673 8443 11690 8495
rect 11742 8443 11759 8495
rect 11811 8443 11828 8495
rect 11884 8465 11897 8495
rect 11957 8465 11996 8499
rect 12030 8465 12069 8499
rect 12103 8465 12142 8499
rect 12176 8465 12215 8499
rect 12249 8465 12288 8499
rect 12322 8465 12361 8499
rect 12395 8465 12434 8499
rect 12468 8465 12507 8499
rect 12541 8465 12580 8499
rect 12614 8465 12653 8499
rect 12687 8465 12726 8499
rect 12760 8465 12799 8499
rect 12833 8465 12872 8499
rect 12906 8465 12945 8499
rect 12979 8465 13018 8499
rect 13052 8465 13091 8499
rect 11880 8443 11897 8465
rect 11949 8443 13091 8465
rect 10458 8427 13091 8443
rect 10458 8426 10536 8427
rect 10458 8392 10464 8426
rect 10498 8393 10536 8426
rect 10570 8393 10609 8427
rect 10643 8393 10682 8427
rect 10716 8393 10755 8427
rect 10789 8393 10828 8427
rect 10862 8393 10901 8427
rect 10935 8393 10974 8427
rect 11008 8393 11047 8427
rect 11081 8393 11120 8427
rect 11154 8393 11193 8427
rect 11227 8393 11266 8427
rect 11300 8393 11339 8427
rect 11373 8393 11412 8427
rect 11446 8393 11485 8427
rect 11519 8393 11558 8427
rect 11592 8393 11631 8427
rect 11665 8393 11704 8427
rect 11738 8393 11777 8427
rect 11811 8393 11850 8427
rect 11884 8393 11923 8427
rect 11957 8393 11996 8427
rect 12030 8393 12069 8427
rect 12103 8393 12142 8427
rect 12176 8393 12215 8427
rect 12249 8393 12288 8427
rect 12322 8393 12361 8427
rect 12395 8393 12434 8427
rect 12468 8393 12507 8427
rect 12541 8393 12580 8427
rect 12614 8393 12653 8427
rect 12687 8393 12726 8427
rect 12760 8393 12799 8427
rect 12833 8393 12872 8427
rect 12906 8393 12945 8427
rect 12979 8393 13018 8427
rect 13052 8393 13091 8427
rect 13701 8427 13779 8499
tri 14641 8470 14676 8505 ne
rect 13701 8393 13739 8427
rect 13773 8393 13779 8427
rect 10498 8392 13163 8393
rect 10458 8373 13163 8392
rect 10458 8355 11204 8373
rect 11256 8355 11274 8373
rect 11326 8355 11344 8373
rect 11396 8355 11414 8373
rect 10458 8353 10608 8355
rect 10458 8319 10464 8353
rect 10498 8319 10536 8353
rect 10570 8321 10608 8353
rect 10642 8321 10681 8355
rect 10715 8321 10754 8355
rect 10788 8321 10827 8355
rect 10861 8321 10900 8355
rect 10934 8321 10973 8355
rect 11007 8321 11046 8355
rect 11080 8321 11119 8355
rect 11153 8321 11192 8355
rect 11256 8321 11265 8355
rect 11326 8321 11338 8355
rect 11396 8321 11411 8355
rect 11466 8321 11483 8373
rect 11535 8321 11552 8373
rect 11604 8321 11621 8373
rect 11673 8321 11690 8373
rect 11742 8321 11759 8373
rect 11811 8321 11828 8373
rect 11880 8355 11897 8373
rect 11949 8355 13163 8373
rect 11883 8321 11897 8355
rect 11956 8321 11995 8355
rect 12029 8321 12068 8355
rect 12102 8321 12141 8355
rect 12175 8321 12214 8355
rect 12248 8321 12287 8355
rect 12321 8321 12360 8355
rect 12394 8321 12433 8355
rect 12467 8321 12506 8355
rect 12540 8321 12579 8355
rect 12613 8321 12652 8355
rect 12686 8321 12725 8355
rect 12759 8321 12798 8355
rect 12832 8321 12871 8355
rect 12905 8321 12944 8355
rect 12978 8321 13017 8355
rect 13051 8321 13090 8355
rect 13124 8321 13163 8355
rect 13557 8326 13779 8393
rect 13557 8321 13595 8326
rect 10570 8319 13595 8321
rect 10458 8315 13595 8319
rect 10458 8292 10677 8315
tri 10677 8292 10700 8315 nw
tri 13537 8292 13560 8315 ne
rect 13560 8292 13595 8315
rect 13629 8297 13779 8326
rect 13629 8292 13667 8297
rect 10458 8282 10648 8292
rect 10458 8280 10608 8282
rect 10458 8246 10464 8280
rect 10498 8246 10536 8280
rect 10570 8248 10608 8280
rect 10642 8248 10648 8282
tri 10648 8263 10677 8292 nw
tri 13560 8263 13589 8292 ne
rect 13589 8263 13667 8292
rect 13701 8263 13739 8297
rect 13773 8263 13779 8297
rect 13589 8251 13779 8263
rect 10570 8246 10648 8248
rect 10458 8209 10648 8246
tri 14642 8210 14676 8244 se
rect 14676 8210 14724 8505
rect 10458 8207 10608 8209
rect 10458 8173 10464 8207
rect 10498 8173 10536 8207
rect 10570 8175 10608 8207
rect 10642 8175 10648 8209
rect 10570 8173 10648 8175
rect 10458 8136 10648 8173
rect 10458 8134 10608 8136
rect 10458 8100 10464 8134
rect 10498 8100 10536 8134
rect 10570 8102 10608 8134
rect 10642 8102 10648 8136
rect 10570 8100 10648 8102
rect 10458 8063 10648 8100
rect 10458 8061 10608 8063
rect 10458 8027 10464 8061
rect 10498 8027 10536 8061
rect 10570 8029 10608 8061
rect 10642 8029 10648 8063
rect 10570 8027 10648 8029
rect 10458 7990 10648 8027
rect 10458 7988 10608 7990
rect 10458 7954 10464 7988
rect 10498 7954 10536 7988
rect 10570 7956 10608 7988
rect 10642 7956 10648 7990
rect 10570 7954 10648 7956
rect 620 7917 9646 7923
rect 620 7914 698 7917
rect 732 7914 771 7917
rect 805 7914 844 7917
rect 878 7914 917 7917
rect 951 7914 990 7917
rect 1024 7914 1063 7917
rect 1097 7914 1136 7917
rect 1170 7914 1209 7917
rect 1243 7914 1282 7917
rect 1316 7914 1355 7917
rect 1389 7914 1428 7917
rect 1462 7914 1501 7917
rect 1535 7914 1574 7917
rect 1608 7914 1647 7917
rect 1681 7914 1720 7917
rect 1754 7914 1793 7917
rect 1827 7914 1866 7917
rect 1900 7914 1939 7917
rect 1973 7914 2012 7917
rect 2046 7914 2085 7917
rect 2119 7914 2158 7917
rect 2192 7914 2231 7917
rect 2265 7914 2304 7917
rect 2338 7914 2377 7917
rect 2411 7914 2450 7917
rect 2484 7914 2523 7917
rect 2557 7914 2596 7917
rect 2630 7914 2669 7917
rect 2703 7914 2742 7917
rect 2776 7914 2815 7917
rect 2849 7914 2888 7917
rect 2922 7914 2961 7917
rect 2995 7914 3034 7917
rect 3068 7914 3107 7917
rect 3141 7914 3180 7917
rect 3214 7914 3253 7917
rect 3287 7914 3326 7917
rect 3360 7914 3399 7917
rect 3433 7914 3472 7917
rect 3506 7914 3545 7917
rect 3579 7914 3618 7917
rect 620 7862 695 7914
rect 747 7862 761 7914
rect 813 7862 827 7914
rect 879 7862 893 7914
rect 951 7883 959 7914
rect 1024 7883 1025 7914
rect 1275 7883 1282 7914
rect 945 7862 959 7883
rect 1011 7862 1025 7883
rect 1077 7862 1091 7883
rect 1143 7862 1157 7883
rect 1209 7862 1223 7883
rect 1275 7862 1289 7883
rect 1341 7862 1355 7914
rect 1407 7862 1421 7914
rect 1473 7862 1487 7914
rect 1539 7862 1553 7914
rect 1608 7883 1619 7914
rect 1681 7883 1684 7914
rect 1931 7883 1939 7914
rect 1605 7862 1619 7883
rect 1671 7862 1684 7883
rect 1736 7862 1749 7883
rect 1801 7862 1814 7883
rect 1866 7862 1879 7883
rect 1931 7862 1944 7883
rect 1996 7862 2009 7914
rect 2061 7862 2074 7914
rect 2126 7862 2139 7914
rect 2192 7883 2204 7914
rect 2265 7883 2269 7914
rect 2516 7883 2523 7914
rect 2191 7862 2204 7883
rect 2256 7862 2269 7883
rect 2321 7862 2334 7883
rect 2386 7862 2399 7883
rect 2451 7862 2464 7883
rect 2516 7862 2529 7883
rect 2581 7862 2594 7914
rect 2646 7862 2659 7914
rect 2711 7862 2724 7914
rect 2776 7862 2789 7914
rect 2849 7883 2854 7914
rect 3101 7883 3107 7914
rect 2841 7862 2854 7883
rect 2906 7862 2919 7883
rect 2971 7862 2984 7883
rect 3036 7862 3049 7883
rect 3101 7862 3114 7883
rect 3166 7862 3179 7914
rect 3231 7862 3244 7914
rect 3296 7862 3309 7914
rect 3361 7862 3374 7914
rect 3433 7883 3439 7914
rect 3652 7883 3691 7917
rect 3725 7883 3764 7917
rect 3798 7883 3837 7917
rect 3871 7883 3910 7917
rect 3944 7883 3983 7917
rect 4017 7883 4056 7917
rect 4090 7883 4129 7917
rect 4163 7883 4202 7917
rect 4236 7883 4275 7917
rect 4309 7883 4348 7917
rect 4382 7883 4421 7917
rect 4455 7883 4494 7917
rect 3426 7862 3439 7883
rect 3491 7862 3504 7883
rect 3556 7862 3569 7883
rect 3621 7862 4494 7883
rect 620 7850 4494 7862
rect 620 7845 631 7850
rect 683 7845 4494 7850
rect 620 6011 626 7845
rect 732 7811 771 7845
rect 805 7811 844 7845
rect 878 7811 917 7845
rect 951 7811 990 7845
rect 1024 7811 1063 7845
rect 1097 7811 1136 7845
rect 1170 7811 1209 7845
rect 1243 7811 1282 7845
rect 1316 7811 1355 7845
rect 1389 7811 1428 7845
rect 1462 7811 1501 7845
rect 1535 7811 1574 7845
rect 1608 7811 1647 7845
rect 1681 7811 1720 7845
rect 1754 7811 1793 7845
rect 1827 7811 1866 7845
rect 1900 7811 1939 7845
rect 1973 7811 2012 7845
rect 2046 7811 2085 7845
rect 2119 7811 2158 7845
rect 2192 7811 2231 7845
rect 2265 7811 2304 7845
rect 2338 7811 2377 7845
rect 2411 7811 2450 7845
rect 2484 7811 2523 7845
rect 2557 7811 2596 7845
rect 2630 7811 2669 7845
rect 2703 7811 2742 7845
rect 2776 7811 2815 7845
rect 2849 7811 2888 7845
rect 2922 7811 2961 7845
rect 2995 7811 3034 7845
rect 3068 7811 3107 7845
rect 3141 7811 3180 7845
rect 3214 7811 3253 7845
rect 3287 7811 3326 7845
rect 3360 7811 3399 7845
rect 3433 7811 3472 7845
rect 3506 7811 3545 7845
rect 3579 7811 3618 7845
rect 3652 7811 3691 7845
rect 3725 7811 3764 7845
rect 3798 7811 3837 7845
rect 3871 7811 3910 7845
rect 3944 7811 3983 7845
rect 4017 7811 4056 7845
rect 4090 7811 4129 7845
rect 4163 7811 4202 7845
rect 4236 7811 4275 7845
rect 4309 7811 4348 7845
rect 4382 7811 4421 7845
rect 4455 7811 4494 7845
rect 9568 7845 9646 7917
rect 9568 7811 9606 7845
rect 9640 7811 9646 7845
rect 732 7796 4566 7811
rect 732 7773 749 7796
rect 801 7773 814 7796
rect 866 7773 879 7796
rect 931 7773 944 7796
rect 996 7773 1009 7796
rect 1061 7773 1073 7796
rect 1125 7773 1137 7796
rect 804 7744 814 7773
rect 877 7744 879 7773
rect 1061 7744 1062 7773
rect 1125 7744 1135 7773
rect 1189 7744 1201 7796
rect 1253 7744 1265 7796
rect 1317 7744 1329 7796
rect 1381 7773 1393 7796
rect 1445 7773 1457 7796
rect 1509 7773 1521 7796
rect 1573 7773 1585 7796
rect 1637 7773 1649 7796
rect 1388 7744 1393 7773
rect 1637 7744 1646 7773
rect 1701 7744 1713 7796
rect 1765 7744 1777 7796
rect 1829 7744 1841 7796
rect 1893 7773 1905 7796
rect 1957 7773 1969 7796
rect 2021 7773 2033 7796
rect 2085 7773 2097 7796
rect 2149 7773 2161 7796
rect 1899 7744 1905 7773
rect 2149 7744 2157 7773
rect 2213 7744 2225 7796
rect 2277 7744 2289 7796
rect 2341 7744 2353 7796
rect 2405 7773 2417 7796
rect 2469 7773 2481 7796
rect 2533 7773 2545 7796
rect 2597 7773 2609 7796
rect 2661 7773 2673 7796
rect 2410 7744 2417 7773
rect 2661 7744 2668 7773
rect 2725 7744 2737 7796
rect 2789 7744 2801 7796
rect 2853 7744 2865 7796
rect 2917 7773 2929 7796
rect 2981 7773 2993 7796
rect 3045 7773 3057 7796
rect 3109 7773 3121 7796
rect 3173 7773 3185 7796
rect 2921 7744 2929 7773
rect 3173 7744 3179 7773
rect 3237 7744 3249 7796
rect 3301 7744 3313 7796
rect 3365 7744 3377 7796
rect 3429 7773 3441 7796
rect 3493 7773 3505 7796
rect 3557 7773 3569 7796
rect 3621 7773 4566 7796
rect 3432 7744 3441 7773
rect 804 7739 843 7744
rect 877 7739 916 7744
rect 950 7739 989 7744
rect 1023 7739 1062 7744
rect 1096 7739 1135 7744
rect 1169 7739 1208 7744
rect 1242 7739 1281 7744
rect 1315 7739 1354 7744
rect 1388 7739 1427 7744
rect 1461 7739 1500 7744
rect 1534 7739 1573 7744
rect 1607 7739 1646 7744
rect 1680 7739 1719 7744
rect 1753 7739 1792 7744
rect 1826 7739 1865 7744
rect 1899 7739 1938 7744
rect 1972 7739 2011 7744
rect 2045 7739 2084 7744
rect 2118 7739 2157 7744
rect 2191 7739 2230 7744
rect 2264 7739 2303 7744
rect 2337 7739 2376 7744
rect 2410 7739 2449 7744
rect 2483 7739 2522 7744
rect 2556 7739 2595 7744
rect 2629 7739 2668 7744
rect 2702 7739 2741 7744
rect 2775 7739 2814 7744
rect 2848 7739 2887 7744
rect 2921 7739 2960 7744
rect 2994 7739 3033 7744
rect 3067 7739 3106 7744
rect 3140 7739 3179 7744
rect 3213 7739 3252 7744
rect 3286 7739 3325 7744
rect 3359 7739 3398 7744
rect 3432 7739 3471 7744
rect 3505 7739 3544 7744
rect 3578 7739 3617 7744
rect 3651 7739 3690 7773
rect 3724 7739 3763 7773
rect 3797 7739 3836 7773
rect 3870 7739 3909 7773
rect 3943 7739 3982 7773
rect 4016 7739 4055 7773
rect 4089 7739 4128 7773
rect 4162 7739 4201 7773
rect 4235 7739 4274 7773
rect 4308 7739 4347 7773
rect 4381 7739 4420 7773
rect 4454 7739 4493 7773
rect 4527 7739 4566 7773
rect 9496 7771 9646 7811
rect 9496 7739 9534 7771
rect 804 7737 9534 7739
rect 9568 7737 9606 7771
rect 9640 7737 9646 7771
rect 804 7733 9646 7737
rect 804 7712 836 7733
tri 836 7712 857 7733 nw
tri 9402 7712 9423 7733 ne
rect 9423 7712 9646 7733
rect 804 7710 834 7712
tri 834 7710 836 7712 nw
tri 9423 7710 9425 7712 ne
rect 9425 7710 9646 7712
rect 804 7699 823 7710
tri 823 7699 834 7710 nw
tri 9425 7699 9436 7710 ne
rect 9436 7699 9646 7710
rect 804 6083 810 7699
tri 810 7686 823 7699 nw
tri 9436 7686 9449 7699 ne
rect 9449 7686 9462 7699
tri 9449 7679 9456 7686 ne
rect 9456 7665 9462 7686
rect 9496 7697 9646 7699
rect 9496 7665 9534 7697
rect 9456 7663 9534 7665
rect 9568 7663 9606 7697
rect 9640 7663 9646 7697
rect 9456 7625 9646 7663
rect 9456 7591 9462 7625
rect 9496 7623 9646 7625
rect 9496 7591 9534 7623
rect 9456 7589 9534 7591
rect 9568 7589 9606 7623
rect 9640 7589 9646 7623
rect 9456 7551 9646 7589
rect 732 6061 749 6083
rect 801 6061 810 6083
rect 732 6048 810 6061
rect 732 6011 749 6048
rect 801 6044 810 6048
rect 620 6006 631 6011
rect 683 6006 749 6011
rect 804 6010 810 6044
rect 620 5996 749 6006
rect 801 5996 810 6010
rect 620 5994 810 5996
rect 620 5972 631 5994
rect 683 5983 810 5994
rect 683 5972 749 5983
rect 620 5938 626 5972
rect 683 5942 698 5972
rect 660 5938 698 5942
rect 732 5938 749 5972
rect 801 5971 810 5983
rect 620 5931 749 5938
rect 804 5937 810 5971
rect 801 5931 810 5937
rect 620 5929 810 5931
rect 620 5899 631 5929
rect 683 5918 810 5929
rect 683 5899 749 5918
rect 620 5865 626 5899
rect 683 5877 698 5899
rect 660 5865 698 5877
rect 732 5866 749 5899
rect 801 5898 810 5918
rect 732 5865 770 5866
rect 620 5864 770 5865
rect 804 5864 810 5898
rect 620 5826 631 5864
rect 683 5853 810 5864
rect 683 5826 749 5853
rect 620 5792 626 5826
rect 683 5812 698 5826
rect 660 5799 698 5812
rect 683 5792 698 5799
rect 732 5801 749 5826
rect 801 5825 810 5853
rect 941 7519 9197 7525
rect 941 7485 1019 7519
rect 1053 7485 1091 7519
rect 1125 7485 1163 7519
rect 1197 7485 1235 7519
rect 1269 7485 1307 7519
rect 1341 7485 1379 7519
rect 1413 7485 1451 7519
rect 1485 7485 1523 7519
rect 1557 7485 1595 7519
rect 1629 7485 1667 7519
rect 1701 7485 1739 7519
rect 1773 7485 1811 7519
rect 1845 7485 1883 7519
rect 1917 7485 1955 7519
rect 1989 7485 2027 7519
rect 2061 7485 2099 7519
rect 2133 7485 2171 7519
rect 2205 7485 2243 7519
rect 2277 7485 2315 7519
rect 2349 7485 2387 7519
rect 2421 7485 2459 7519
rect 2493 7485 2531 7519
rect 2565 7485 2603 7519
rect 2637 7485 2675 7519
rect 2709 7485 2747 7519
rect 2781 7485 2819 7519
rect 2853 7485 2891 7519
rect 2925 7485 2963 7519
rect 2997 7485 3035 7519
rect 3069 7485 3107 7519
rect 3141 7485 3179 7519
rect 3213 7485 3251 7519
rect 3285 7485 3323 7519
rect 3357 7485 3395 7519
rect 3429 7485 3467 7519
rect 3501 7485 3539 7519
rect 3573 7485 3611 7519
rect 3645 7485 3683 7519
rect 3717 7485 3755 7519
rect 3789 7485 3827 7519
rect 3861 7485 3899 7519
rect 3933 7485 3971 7519
rect 4005 7485 4043 7519
rect 4077 7485 4115 7519
rect 4149 7485 4187 7519
rect 4221 7485 4259 7519
rect 4293 7485 4331 7519
rect 4365 7485 4403 7519
rect 4437 7485 4475 7519
rect 4509 7485 4547 7519
rect 4581 7485 4619 7519
rect 4653 7485 4691 7519
rect 4725 7485 4763 7519
rect 4797 7485 4835 7519
rect 4869 7485 4907 7519
rect 4941 7485 4979 7519
rect 5013 7485 5051 7519
rect 5085 7485 5123 7519
rect 5157 7485 5195 7519
rect 5229 7485 5267 7519
rect 5301 7485 5339 7519
rect 5373 7485 5411 7519
rect 5445 7485 5483 7519
rect 5517 7485 5555 7519
rect 5589 7485 5627 7519
rect 5661 7485 5699 7519
rect 5733 7485 5771 7519
rect 5805 7485 5843 7519
rect 5877 7485 5915 7519
rect 5949 7485 5987 7519
rect 6021 7485 6059 7519
rect 6093 7485 6131 7519
rect 6165 7485 6203 7519
rect 6237 7485 6275 7519
rect 6309 7485 6347 7519
rect 6381 7485 6419 7519
rect 6453 7485 6491 7519
rect 6525 7485 6563 7519
rect 6597 7485 6635 7519
rect 6669 7485 6707 7519
rect 6741 7485 6779 7519
rect 6813 7485 6851 7519
rect 6885 7485 6923 7519
rect 6957 7485 6995 7519
rect 7029 7485 7067 7519
rect 7101 7485 7139 7519
rect 7173 7485 7211 7519
rect 7245 7485 7283 7519
rect 7317 7485 7355 7519
rect 7389 7485 7427 7519
rect 7461 7485 7499 7519
rect 7533 7485 7571 7519
rect 7605 7485 7643 7519
rect 7677 7485 7715 7519
rect 7749 7485 7787 7519
rect 7821 7485 7859 7519
rect 7893 7485 7931 7519
rect 7965 7485 8003 7519
rect 8037 7485 8075 7519
rect 8109 7485 8147 7519
rect 8181 7485 8219 7519
rect 8253 7485 8291 7519
rect 8325 7485 8363 7519
rect 8397 7485 8435 7519
rect 8469 7485 8507 7519
rect 8541 7485 8579 7519
rect 8613 7485 8651 7519
rect 8685 7485 8723 7519
rect 8757 7485 8795 7519
rect 8829 7485 8867 7519
rect 8901 7485 8939 7519
rect 8973 7485 9012 7519
rect 9046 7485 9085 7519
rect 9119 7485 9197 7519
rect 941 7479 9197 7485
rect 941 7477 1025 7479
tri 1025 7477 1027 7479 nw
tri 9121 7477 9123 7479 ne
rect 9123 7477 9197 7479
rect 941 7447 993 7477
rect 941 7413 947 7447
rect 981 7445 993 7447
tri 993 7445 1025 7477 nw
tri 9123 7449 9151 7477 ne
rect 9151 7445 9197 7477
rect 981 7413 987 7445
tri 987 7439 993 7445 nw
rect 941 7372 987 7413
rect 1257 7428 8895 7434
rect 1257 7394 1269 7428
rect 1303 7394 1342 7428
rect 1376 7394 1415 7428
rect 1449 7394 1488 7428
rect 1522 7394 1561 7428
rect 1595 7394 1634 7428
rect 1668 7394 1707 7428
rect 1741 7394 1780 7428
rect 1814 7394 1853 7428
rect 1887 7394 1926 7428
rect 1960 7394 1999 7428
rect 2033 7394 2072 7428
rect 2106 7394 2145 7428
rect 2179 7394 2218 7428
rect 2252 7394 2291 7428
rect 2325 7394 2364 7428
rect 2398 7394 2437 7428
rect 2471 7394 2510 7428
rect 2544 7394 2583 7428
rect 2617 7394 2656 7428
rect 2690 7394 2729 7428
rect 2763 7394 2802 7428
rect 2836 7394 2875 7428
rect 2909 7394 2948 7428
rect 2982 7394 3021 7428
rect 3055 7394 3094 7428
rect 3128 7394 3167 7428
rect 3201 7394 3240 7428
rect 3274 7394 3313 7428
rect 3347 7394 3386 7428
rect 3420 7394 3459 7428
rect 3493 7394 3532 7428
rect 3566 7394 3605 7428
rect 3639 7394 3678 7428
rect 3712 7394 3751 7428
rect 3785 7394 3824 7428
rect 3858 7394 3897 7428
rect 3931 7394 3970 7428
rect 4004 7394 4043 7428
rect 4077 7394 4116 7428
rect 4150 7394 4189 7428
rect 4223 7394 4262 7428
rect 4296 7394 4335 7428
rect 4369 7394 4408 7428
rect 4442 7394 4481 7428
rect 4515 7394 4554 7428
rect 4588 7394 4627 7428
rect 4661 7394 4700 7428
rect 4734 7394 4773 7428
rect 4807 7394 4846 7428
rect 4880 7394 4919 7428
rect 4953 7394 4992 7428
rect 5026 7394 5065 7428
rect 5099 7394 5138 7428
rect 5172 7394 5211 7428
rect 5245 7394 5284 7428
rect 5318 7394 5357 7428
rect 5391 7394 5430 7428
rect 5464 7394 5503 7428
rect 5537 7394 5576 7428
rect 5610 7394 5649 7428
rect 5683 7394 5722 7428
rect 5756 7394 5795 7428
rect 5829 7394 5868 7428
rect 5902 7394 5941 7428
rect 5975 7394 6014 7428
rect 6048 7394 6087 7428
rect 6121 7394 6160 7428
rect 6194 7394 6233 7428
rect 6267 7394 6306 7428
rect 6340 7394 6379 7428
rect 6413 7394 6451 7428
rect 6485 7394 6523 7428
rect 6557 7394 6595 7428
rect 6629 7394 6667 7428
rect 6701 7394 6739 7428
rect 6773 7394 6811 7428
rect 6845 7394 6883 7428
rect 6917 7394 6955 7428
rect 6989 7394 7027 7428
rect 7061 7394 7099 7428
rect 7133 7394 7171 7428
rect 7205 7394 7243 7428
rect 7277 7394 7315 7428
rect 7349 7394 7387 7428
rect 7421 7394 7459 7428
rect 7493 7394 7531 7428
rect 7565 7394 7603 7428
rect 7637 7394 7675 7428
rect 7709 7394 7747 7428
rect 7781 7394 7819 7428
rect 7853 7394 7891 7428
rect 7925 7394 7963 7428
rect 7997 7394 8035 7428
rect 8069 7394 8107 7428
rect 8141 7394 8179 7428
rect 8213 7394 8251 7428
rect 8285 7394 8323 7428
rect 8357 7394 8395 7428
rect 8429 7394 8467 7428
rect 8501 7394 8539 7428
rect 8573 7394 8611 7428
rect 8645 7394 8683 7428
rect 8717 7394 8755 7428
rect 8789 7394 8827 7428
rect 8861 7394 8895 7428
rect 1257 7388 8895 7394
tri 8883 7382 8889 7388 ne
rect 8889 7382 8895 7388
rect 8947 7382 8959 7434
rect 9011 7382 9017 7434
rect 9151 7411 9157 7445
rect 9191 7411 9197 7445
rect 941 7338 947 7372
rect 981 7338 987 7372
rect 9151 7371 9197 7411
rect 941 7337 987 7338
tri 987 7337 994 7344 sw
tri 9144 7337 9151 7344 se
rect 9151 7337 9157 7371
rect 9191 7337 9197 7371
rect 941 7333 994 7337
tri 994 7333 998 7337 sw
tri 9140 7333 9144 7337 se
rect 9144 7333 9197 7337
rect 941 7331 998 7333
tri 998 7331 1000 7333 sw
tri 9138 7331 9140 7333 se
rect 9140 7331 9197 7333
rect 941 7329 1000 7331
tri 1000 7329 1002 7331 sw
tri 9136 7329 9138 7331 se
rect 9138 7329 9197 7331
rect 941 7310 1002 7329
tri 1002 7310 1021 7329 sw
tri 9117 7310 9136 7329 se
rect 9136 7310 9197 7329
rect 941 7298 9197 7310
rect 941 7297 1223 7298
rect 941 7263 947 7297
rect 981 7264 1223 7297
rect 1257 7264 1535 7298
rect 1569 7264 1847 7298
rect 1881 7264 2159 7298
rect 2193 7264 2471 7298
rect 2505 7264 2783 7298
rect 2817 7264 3095 7298
rect 3129 7264 3407 7298
rect 3441 7295 3719 7298
rect 3753 7295 4031 7298
rect 4065 7295 4343 7298
rect 4377 7295 4655 7298
rect 4689 7295 4967 7298
rect 5001 7295 5279 7298
rect 5313 7295 5591 7298
rect 5625 7295 5903 7298
rect 5937 7295 6215 7298
rect 6249 7295 6527 7298
rect 6561 7295 6839 7298
rect 6873 7295 7151 7298
rect 7185 7295 7463 7298
rect 7497 7295 7775 7298
rect 7809 7295 8087 7298
rect 8121 7295 8399 7298
rect 8433 7295 8711 7298
rect 8745 7295 9023 7298
rect 9057 7297 9197 7298
rect 9057 7295 9157 7297
rect 3441 7264 3446 7295
rect 981 7263 3446 7264
rect 941 7243 3446 7263
rect 3498 7243 3511 7295
rect 3563 7243 3576 7295
rect 3628 7243 3641 7295
rect 3693 7243 3706 7295
rect 3758 7243 3771 7295
rect 3823 7243 3836 7295
rect 3888 7243 3901 7295
rect 3953 7243 3966 7295
rect 4018 7243 4031 7295
rect 4083 7243 4096 7295
rect 4148 7243 4161 7295
rect 4213 7243 4226 7295
rect 4278 7243 4291 7295
rect 4343 7243 4356 7264
rect 4408 7243 4421 7295
rect 4473 7243 4486 7295
rect 4538 7243 4551 7295
rect 4603 7243 4616 7295
rect 4668 7243 4681 7264
rect 4733 7243 4746 7295
rect 4798 7243 4811 7295
rect 4863 7243 4876 7295
rect 4928 7243 4941 7295
rect 5001 7264 5006 7295
rect 4993 7243 5006 7264
rect 5058 7243 5071 7295
rect 5123 7243 5136 7295
rect 5188 7243 5201 7295
rect 5253 7243 5266 7295
rect 5318 7243 5331 7295
rect 5383 7243 5396 7295
rect 5448 7243 5461 7295
rect 5513 7243 5526 7295
rect 5578 7243 5591 7295
rect 941 7231 5591 7243
rect 941 7224 3446 7231
rect 941 7222 1223 7224
rect 941 7188 947 7222
rect 981 7190 1223 7222
rect 1257 7190 1535 7224
rect 1569 7190 1847 7224
rect 1881 7190 2159 7224
rect 2193 7190 2471 7224
rect 2505 7190 2783 7224
rect 2817 7190 3095 7224
rect 3129 7190 3407 7224
rect 3441 7190 3446 7224
rect 981 7188 3446 7190
rect 941 7179 3446 7188
rect 3498 7179 3511 7231
rect 3563 7179 3576 7231
rect 3628 7179 3641 7231
rect 3693 7179 3706 7231
rect 3758 7179 3771 7231
rect 3823 7179 3836 7231
rect 3888 7179 3901 7231
rect 3953 7179 3966 7231
rect 4018 7179 4031 7231
rect 4083 7179 4096 7231
rect 4148 7179 4161 7231
rect 4213 7179 4226 7231
rect 4278 7179 4291 7231
rect 4343 7224 4356 7231
rect 4343 7179 4356 7190
rect 4408 7179 4421 7231
rect 4473 7179 4486 7231
rect 4538 7179 4551 7231
rect 4603 7179 4616 7231
rect 4668 7224 4681 7231
rect 4668 7179 4681 7190
rect 4733 7179 4746 7231
rect 4798 7179 4811 7231
rect 4863 7179 4876 7231
rect 4928 7179 4941 7231
rect 4993 7224 5006 7231
rect 5001 7190 5006 7224
rect 4993 7179 5006 7190
rect 5058 7179 5071 7231
rect 5123 7179 5136 7231
rect 5188 7179 5201 7231
rect 5253 7179 5266 7231
rect 5318 7179 5331 7231
rect 5383 7179 5396 7231
rect 5448 7179 5461 7231
rect 5513 7179 5526 7231
rect 5578 7179 5591 7231
rect 9099 7263 9157 7295
rect 9191 7263 9197 7297
rect 9099 7223 9197 7263
rect 941 7167 5591 7179
rect 941 7150 3446 7167
rect 941 7147 1223 7150
rect 941 7113 947 7147
rect 981 7116 1223 7147
rect 1257 7116 1535 7150
rect 1569 7116 1847 7150
rect 1881 7116 2159 7150
rect 2193 7116 2471 7150
rect 2505 7116 2783 7150
rect 2817 7116 3095 7150
rect 3129 7116 3407 7150
rect 3441 7116 3446 7150
rect 981 7115 3446 7116
rect 3498 7115 3511 7167
rect 3563 7115 3576 7167
rect 3628 7115 3641 7167
rect 3693 7115 3706 7167
rect 3758 7115 3771 7167
rect 3823 7115 3836 7167
rect 3888 7115 3901 7167
rect 3953 7115 3966 7167
rect 4018 7115 4031 7167
rect 4083 7115 4096 7167
rect 4148 7115 4161 7167
rect 4213 7115 4226 7167
rect 4278 7115 4291 7167
rect 4343 7150 4356 7167
rect 4343 7115 4356 7116
rect 4408 7115 4421 7167
rect 4473 7115 4486 7167
rect 4538 7115 4551 7167
rect 4603 7115 4616 7167
rect 4668 7150 4681 7167
rect 4668 7115 4681 7116
rect 4733 7115 4746 7167
rect 4798 7115 4811 7167
rect 4863 7115 4876 7167
rect 4928 7115 4941 7167
rect 4993 7150 5006 7167
rect 5001 7116 5006 7150
rect 4993 7115 5006 7116
rect 5058 7115 5071 7167
rect 5123 7115 5136 7167
rect 5188 7115 5201 7167
rect 5253 7115 5266 7167
rect 5318 7115 5331 7167
rect 5383 7115 5396 7167
rect 5448 7115 5461 7167
rect 5513 7115 5526 7167
rect 5578 7115 5591 7167
rect 9099 7189 9157 7223
rect 9191 7189 9197 7223
rect 9099 7149 9197 7189
rect 981 7113 5591 7115
rect 941 7103 5591 7113
rect 941 7076 3446 7103
rect 941 7072 1223 7076
rect 941 7038 947 7072
rect 981 7042 1223 7072
rect 1257 7042 1535 7076
rect 1569 7042 1847 7076
rect 1881 7042 2159 7076
rect 2193 7042 2471 7076
rect 2505 7042 2783 7076
rect 2817 7042 3095 7076
rect 3129 7042 3407 7076
rect 3441 7051 3446 7076
rect 3498 7051 3511 7103
rect 3563 7051 3576 7103
rect 3628 7051 3641 7103
rect 3693 7051 3706 7103
rect 3758 7051 3771 7103
rect 3823 7051 3836 7103
rect 3888 7051 3901 7103
rect 3953 7051 3966 7103
rect 4018 7051 4031 7103
rect 4083 7051 4096 7103
rect 4148 7051 4161 7103
rect 4213 7051 4226 7103
rect 4278 7051 4291 7103
rect 4343 7076 4356 7103
rect 4408 7051 4421 7103
rect 4473 7051 4486 7103
rect 4538 7051 4551 7103
rect 4603 7051 4616 7103
rect 4668 7076 4681 7103
rect 4733 7051 4746 7103
rect 4798 7051 4811 7103
rect 4863 7051 4876 7103
rect 4928 7051 4941 7103
rect 4993 7076 5006 7103
rect 5001 7051 5006 7076
rect 5058 7051 5071 7103
rect 5123 7051 5136 7103
rect 5188 7051 5201 7103
rect 5253 7051 5266 7103
rect 5318 7051 5331 7103
rect 5383 7051 5396 7103
rect 5448 7051 5461 7103
rect 5513 7051 5526 7103
rect 5578 7051 5591 7103
rect 9099 7115 9157 7149
rect 9191 7115 9197 7149
rect 3441 7042 3719 7051
rect 3753 7042 4031 7051
rect 4065 7042 4343 7051
rect 4377 7042 4655 7051
rect 4689 7042 4967 7051
rect 5001 7042 5279 7051
rect 5313 7042 5591 7051
rect 9099 7075 9197 7115
rect 981 7039 5591 7042
rect 981 7038 3446 7039
rect 941 7002 3446 7038
rect 941 6997 1223 7002
rect 941 6963 947 6997
rect 981 6968 1223 6997
rect 1257 7001 1847 7002
rect 1257 6968 1535 7001
rect 981 6967 1535 6968
rect 1569 6968 1847 7001
rect 1881 7001 2471 7002
rect 1881 6968 2159 7001
rect 1569 6967 2159 6968
rect 2193 6968 2471 7001
rect 2505 7001 3095 7002
rect 2505 6968 2783 7001
rect 2193 6967 2783 6968
rect 2817 6968 3095 7001
rect 3129 7001 3446 7002
rect 3129 6968 3407 7001
rect 2817 6967 3407 6968
rect 3441 6987 3446 7001
rect 3498 6987 3511 7039
rect 3563 6987 3576 7039
rect 3628 6987 3641 7039
rect 3693 6987 3706 7039
rect 3758 6987 3771 7039
rect 3823 6987 3836 7039
rect 3888 6987 3901 7039
rect 3953 6987 3966 7039
rect 4018 6987 4031 7039
rect 4083 6987 4096 7039
rect 4148 6987 4161 7039
rect 4213 6987 4226 7039
rect 4278 6987 4291 7039
rect 4343 7002 4356 7039
rect 4408 6987 4421 7039
rect 4473 6987 4486 7039
rect 4538 6987 4551 7039
rect 4603 6987 4616 7039
rect 4668 7001 4681 7039
rect 4733 6987 4746 7039
rect 4798 6987 4811 7039
rect 4863 6987 4876 7039
rect 4928 6987 4941 7039
rect 4993 7002 5006 7039
rect 5001 6987 5006 7002
rect 5058 6987 5071 7039
rect 5123 6987 5136 7039
rect 5188 6987 5201 7039
rect 5253 6987 5266 7039
rect 5318 6987 5331 7039
rect 5383 6987 5396 7039
rect 5448 6987 5461 7039
rect 5513 6987 5526 7039
rect 5578 6987 5591 7039
rect 9099 7041 9157 7075
rect 9191 7041 9197 7075
rect 3441 6975 3719 6987
rect 3753 6975 4031 6987
rect 4065 6975 4343 6987
rect 4377 6975 4655 6987
rect 4689 6975 4967 6987
rect 5001 6975 5279 6987
rect 5313 6975 5591 6987
rect 3441 6967 3446 6975
rect 981 6963 3446 6967
rect 941 6927 3446 6963
rect 941 6922 1223 6927
rect 941 6888 947 6922
rect 981 6893 1223 6922
rect 1257 6926 1847 6927
rect 1257 6893 1535 6926
rect 981 6892 1535 6893
rect 1569 6893 1847 6926
rect 1881 6926 2471 6927
rect 1881 6893 2159 6926
rect 1569 6892 2159 6893
rect 2193 6893 2471 6926
rect 2505 6926 3095 6927
rect 2505 6893 2783 6926
rect 2193 6892 2783 6893
rect 2817 6893 3095 6926
rect 3129 6926 3446 6927
rect 3129 6893 3407 6926
rect 2817 6892 3407 6893
rect 3441 6923 3446 6926
rect 3498 6923 3511 6975
rect 3563 6923 3576 6975
rect 3628 6923 3641 6975
rect 3693 6923 3706 6975
rect 3758 6923 3771 6975
rect 3823 6923 3836 6975
rect 3888 6923 3901 6975
rect 3953 6923 3966 6975
rect 4018 6923 4031 6975
rect 4083 6923 4096 6975
rect 4148 6923 4161 6975
rect 4213 6923 4226 6975
rect 4278 6923 4291 6975
rect 4343 6927 4356 6968
rect 4408 6923 4421 6975
rect 4473 6923 4486 6975
rect 4538 6923 4551 6975
rect 4603 6923 4616 6975
rect 4668 6926 4681 6967
rect 4733 6923 4746 6975
rect 4798 6923 4811 6975
rect 4863 6923 4876 6975
rect 4928 6923 4941 6975
rect 5001 6968 5006 6975
rect 4993 6927 5006 6968
rect 5001 6923 5006 6927
rect 5058 6923 5071 6975
rect 5123 6923 5136 6975
rect 5188 6923 5201 6975
rect 5253 6923 5266 6975
rect 5318 6923 5331 6975
rect 5383 6923 5396 6975
rect 5448 6923 5461 6975
rect 5513 6923 5526 6975
rect 5578 6923 5591 6975
rect 9099 7001 9197 7041
rect 9099 6967 9157 7001
rect 9191 6967 9197 7001
rect 3441 6911 3719 6923
rect 3753 6911 4031 6923
rect 4065 6911 4343 6923
rect 4377 6911 4655 6923
rect 4689 6911 4967 6923
rect 5001 6911 5279 6923
rect 5313 6911 5591 6923
rect 3441 6892 3446 6911
rect 981 6888 3446 6892
rect 941 6859 3446 6888
rect 3498 6859 3511 6911
rect 3563 6859 3576 6911
rect 3628 6859 3641 6911
rect 3693 6859 3706 6911
rect 3758 6859 3771 6911
rect 3823 6859 3836 6911
rect 3888 6859 3901 6911
rect 3953 6859 3966 6911
rect 4018 6859 4031 6911
rect 4083 6859 4096 6911
rect 4148 6859 4161 6911
rect 4213 6859 4226 6911
rect 4278 6859 4291 6911
rect 4343 6859 4356 6893
rect 4408 6859 4421 6911
rect 4473 6859 4486 6911
rect 4538 6859 4551 6911
rect 4603 6859 4616 6911
rect 4668 6859 4681 6892
rect 4733 6859 4746 6911
rect 4798 6859 4811 6911
rect 4863 6859 4876 6911
rect 4928 6859 4941 6911
rect 5001 6893 5006 6911
rect 4993 6859 5006 6893
rect 5058 6859 5071 6911
rect 5123 6859 5136 6911
rect 5188 6859 5201 6911
rect 5253 6859 5266 6911
rect 5318 6859 5331 6911
rect 5383 6859 5396 6911
rect 5448 6859 5461 6911
rect 5513 6859 5526 6911
rect 5578 6859 5591 6911
rect 9099 6926 9197 6967
rect 9099 6892 9157 6926
rect 9191 6892 9197 6926
rect 941 6852 5591 6859
rect 941 6847 1223 6852
rect 941 6813 947 6847
rect 981 6818 1223 6847
rect 1257 6851 1847 6852
rect 1257 6818 1535 6851
rect 981 6817 1535 6818
rect 1569 6818 1847 6851
rect 1881 6851 2471 6852
rect 1881 6818 2159 6851
rect 1569 6817 2159 6818
rect 2193 6818 2471 6851
rect 2505 6851 3095 6852
rect 2505 6818 2783 6851
rect 2193 6817 2783 6818
rect 2817 6818 3095 6851
rect 3129 6851 3719 6852
rect 3129 6818 3407 6851
rect 2817 6817 3407 6818
rect 3441 6847 3719 6851
rect 3753 6851 4343 6852
rect 3753 6847 4031 6851
rect 4065 6847 4343 6851
rect 4377 6851 4967 6852
rect 4377 6847 4655 6851
rect 4689 6847 4967 6851
rect 5001 6851 5591 6852
rect 5001 6847 5279 6851
rect 5313 6847 5591 6851
rect 3441 6817 3446 6847
rect 981 6813 3446 6817
rect 941 6795 3446 6813
rect 3498 6795 3511 6847
rect 3563 6795 3576 6847
rect 3628 6795 3641 6847
rect 3693 6795 3706 6847
rect 3758 6795 3771 6847
rect 3823 6795 3836 6847
rect 3888 6795 3901 6847
rect 3953 6795 3966 6847
rect 4018 6795 4031 6847
rect 4083 6795 4096 6847
rect 4148 6795 4161 6847
rect 4213 6795 4226 6847
rect 4278 6795 4291 6847
rect 4343 6795 4356 6818
rect 4408 6795 4421 6847
rect 4473 6795 4486 6847
rect 4538 6795 4551 6847
rect 4603 6795 4616 6847
rect 4668 6795 4681 6817
rect 4733 6795 4746 6847
rect 4798 6795 4811 6847
rect 4863 6795 4876 6847
rect 4928 6795 4941 6847
rect 5001 6818 5006 6847
rect 4993 6795 5006 6818
rect 5058 6795 5071 6847
rect 5123 6795 5136 6847
rect 5188 6795 5201 6847
rect 5253 6795 5266 6847
rect 5318 6795 5331 6847
rect 5383 6795 5396 6847
rect 5448 6795 5461 6847
rect 5513 6795 5526 6847
rect 5578 6795 5591 6847
rect 9099 6851 9197 6892
rect 9099 6817 9157 6851
rect 9191 6817 9197 6851
rect 941 6783 5591 6795
rect 941 6777 3446 6783
rect 941 6772 1223 6777
rect 941 6738 947 6772
rect 981 6743 1223 6772
rect 1257 6776 1847 6777
rect 1257 6743 1535 6776
rect 981 6742 1535 6743
rect 1569 6743 1847 6776
rect 1881 6776 2471 6777
rect 1881 6743 2159 6776
rect 1569 6742 2159 6743
rect 2193 6743 2471 6776
rect 2505 6776 3095 6777
rect 2505 6743 2783 6776
rect 2193 6742 2783 6743
rect 2817 6743 3095 6776
rect 3129 6776 3446 6777
rect 3129 6743 3407 6776
rect 2817 6742 3407 6743
rect 3441 6742 3446 6776
rect 981 6738 3446 6742
rect 941 6731 3446 6738
rect 3498 6731 3511 6783
rect 3563 6731 3576 6783
rect 3628 6731 3641 6783
rect 3693 6731 3706 6783
rect 3758 6731 3771 6783
rect 3823 6731 3836 6783
rect 3888 6731 3901 6783
rect 3953 6731 3966 6783
rect 4018 6731 4031 6783
rect 4083 6731 4096 6783
rect 4148 6731 4161 6783
rect 4213 6731 4226 6783
rect 4278 6731 4291 6783
rect 4343 6777 4356 6783
rect 4343 6731 4356 6743
rect 4408 6731 4421 6783
rect 4473 6731 4486 6783
rect 4538 6731 4551 6783
rect 4603 6731 4616 6783
rect 4668 6776 4681 6783
rect 4668 6731 4681 6742
rect 4733 6731 4746 6783
rect 4798 6731 4811 6783
rect 4863 6731 4876 6783
rect 4928 6731 4941 6783
rect 4993 6777 5006 6783
rect 5001 6743 5006 6777
rect 4993 6731 5006 6743
rect 5058 6731 5071 6783
rect 5123 6731 5136 6783
rect 5188 6731 5201 6783
rect 5253 6731 5266 6783
rect 5318 6731 5331 6783
rect 5383 6731 5396 6783
rect 5448 6731 5461 6783
rect 5513 6731 5526 6783
rect 5578 6731 5591 6783
rect 9099 6776 9197 6817
rect 9099 6742 9157 6776
rect 9191 6742 9197 6776
rect 941 6719 5591 6731
rect 941 6702 3446 6719
rect 941 6697 1223 6702
rect 941 6663 947 6697
rect 981 6668 1223 6697
rect 1257 6701 1847 6702
rect 1257 6668 1535 6701
rect 981 6667 1535 6668
rect 1569 6668 1847 6701
rect 1881 6701 2471 6702
rect 1881 6668 2159 6701
rect 1569 6667 2159 6668
rect 2193 6668 2471 6701
rect 2505 6701 3095 6702
rect 2505 6668 2783 6701
rect 2193 6667 2783 6668
rect 2817 6668 3095 6701
rect 3129 6701 3446 6702
rect 3129 6668 3407 6701
rect 2817 6667 3407 6668
rect 3441 6667 3446 6701
rect 3498 6667 3511 6719
rect 3563 6667 3576 6719
rect 3628 6667 3641 6719
rect 3693 6667 3706 6719
rect 3758 6667 3771 6719
rect 3823 6667 3836 6719
rect 3888 6667 3901 6719
rect 3953 6667 3966 6719
rect 4018 6667 4031 6719
rect 4083 6667 4096 6719
rect 4148 6667 4161 6719
rect 4213 6667 4226 6719
rect 4278 6667 4291 6719
rect 4343 6702 4356 6719
rect 4343 6667 4356 6668
rect 4408 6667 4421 6719
rect 4473 6667 4486 6719
rect 4538 6667 4551 6719
rect 4603 6667 4616 6719
rect 4668 6701 4681 6719
rect 4733 6667 4746 6719
rect 4798 6667 4811 6719
rect 4863 6667 4876 6719
rect 4928 6667 4941 6719
rect 4993 6702 5006 6719
rect 5001 6668 5006 6702
rect 4993 6667 5006 6668
rect 5058 6667 5071 6719
rect 5123 6667 5136 6719
rect 5188 6667 5201 6719
rect 5253 6667 5266 6719
rect 5318 6667 5331 6719
rect 5383 6667 5396 6719
rect 5448 6667 5461 6719
rect 5513 6667 5526 6719
rect 5578 6667 5591 6719
rect 9099 6701 9197 6742
rect 9099 6667 9157 6701
rect 9191 6667 9197 6701
rect 981 6663 9197 6667
rect 941 6655 9197 6663
rect 941 6635 1001 6655
tri 1001 6635 1021 6655 nw
tri 9121 6635 9141 6655 ne
rect 9141 6635 9197 6655
rect 941 6633 999 6635
tri 999 6633 1001 6635 nw
tri 9141 6633 9143 6635 ne
rect 9143 6633 9197 6635
rect 941 6626 992 6633
tri 992 6626 999 6633 nw
tri 9143 6626 9150 6633 ne
rect 9150 6626 9197 6633
rect 941 6622 987 6626
rect 941 6588 947 6622
rect 981 6588 987 6622
tri 987 6621 992 6626 nw
tri 9150 6625 9151 6626 ne
rect 941 6547 987 6588
rect 9151 6592 9157 6626
rect 9191 6592 9197 6626
rect 941 6513 947 6547
rect 981 6513 987 6547
rect 941 6472 987 6513
rect 941 6438 947 6472
rect 981 6438 987 6472
rect 941 6398 987 6438
rect 941 6364 947 6398
rect 981 6364 987 6398
rect 941 6324 987 6364
rect 941 6290 947 6324
rect 981 6290 987 6324
rect 941 6250 987 6290
rect 941 6216 947 6250
rect 981 6216 987 6250
rect 941 6176 987 6216
rect 941 6142 947 6176
rect 981 6142 987 6176
rect 941 6102 987 6142
rect 941 6068 947 6102
rect 981 6068 987 6102
rect 941 6028 987 6068
rect 941 5994 947 6028
rect 981 5994 987 6028
rect 941 5954 987 5994
rect 941 5920 947 5954
rect 981 5920 987 5954
rect 1217 6578 9064 6584
rect 1217 6572 8941 6578
rect 1217 6538 1379 6572
rect 1413 6538 1691 6572
rect 1725 6538 2003 6572
rect 2037 6538 2315 6572
rect 2349 6538 2627 6572
rect 2661 6538 2939 6572
rect 2973 6538 3251 6572
rect 3285 6538 3563 6572
rect 3597 6570 3875 6572
rect 3909 6570 4187 6572
rect 3597 6538 3857 6570
rect 1217 6518 3857 6538
rect 3909 6518 3981 6570
rect 4033 6538 4187 6570
rect 4221 6538 4499 6572
rect 4533 6538 4811 6572
rect 4845 6538 5123 6572
rect 5157 6538 5435 6572
rect 5469 6538 5747 6572
rect 5781 6538 6059 6572
rect 6093 6538 6371 6572
rect 6405 6538 6683 6572
rect 6717 6538 6995 6572
rect 7029 6538 7307 6572
rect 7341 6538 7619 6572
rect 7653 6538 7931 6572
rect 7965 6538 8243 6572
rect 8277 6538 8555 6572
rect 8589 6538 8867 6572
rect 8901 6538 8941 6572
rect 4033 6526 8941 6538
rect 8993 6526 9011 6578
rect 9063 6526 9064 6578
rect 4033 6518 9064 6526
rect 1217 6514 9064 6518
rect 1217 6500 8941 6514
rect 1217 6466 1379 6500
rect 1413 6499 2003 6500
rect 1413 6466 1691 6499
rect 1217 6465 1691 6466
rect 1725 6466 2003 6499
rect 2037 6499 2627 6500
rect 2037 6466 2315 6499
rect 1725 6465 2315 6466
rect 2349 6466 2627 6499
rect 2661 6499 3857 6500
rect 2661 6466 2939 6499
rect 2349 6465 2939 6466
rect 2973 6465 3251 6499
rect 3285 6465 3563 6499
rect 3597 6465 3857 6499
rect 1217 6448 3857 6465
rect 3909 6448 3981 6500
rect 4033 6499 4499 6500
rect 4033 6465 4187 6499
rect 4221 6466 4499 6499
rect 4533 6499 5123 6500
rect 4533 6466 4811 6499
rect 4221 6465 4811 6466
rect 4845 6466 5123 6499
rect 5157 6499 5747 6500
rect 5157 6466 5435 6499
rect 4845 6465 5435 6466
rect 5469 6466 5747 6499
rect 5781 6499 6371 6500
rect 5781 6466 6059 6499
rect 5469 6465 6059 6466
rect 6093 6466 6371 6499
rect 6405 6499 6995 6500
rect 6405 6466 6683 6499
rect 6093 6465 6683 6466
rect 6717 6466 6995 6499
rect 7029 6499 7619 6500
rect 7029 6466 7307 6499
rect 6717 6465 7307 6466
rect 7341 6466 7619 6499
rect 7653 6499 8555 6500
rect 7653 6466 7931 6499
rect 7341 6465 7931 6466
rect 7965 6465 8243 6499
rect 8277 6466 8555 6499
rect 8589 6499 8941 6500
rect 8589 6466 8867 6499
rect 8277 6465 8867 6466
rect 8901 6465 8941 6499
rect 4033 6462 8941 6465
rect 8993 6462 9011 6514
rect 9063 6462 9064 6514
rect 4033 6450 9064 6462
rect 4033 6448 8941 6450
rect 1217 6430 8941 6448
rect 1217 6427 3857 6430
rect 1217 6393 1379 6427
rect 1413 6426 2003 6427
rect 1413 6393 1691 6426
rect 1217 6392 1691 6393
rect 1725 6393 2003 6426
rect 2037 6426 2627 6427
rect 2037 6393 2315 6426
rect 1725 6392 2315 6393
rect 2349 6393 2627 6426
rect 2661 6426 3857 6427
rect 2661 6393 2939 6426
rect 2349 6392 2939 6393
rect 2973 6392 3251 6426
rect 3285 6392 3563 6426
rect 3597 6392 3857 6426
rect 1217 6378 3857 6392
rect 3909 6378 3981 6430
rect 4033 6427 8941 6430
rect 4033 6426 4499 6427
rect 4033 6392 4187 6426
rect 4221 6393 4499 6426
rect 4533 6426 5123 6427
rect 4533 6393 4811 6426
rect 4221 6392 4811 6393
rect 4845 6393 5123 6426
rect 5157 6426 5747 6427
rect 5157 6393 5435 6426
rect 4845 6392 5435 6393
rect 5469 6393 5747 6426
rect 5781 6426 6371 6427
rect 5781 6393 6059 6426
rect 5469 6392 6059 6393
rect 6093 6393 6371 6426
rect 6405 6426 6995 6427
rect 6405 6393 6683 6426
rect 6093 6392 6683 6393
rect 6717 6393 6995 6426
rect 7029 6426 7619 6427
rect 7029 6393 7307 6426
rect 6717 6392 7307 6393
rect 7341 6393 7619 6426
rect 7653 6426 8555 6427
rect 7653 6393 7931 6426
rect 7341 6392 7931 6393
rect 7965 6392 8243 6426
rect 8277 6393 8555 6426
rect 8589 6426 8941 6427
rect 8589 6393 8867 6426
rect 8277 6392 8867 6393
rect 8901 6398 8941 6426
rect 8993 6398 9011 6450
rect 9063 6398 9064 6450
rect 8901 6392 9064 6398
rect 4033 6386 9064 6392
rect 4033 6378 8941 6386
rect 1217 6359 8941 6378
rect 1217 6354 3857 6359
rect 1217 6320 1379 6354
rect 1413 6353 2003 6354
rect 1413 6320 1691 6353
rect 1217 6319 1691 6320
rect 1725 6320 2003 6353
rect 2037 6353 2627 6354
rect 2037 6320 2315 6353
rect 1725 6319 2315 6320
rect 2349 6320 2627 6353
rect 2661 6353 3857 6354
rect 2661 6320 2939 6353
rect 2349 6319 2939 6320
rect 2973 6319 3251 6353
rect 3285 6319 3563 6353
rect 3597 6319 3857 6353
rect 1217 6307 3857 6319
rect 3909 6307 3981 6359
rect 4033 6354 8941 6359
rect 4033 6353 4499 6354
rect 4033 6319 4187 6353
rect 4221 6320 4499 6353
rect 4533 6353 5123 6354
rect 4533 6320 4811 6353
rect 4221 6319 4811 6320
rect 4845 6320 5123 6353
rect 5157 6353 5747 6354
rect 5157 6320 5435 6353
rect 4845 6319 5435 6320
rect 5469 6320 5747 6353
rect 5781 6353 6371 6354
rect 5781 6320 6059 6353
rect 5469 6319 6059 6320
rect 6093 6320 6371 6353
rect 6405 6353 6995 6354
rect 6405 6320 6683 6353
rect 6093 6319 6683 6320
rect 6717 6320 6995 6353
rect 7029 6353 7619 6354
rect 7029 6320 7307 6353
rect 6717 6319 7307 6320
rect 7341 6320 7619 6353
rect 7653 6353 8555 6354
rect 7653 6320 7931 6353
rect 7341 6319 7931 6320
rect 7965 6319 8243 6353
rect 8277 6320 8555 6353
rect 8589 6353 8941 6354
rect 8589 6320 8867 6353
rect 8277 6319 8867 6320
rect 8901 6334 8941 6353
rect 8993 6334 9011 6386
rect 9063 6334 9064 6386
rect 8901 6322 9064 6334
rect 8901 6319 8941 6322
rect 4033 6307 8941 6319
rect 1217 6288 8941 6307
rect 1217 6281 3857 6288
rect 1217 6247 1379 6281
rect 1413 6280 2003 6281
rect 1413 6247 1691 6280
rect 1217 6246 1691 6247
rect 1725 6247 2003 6280
rect 2037 6280 2627 6281
rect 2037 6247 2315 6280
rect 1725 6246 2315 6247
rect 2349 6247 2627 6280
rect 2661 6280 3857 6281
rect 2661 6247 2939 6280
rect 2349 6246 2939 6247
rect 2973 6246 3251 6280
rect 3285 6246 3563 6280
rect 3597 6246 3857 6280
rect 1217 6236 3857 6246
rect 3909 6236 3981 6288
rect 4033 6281 8941 6288
rect 4033 6280 4499 6281
rect 4033 6246 4187 6280
rect 4221 6247 4499 6280
rect 4533 6280 5123 6281
rect 4533 6247 4811 6280
rect 4221 6246 4811 6247
rect 4845 6247 5123 6280
rect 5157 6280 5747 6281
rect 5157 6247 5435 6280
rect 4845 6246 5435 6247
rect 5469 6247 5747 6280
rect 5781 6280 6371 6281
rect 5781 6247 6059 6280
rect 5469 6246 6059 6247
rect 6093 6247 6371 6280
rect 6405 6280 6995 6281
rect 6405 6247 6683 6280
rect 6093 6246 6683 6247
rect 6717 6247 6995 6280
rect 7029 6280 7619 6281
rect 7029 6247 7307 6280
rect 6717 6246 7307 6247
rect 7341 6247 7619 6280
rect 7653 6280 8555 6281
rect 7653 6247 7931 6280
rect 7341 6246 7931 6247
rect 7965 6246 8243 6280
rect 8277 6247 8555 6280
rect 8589 6280 8941 6281
rect 8589 6247 8867 6280
rect 8277 6246 8867 6247
rect 8901 6270 8941 6280
rect 8993 6270 9011 6322
rect 9063 6270 9064 6322
rect 8901 6258 9064 6270
rect 8901 6246 8941 6258
rect 4033 6236 8941 6246
rect 1217 6217 8941 6236
rect 1217 6208 3857 6217
rect 1217 6174 1379 6208
rect 1413 6207 2003 6208
rect 1413 6174 1691 6207
rect 1217 6173 1691 6174
rect 1725 6174 2003 6207
rect 2037 6207 2627 6208
rect 2037 6174 2315 6207
rect 1725 6173 2315 6174
rect 2349 6174 2627 6207
rect 2661 6207 3857 6208
rect 2661 6174 2939 6207
rect 2349 6173 2939 6174
rect 2973 6173 3251 6207
rect 3285 6173 3563 6207
rect 3597 6173 3857 6207
rect 1217 6165 3857 6173
rect 3909 6165 3981 6217
rect 4033 6208 8941 6217
rect 4033 6207 4499 6208
rect 4033 6173 4187 6207
rect 4221 6174 4499 6207
rect 4533 6207 5123 6208
rect 4533 6174 4811 6207
rect 4221 6173 4811 6174
rect 4845 6174 5123 6207
rect 5157 6207 5747 6208
rect 5157 6174 5435 6207
rect 4845 6173 5435 6174
rect 5469 6174 5747 6207
rect 5781 6207 6371 6208
rect 5781 6174 6059 6207
rect 5469 6173 6059 6174
rect 6093 6174 6371 6207
rect 6405 6207 6995 6208
rect 6405 6174 6683 6207
rect 6093 6173 6683 6174
rect 6717 6174 6995 6207
rect 7029 6207 7619 6208
rect 7029 6174 7307 6207
rect 6717 6173 7307 6174
rect 7341 6174 7619 6207
rect 7653 6207 8555 6208
rect 7653 6174 7931 6207
rect 7341 6173 7931 6174
rect 7965 6173 8243 6207
rect 8277 6174 8555 6207
rect 8589 6207 8941 6208
rect 8589 6174 8867 6207
rect 8277 6173 8867 6174
rect 8901 6206 8941 6207
rect 8993 6206 9011 6258
rect 9063 6206 9064 6258
rect 8901 6194 9064 6206
rect 8901 6173 8941 6194
rect 4033 6165 8941 6173
rect 1217 6146 8941 6165
rect 1217 6135 3857 6146
rect 1217 6101 1379 6135
rect 1413 6134 2003 6135
rect 1413 6101 1691 6134
rect 1217 6100 1691 6101
rect 1725 6101 2003 6134
rect 2037 6134 2627 6135
rect 2037 6101 2315 6134
rect 1725 6100 2315 6101
rect 2349 6101 2627 6134
rect 2661 6134 3857 6135
rect 2661 6101 2939 6134
rect 2349 6100 2939 6101
rect 2973 6100 3251 6134
rect 3285 6100 3563 6134
rect 3597 6100 3857 6134
rect 1217 6094 3857 6100
rect 3909 6094 3981 6146
rect 4033 6142 8941 6146
rect 8993 6142 9011 6194
rect 9063 6142 9064 6194
rect 4033 6135 9064 6142
rect 4033 6134 4499 6135
rect 4033 6100 4187 6134
rect 4221 6101 4499 6134
rect 4533 6134 5123 6135
rect 4533 6101 4811 6134
rect 4221 6100 4811 6101
rect 4845 6101 5123 6134
rect 5157 6134 5747 6135
rect 5157 6101 5435 6134
rect 4845 6100 5435 6101
rect 5469 6101 5747 6134
rect 5781 6134 6371 6135
rect 5781 6101 6059 6134
rect 5469 6100 6059 6101
rect 6093 6101 6371 6134
rect 6405 6134 6995 6135
rect 6405 6101 6683 6134
rect 6093 6100 6683 6101
rect 6717 6101 6995 6134
rect 7029 6134 7619 6135
rect 7029 6101 7307 6134
rect 6717 6100 7307 6101
rect 7341 6101 7619 6134
rect 7653 6134 8555 6135
rect 7653 6101 7931 6134
rect 7341 6100 7931 6101
rect 7965 6100 8243 6134
rect 8277 6101 8555 6134
rect 8589 6134 9064 6135
rect 8589 6101 8867 6134
rect 8277 6100 8867 6101
rect 8901 6130 9064 6134
rect 8901 6100 8941 6130
rect 4033 6094 8941 6100
rect 1217 6078 8941 6094
rect 8993 6078 9011 6130
rect 9063 6078 9064 6130
rect 1217 6075 9064 6078
rect 1217 6062 3857 6075
rect 1217 6028 1379 6062
rect 1413 6061 2003 6062
rect 1413 6028 1691 6061
rect 1217 6027 1691 6028
rect 1725 6028 2003 6061
rect 2037 6061 2627 6062
rect 2037 6028 2315 6061
rect 1725 6027 2315 6028
rect 2349 6028 2627 6061
rect 2661 6061 3857 6062
rect 2661 6028 2939 6061
rect 2349 6027 2939 6028
rect 2973 6027 3251 6061
rect 3285 6027 3563 6061
rect 3597 6027 3857 6061
rect 1217 6023 3857 6027
rect 3909 6023 3981 6075
rect 4033 6065 9064 6075
rect 4033 6062 8941 6065
rect 4033 6061 4499 6062
rect 4033 6027 4187 6061
rect 4221 6028 4499 6061
rect 4533 6061 5123 6062
rect 4533 6028 4811 6061
rect 4221 6027 4811 6028
rect 4845 6028 5123 6061
rect 5157 6061 5747 6062
rect 5157 6028 5435 6061
rect 4845 6027 5435 6028
rect 5469 6028 5747 6061
rect 5781 6061 6371 6062
rect 5781 6028 6059 6061
rect 5469 6027 6059 6028
rect 6093 6028 6371 6061
rect 6405 6061 6995 6062
rect 6405 6028 6683 6061
rect 6093 6027 6683 6028
rect 6717 6028 6995 6061
rect 7029 6061 7619 6062
rect 7029 6028 7307 6061
rect 6717 6027 7307 6028
rect 7341 6028 7619 6061
rect 7653 6061 8555 6062
rect 7653 6028 7931 6061
rect 7341 6027 7931 6028
rect 7965 6027 8243 6061
rect 8277 6028 8555 6061
rect 8589 6061 8941 6062
rect 8589 6028 8867 6061
rect 8277 6027 8867 6028
rect 8901 6027 8941 6061
rect 4033 6023 8941 6027
rect 1217 6013 8941 6023
rect 8993 6013 9011 6065
rect 9063 6013 9064 6065
rect 1217 6004 9064 6013
rect 1217 5989 3857 6004
rect 1217 5955 1379 5989
rect 1413 5988 2003 5989
rect 1413 5955 1691 5988
rect 1217 5954 1691 5955
rect 1725 5955 2003 5988
rect 2037 5988 2627 5989
rect 2037 5955 2315 5988
rect 1725 5954 2315 5955
rect 2349 5955 2627 5988
rect 2661 5988 3857 5989
rect 2661 5955 2939 5988
rect 2349 5954 2939 5955
rect 2973 5954 3251 5988
rect 3285 5954 3563 5988
rect 3597 5954 3857 5988
rect 1217 5952 3857 5954
rect 3909 5952 3981 6004
rect 4033 6000 9064 6004
rect 4033 5989 8941 6000
rect 4033 5988 4499 5989
rect 4033 5954 4187 5988
rect 4221 5955 4499 5988
rect 4533 5988 5123 5989
rect 4533 5955 4811 5988
rect 4221 5954 4811 5955
rect 4845 5955 5123 5988
rect 5157 5988 5747 5989
rect 5157 5955 5435 5988
rect 4845 5954 5435 5955
rect 5469 5955 5747 5988
rect 5781 5988 6371 5989
rect 5781 5955 6059 5988
rect 5469 5954 6059 5955
rect 6093 5955 6371 5988
rect 6405 5988 6995 5989
rect 6405 5955 6683 5988
rect 6093 5954 6683 5955
rect 6717 5955 6995 5988
rect 7029 5988 7619 5989
rect 7029 5955 7307 5988
rect 6717 5954 7307 5955
rect 7341 5955 7619 5988
rect 7653 5988 8555 5989
rect 7653 5955 7931 5988
rect 7341 5954 7931 5955
rect 7965 5954 8243 5988
rect 8277 5955 8555 5988
rect 8589 5988 8941 5989
rect 8589 5955 8867 5988
rect 8277 5954 8867 5955
rect 8901 5954 8941 5988
rect 4033 5952 8941 5954
rect 1217 5948 8941 5952
rect 8993 5948 9011 6000
rect 9063 5948 9064 6000
rect 1217 5942 9064 5948
rect 9151 6551 9197 6592
rect 9151 6517 9157 6551
rect 9191 6517 9197 6551
rect 9151 6476 9197 6517
rect 9151 6442 9157 6476
rect 9191 6442 9197 6476
rect 9151 6401 9197 6442
rect 9151 6367 9157 6401
rect 9191 6367 9197 6401
rect 9151 6326 9197 6367
rect 9151 6292 9157 6326
rect 9191 6292 9197 6326
rect 9151 6251 9197 6292
rect 9151 6217 9157 6251
rect 9191 6217 9197 6251
rect 9151 6176 9197 6217
rect 9151 6142 9157 6176
rect 9191 6142 9197 6176
rect 9151 6101 9197 6142
rect 9151 6067 9157 6101
rect 9191 6067 9197 6101
rect 9151 6026 9197 6067
rect 9151 5992 9157 6026
rect 9191 5992 9197 6026
rect 9151 5951 9197 5992
tri 9145 5920 9151 5926 se
rect 9151 5920 9157 5951
rect 941 5917 987 5920
tri 987 5917 990 5920 sw
tri 9142 5917 9145 5920 se
rect 9145 5917 9157 5920
rect 9191 5917 9197 5951
rect 941 5905 990 5917
tri 990 5905 1002 5917 sw
tri 9130 5905 9142 5917 se
rect 9142 5905 9197 5917
rect 941 5886 1002 5905
tri 1002 5886 1021 5905 sw
tri 9111 5886 9130 5905 se
rect 9130 5886 9197 5905
rect 941 5880 9197 5886
rect 941 5846 1019 5880
rect 1053 5846 1092 5880
rect 1126 5846 1165 5880
rect 1199 5846 1237 5880
rect 1271 5846 1309 5880
rect 1343 5846 1381 5880
rect 1415 5846 1453 5880
rect 1487 5846 1525 5880
rect 1559 5846 1597 5880
rect 1631 5846 1669 5880
rect 1703 5846 1741 5880
rect 1775 5846 1813 5880
rect 1847 5846 1885 5880
rect 1919 5846 1957 5880
rect 1991 5846 2029 5880
rect 2063 5846 2101 5880
rect 2135 5846 2173 5880
rect 2207 5846 2245 5880
rect 2279 5846 2317 5880
rect 2351 5846 2389 5880
rect 2423 5846 2461 5880
rect 2495 5846 2533 5880
rect 2567 5846 2605 5880
rect 2639 5846 2677 5880
rect 2711 5846 2749 5880
rect 2783 5846 2821 5880
rect 2855 5846 2893 5880
rect 2927 5846 2965 5880
rect 2999 5846 3037 5880
rect 3071 5846 3109 5880
rect 3143 5846 3181 5880
rect 3215 5846 3253 5880
rect 3287 5846 3325 5880
rect 3359 5846 3397 5880
rect 3431 5846 3469 5880
rect 3503 5846 3541 5880
rect 3575 5846 3613 5880
rect 3647 5846 3685 5880
rect 3719 5846 3757 5880
rect 3791 5846 3829 5880
rect 3863 5846 3901 5880
rect 3935 5846 3973 5880
rect 4007 5846 4045 5880
rect 4079 5846 4117 5880
rect 4151 5846 4189 5880
rect 4223 5846 4261 5880
rect 4295 5846 4333 5880
rect 4367 5846 4405 5880
rect 4439 5846 4477 5880
rect 4511 5846 4549 5880
rect 4583 5846 4621 5880
rect 4655 5846 4693 5880
rect 4727 5846 4765 5880
rect 4799 5846 4837 5880
rect 4871 5846 4909 5880
rect 4943 5846 4981 5880
rect 5015 5846 5053 5880
rect 5087 5846 5125 5880
rect 5159 5846 5197 5880
rect 5231 5846 5269 5880
rect 5303 5846 5341 5880
rect 5375 5846 5413 5880
rect 5447 5846 5485 5880
rect 5519 5846 5557 5880
rect 5591 5846 5629 5880
rect 5663 5846 5701 5880
rect 5735 5846 5773 5880
rect 5807 5846 5845 5880
rect 5879 5846 5917 5880
rect 5951 5846 5989 5880
rect 6023 5846 6061 5880
rect 6095 5846 6133 5880
rect 6167 5846 6205 5880
rect 6239 5846 6277 5880
rect 6311 5846 6349 5880
rect 6383 5846 6421 5880
rect 6455 5846 6493 5880
rect 6527 5846 6565 5880
rect 6599 5846 6637 5880
rect 6671 5846 6709 5880
rect 6743 5846 6781 5880
rect 6815 5846 6853 5880
rect 6887 5846 6925 5880
rect 6959 5846 6997 5880
rect 7031 5846 7069 5880
rect 7103 5846 7141 5880
rect 7175 5846 7213 5880
rect 7247 5846 7285 5880
rect 7319 5846 7357 5880
rect 7391 5846 7429 5880
rect 7463 5846 7501 5880
rect 7535 5846 7573 5880
rect 7607 5846 7645 5880
rect 7679 5846 7717 5880
rect 7751 5846 7789 5880
rect 7823 5846 7861 5880
rect 7895 5846 7933 5880
rect 7967 5846 8005 5880
rect 8039 5846 8077 5880
rect 8111 5846 8149 5880
rect 8183 5846 8221 5880
rect 8255 5846 8293 5880
rect 8327 5846 8365 5880
rect 8399 5846 8437 5880
rect 8471 5846 8509 5880
rect 8543 5846 8581 5880
rect 8615 5846 8653 5880
rect 8687 5846 8725 5880
rect 8759 5846 8797 5880
rect 8831 5846 8869 5880
rect 8903 5846 8941 5880
rect 8975 5846 9013 5880
rect 9047 5846 9085 5880
rect 9119 5846 9197 5880
rect 941 5840 9197 5846
rect 9456 7517 9462 7551
rect 9496 7549 9646 7551
rect 9496 7517 9534 7549
rect 9456 7515 9534 7517
rect 9568 7515 9606 7549
rect 9640 7515 9646 7549
rect 9456 7477 9646 7515
rect 9456 7443 9462 7477
rect 9496 7475 9646 7477
rect 9496 7443 9534 7475
rect 9456 7441 9534 7443
rect 9568 7441 9606 7475
rect 9640 7441 9646 7475
rect 9456 7403 9646 7441
rect 9456 7369 9462 7403
rect 9496 7401 9646 7403
rect 9496 7369 9534 7401
rect 9456 7367 9534 7369
rect 9568 7367 9606 7401
rect 9640 7367 9646 7401
rect 9456 7329 9646 7367
rect 9456 7295 9462 7329
rect 9496 7327 9646 7329
rect 9496 7295 9534 7327
rect 9456 7293 9534 7295
rect 9568 7293 9606 7327
rect 9640 7293 9646 7327
rect 9456 7255 9646 7293
rect 9456 7221 9462 7255
rect 9496 7253 9646 7255
rect 9496 7221 9534 7253
rect 9456 7219 9534 7221
rect 9568 7219 9606 7253
rect 9640 7219 9646 7253
rect 9456 7181 9646 7219
rect 9456 7147 9462 7181
rect 9496 7180 9646 7181
rect 9496 7147 9534 7180
rect 9456 7146 9534 7147
rect 9568 7146 9606 7180
rect 9640 7146 9646 7180
rect 9456 7107 9646 7146
rect 9456 7073 9462 7107
rect 9496 7073 9534 7107
rect 9568 7073 9606 7107
rect 9640 7073 9646 7107
rect 9456 7034 9646 7073
rect 9456 7000 9462 7034
rect 9496 7000 9534 7034
rect 9568 7000 9606 7034
rect 9640 7000 9646 7034
rect 9456 6961 9646 7000
rect 9456 6927 9462 6961
rect 9496 6927 9534 6961
rect 9568 6927 9606 6961
rect 9640 6927 9646 6961
rect 9456 6888 9646 6927
rect 9456 6854 9462 6888
rect 9496 6854 9534 6888
rect 9568 6854 9606 6888
rect 9640 6854 9646 6888
rect 9456 6815 9646 6854
rect 9456 6781 9462 6815
rect 9496 6781 9534 6815
rect 9568 6781 9606 6815
rect 9640 6781 9646 6815
rect 9456 6742 9646 6781
rect 9456 6708 9462 6742
rect 9496 6708 9534 6742
rect 9568 6708 9606 6742
rect 9640 6708 9646 6742
rect 9456 6669 9646 6708
rect 9456 6635 9462 6669
rect 9496 6635 9534 6669
rect 9568 6635 9606 6669
rect 9640 6635 9646 6669
rect 9456 6596 9646 6635
rect 9456 6562 9462 6596
rect 9496 6562 9534 6596
rect 9568 6562 9606 6596
rect 9640 6562 9646 6596
rect 9456 6523 9646 6562
rect 9456 6489 9462 6523
rect 9496 6489 9534 6523
rect 9568 6489 9606 6523
rect 9640 6489 9646 6523
rect 9456 6450 9646 6489
rect 9456 6416 9462 6450
rect 9496 6416 9534 6450
rect 9568 6416 9606 6450
rect 9640 6416 9646 6450
rect 9456 6377 9646 6416
rect 9456 6343 9462 6377
rect 9496 6343 9534 6377
rect 9568 6343 9606 6377
rect 9640 6343 9646 6377
rect 9456 6304 9646 6343
rect 9456 6270 9462 6304
rect 9496 6270 9534 6304
rect 9568 6270 9606 6304
rect 9640 6270 9646 6304
rect 9456 6231 9646 6270
rect 9456 6197 9462 6231
rect 9496 6197 9534 6231
rect 9568 6197 9606 6231
rect 9640 6197 9646 6231
rect 9456 6158 9646 6197
rect 9456 6124 9462 6158
rect 9496 6124 9534 6158
rect 9568 6124 9606 6158
rect 9640 6124 9646 6158
rect 9456 6085 9646 6124
rect 9456 6051 9462 6085
rect 9496 6051 9534 6085
rect 9568 6051 9606 6085
rect 9640 6051 9646 6085
rect 9456 6012 9646 6051
rect 9456 5978 9462 6012
rect 9496 5978 9534 6012
rect 9568 5978 9606 6012
rect 9640 5978 9646 6012
rect 9456 5939 9646 5978
rect 9456 5905 9462 5939
rect 9496 5905 9534 5939
rect 9568 5905 9606 5939
rect 9640 5905 9646 5939
rect 9456 5843 9646 5905
rect 732 5792 770 5801
rect 620 5753 631 5792
rect 683 5791 770 5792
rect 804 5791 810 5825
rect 683 5788 810 5791
rect 683 5753 749 5788
rect 620 5719 626 5753
rect 683 5747 698 5753
rect 660 5734 698 5747
rect 683 5719 698 5734
rect 732 5736 749 5753
rect 801 5752 810 5788
rect 732 5723 770 5736
rect 732 5719 749 5723
rect 620 5682 631 5719
rect 683 5682 749 5719
rect 804 5718 810 5752
rect 620 5680 749 5682
rect 620 5646 626 5680
rect 660 5669 698 5680
rect 683 5646 698 5669
rect 732 5671 749 5680
rect 801 5679 810 5718
rect 732 5658 770 5671
rect 732 5646 749 5658
rect 620 5617 631 5646
rect 683 5617 749 5646
rect 804 5651 810 5679
rect 9456 5809 9462 5843
rect 9496 5809 9534 5843
rect 9568 5809 9606 5843
rect 9640 5809 9646 5843
rect 9456 5766 9646 5809
rect 10458 7917 10648 7954
rect 10458 7915 10608 7917
rect 10458 7881 10464 7915
rect 10498 7881 10536 7915
rect 10570 7883 10608 7915
rect 10642 7883 10648 7917
rect 10570 7881 10648 7883
rect 10458 7844 10648 7881
rect 10458 7842 10608 7844
rect 10458 7808 10464 7842
rect 10498 7808 10536 7842
rect 10570 7810 10608 7842
rect 10642 7810 10648 7844
rect 10570 7808 10648 7810
rect 10458 7771 10648 7808
rect 10458 7769 10608 7771
rect 10458 7735 10464 7769
rect 10498 7735 10536 7769
rect 10570 7737 10608 7769
rect 10642 7737 10648 7771
rect 10683 8162 14724 8210
rect 10683 8007 10731 8162
tri 10731 8128 10765 8162 nw
tri 14642 8128 14676 8162 ne
rect 10786 8116 13427 8122
rect 10786 8082 10864 8116
rect 10898 8082 10936 8116
rect 10970 8082 11008 8116
rect 11042 8082 11080 8116
rect 11114 8082 11152 8116
rect 11186 8082 11224 8116
rect 11258 8082 11296 8116
rect 11330 8082 11368 8116
rect 11402 8082 11440 8116
rect 11474 8082 11512 8116
rect 11546 8082 11584 8116
rect 11618 8082 11656 8116
rect 11690 8082 11728 8116
rect 11762 8082 11800 8116
rect 11834 8082 11872 8116
rect 11906 8082 11944 8116
rect 11978 8082 12016 8116
rect 12050 8082 12088 8116
rect 12122 8082 12160 8116
rect 12194 8082 12232 8116
rect 12266 8082 12304 8116
rect 12338 8082 12376 8116
rect 12410 8082 12448 8116
rect 12482 8082 12520 8116
rect 12554 8082 12592 8116
rect 12626 8082 12664 8116
rect 12698 8082 12736 8116
rect 12770 8082 12808 8116
rect 12842 8082 12880 8116
rect 12914 8082 12952 8116
rect 12986 8082 13024 8116
rect 13058 8082 13096 8116
rect 13130 8082 13169 8116
rect 13203 8082 13242 8116
rect 13276 8082 13315 8116
rect 13349 8082 13427 8116
rect 10786 8076 13427 8082
rect 10786 8062 10845 8076
tri 10845 8062 10859 8076 nw
tri 13329 8062 13343 8076 ne
rect 13343 8062 13427 8076
rect 10786 8049 10832 8062
tri 10832 8049 10845 8062 nw
tri 13343 8049 13356 8062 ne
rect 13356 8049 13427 8062
tri 13356 8041 13364 8049 ne
rect 13364 8041 13427 8049
tri 13364 8028 13377 8041 ne
rect 13377 8028 13387 8041
tri 10731 8007 10752 8028 sw
tri 13377 8024 13381 8028 ne
rect 13381 8007 13387 8028
rect 13421 8007 13427 8041
rect 10683 7994 10752 8007
tri 10752 7994 10765 8007 sw
rect 10683 7988 13267 7994
rect 10683 7954 10995 7988
rect 11029 7954 11070 7988
rect 11104 7954 11145 7988
rect 11179 7954 11220 7988
rect 11254 7954 11295 7988
rect 11329 7954 11370 7988
rect 11404 7954 11445 7988
rect 11479 7954 11519 7988
rect 11553 7954 11593 7988
rect 11627 7954 11667 7988
rect 11701 7954 11741 7988
rect 11775 7954 11815 7988
rect 11849 7954 11889 7988
rect 11923 7954 11963 7988
rect 11997 7954 12037 7988
rect 12071 7954 12111 7988
rect 12145 7954 12185 7988
rect 12219 7954 12259 7988
rect 12293 7954 12333 7988
rect 12367 7954 12407 7988
rect 12441 7954 12481 7988
rect 12515 7954 12555 7988
rect 12589 7954 12629 7988
rect 12663 7954 12703 7988
rect 12737 7954 12777 7988
rect 12811 7954 12851 7988
rect 12885 7954 12925 7988
rect 12959 7954 12999 7988
rect 13033 7954 13073 7988
rect 13107 7954 13147 7988
rect 13181 7954 13221 7988
rect 13255 7954 13267 7988
rect 10683 7948 13267 7954
rect 13381 7966 13427 8007
rect 10683 7932 10747 7948
tri 10747 7932 10763 7948 nw
rect 13381 7932 13387 7966
rect 13421 7932 13427 7966
rect 10570 7735 10648 7737
rect 10458 7698 10648 7735
rect 10458 7696 10608 7698
rect 10458 7662 10464 7696
rect 10498 7662 10536 7696
rect 10570 7664 10608 7696
rect 10642 7664 10648 7698
rect 10570 7662 10648 7664
rect 10458 7625 10648 7662
tri 10677 7756 10683 7762 se
rect 10683 7756 10729 7932
tri 10729 7914 10747 7932 nw
tri 13367 7914 13381 7928 se
rect 13381 7914 13427 7932
tri 13344 7891 13367 7914 se
rect 13367 7891 13427 7914
tri 13323 7870 13344 7891 se
rect 13344 7870 13387 7891
rect 10677 7750 10729 7756
rect 10677 7686 10729 7698
rect 10677 7628 10729 7634
rect 10786 7864 13387 7870
rect 10786 7858 10934 7864
rect 10786 7824 10792 7858
rect 10826 7824 10934 7858
rect 10786 7812 10934 7824
rect 10986 7812 11000 7864
rect 11052 7812 11066 7864
rect 11118 7812 11132 7864
rect 11184 7812 11198 7864
rect 11250 7858 11264 7864
rect 11250 7824 11251 7858
rect 11250 7812 11264 7824
rect 11316 7812 11330 7864
rect 11382 7858 13387 7864
rect 11382 7824 11563 7858
rect 11597 7824 11875 7858
rect 11909 7824 12187 7858
rect 12221 7824 12499 7858
rect 12533 7824 12811 7858
rect 12845 7824 13123 7858
rect 13157 7857 13387 7858
rect 13421 7857 13427 7891
rect 13157 7824 13427 7857
rect 11382 7816 13427 7824
rect 11382 7812 13387 7816
rect 10786 7793 13387 7812
rect 10786 7784 10934 7793
rect 10786 7750 10792 7784
rect 10826 7750 10934 7784
rect 10786 7741 10934 7750
rect 10986 7741 11000 7793
rect 11052 7741 11066 7793
rect 11118 7741 11132 7793
rect 11184 7741 11198 7793
rect 11250 7785 11264 7793
rect 11250 7751 11251 7785
rect 11250 7741 11264 7751
rect 11316 7741 11330 7793
rect 11382 7785 13387 7793
rect 11382 7751 11563 7785
rect 11597 7751 11875 7785
rect 11909 7751 12187 7785
rect 12221 7751 12499 7785
rect 12533 7751 12811 7785
rect 12845 7751 13123 7785
rect 13157 7782 13387 7785
rect 13421 7782 13427 7816
rect 13157 7751 13427 7782
rect 11382 7741 13427 7751
rect 10786 7722 13387 7741
rect 10786 7710 10934 7722
rect 10786 7676 10792 7710
rect 10826 7676 10934 7710
rect 10786 7670 10934 7676
rect 10986 7670 11000 7722
rect 11052 7670 11066 7722
rect 11118 7670 11132 7722
rect 11184 7670 11198 7722
rect 11250 7712 11264 7722
rect 11250 7678 11251 7712
rect 11250 7670 11264 7678
rect 11316 7670 11330 7722
rect 11382 7712 13387 7722
rect 11382 7678 11563 7712
rect 11597 7678 11875 7712
rect 11909 7678 12187 7712
rect 12221 7678 12499 7712
rect 12533 7678 12811 7712
rect 12845 7678 13123 7712
rect 13157 7707 13387 7712
rect 13421 7707 13427 7741
rect 13157 7678 13427 7707
rect 11382 7670 13427 7678
rect 10786 7666 13427 7670
rect 10786 7651 13387 7666
rect 10786 7636 10934 7651
rect 10458 7623 10608 7625
rect 10458 7589 10464 7623
rect 10498 7589 10536 7623
rect 10570 7591 10608 7623
rect 10642 7591 10648 7625
rect 10570 7589 10648 7591
rect 10458 7552 10648 7589
rect 10458 7550 10608 7552
rect 10458 7516 10464 7550
rect 10498 7516 10536 7550
rect 10570 7518 10608 7550
rect 10642 7518 10648 7552
rect 10570 7516 10648 7518
rect 10458 7479 10648 7516
rect 10458 7477 10608 7479
rect 10458 7443 10464 7477
rect 10498 7443 10536 7477
rect 10570 7445 10608 7477
rect 10642 7445 10648 7479
rect 10570 7443 10648 7445
rect 10458 7406 10648 7443
rect 10458 7404 10608 7406
rect 10458 7370 10464 7404
rect 10498 7370 10536 7404
rect 10570 7372 10608 7404
rect 10642 7372 10648 7406
rect 10570 7370 10648 7372
rect 10458 7333 10648 7370
rect 10458 7331 10608 7333
rect 10458 7297 10464 7331
rect 10498 7297 10536 7331
rect 10570 7299 10608 7331
rect 10642 7299 10648 7333
rect 10570 7297 10648 7299
rect 10458 7260 10648 7297
rect 10458 7258 10608 7260
rect 10458 7224 10464 7258
rect 10498 7224 10536 7258
rect 10570 7226 10608 7258
rect 10642 7226 10648 7260
rect 10570 7224 10648 7226
rect 10786 7602 10792 7636
rect 10826 7602 10934 7636
rect 10786 7599 10934 7602
rect 10986 7599 11000 7651
rect 11052 7599 11066 7651
rect 11118 7599 11132 7651
rect 11184 7599 11198 7651
rect 11250 7639 11264 7651
rect 11250 7605 11251 7639
rect 11250 7599 11264 7605
rect 11316 7599 11330 7651
rect 11382 7639 13387 7651
rect 11382 7605 11563 7639
rect 11597 7605 11875 7639
rect 11909 7605 12187 7639
rect 12221 7605 12499 7639
rect 12533 7605 12811 7639
rect 12845 7605 13123 7639
rect 13157 7632 13387 7639
rect 13421 7632 13427 7666
rect 13157 7605 13427 7632
rect 11382 7599 13427 7605
rect 10786 7591 13427 7599
rect 10786 7579 13387 7591
rect 10786 7563 10934 7579
rect 10786 7529 10792 7563
rect 10826 7529 10934 7563
rect 10786 7527 10934 7529
rect 10986 7527 11000 7579
rect 11052 7527 11066 7579
rect 11118 7527 11132 7579
rect 11184 7527 11198 7579
rect 11250 7566 11264 7579
rect 11250 7532 11251 7566
rect 11250 7527 11264 7532
rect 11316 7527 11330 7579
rect 11382 7566 13387 7579
rect 11382 7532 11563 7566
rect 11597 7532 11875 7566
rect 11909 7532 12187 7566
rect 12221 7532 12499 7566
rect 12533 7532 12811 7566
rect 12845 7532 13123 7566
rect 13157 7557 13387 7566
rect 13421 7557 13427 7591
rect 13157 7532 13427 7557
rect 11382 7527 13427 7532
rect 10786 7516 13427 7527
rect 10786 7507 13387 7516
rect 10786 7490 10934 7507
rect 10786 7456 10792 7490
rect 10826 7456 10934 7490
rect 10786 7455 10934 7456
rect 10986 7455 11000 7507
rect 11052 7455 11066 7507
rect 11118 7455 11132 7507
rect 11184 7455 11198 7507
rect 11250 7493 11264 7507
rect 11250 7459 11251 7493
rect 11250 7455 11264 7459
rect 11316 7455 11330 7507
rect 11382 7493 13387 7507
rect 11382 7459 11563 7493
rect 11597 7459 11875 7493
rect 11909 7459 12187 7493
rect 12221 7459 12499 7493
rect 12533 7459 12811 7493
rect 12845 7459 13123 7493
rect 13157 7482 13387 7493
rect 13421 7482 13427 7516
rect 13157 7459 13427 7482
rect 11382 7455 13427 7459
rect 10786 7441 13427 7455
rect 10786 7435 13387 7441
rect 10786 7417 10934 7435
rect 10786 7383 10792 7417
rect 10826 7383 10934 7417
rect 10986 7383 11000 7435
rect 11052 7383 11066 7435
rect 11118 7383 11132 7435
rect 11184 7383 11198 7435
rect 11250 7420 11264 7435
rect 11250 7386 11251 7420
rect 11250 7383 11264 7386
rect 11316 7383 11330 7435
rect 11382 7420 13387 7435
rect 11382 7386 11563 7420
rect 11597 7386 11875 7420
rect 11909 7386 12187 7420
rect 12221 7386 12499 7420
rect 12533 7386 12811 7420
rect 12845 7386 13123 7420
rect 13157 7407 13387 7420
rect 13421 7407 13427 7441
rect 13157 7386 13427 7407
rect 11382 7383 13427 7386
rect 10786 7365 13427 7383
rect 10786 7363 13387 7365
rect 10786 7344 10934 7363
rect 10786 7310 10792 7344
rect 10826 7311 10934 7344
rect 10986 7311 11000 7363
rect 11052 7311 11066 7363
rect 11118 7311 11132 7363
rect 11184 7311 11198 7363
rect 11250 7346 11264 7363
rect 11250 7312 11251 7346
rect 11250 7311 11264 7312
rect 11316 7311 11330 7363
rect 11382 7346 13387 7363
rect 11382 7312 11563 7346
rect 11597 7312 11875 7346
rect 11909 7312 12187 7346
rect 12221 7312 12499 7346
rect 12533 7312 12811 7346
rect 12845 7312 13123 7346
rect 13157 7331 13387 7346
rect 13421 7331 13427 7365
rect 13157 7312 13427 7331
rect 11382 7311 13427 7312
rect 10826 7310 13427 7311
rect 10786 7291 13427 7310
rect 10786 7271 10934 7291
rect 10786 7237 10792 7271
rect 10826 7239 10934 7271
rect 10986 7239 11000 7291
rect 11052 7239 11066 7291
rect 11118 7239 11132 7291
rect 11184 7239 11198 7291
rect 11250 7272 11264 7291
rect 11250 7239 11251 7272
rect 11316 7239 11330 7291
rect 11382 7289 13427 7291
rect 11382 7272 13387 7289
rect 11382 7239 11563 7272
rect 10826 7238 10939 7239
rect 10973 7238 11251 7239
rect 11285 7238 11563 7239
rect 11597 7238 11875 7272
rect 11909 7238 12187 7272
rect 12221 7238 12499 7272
rect 12533 7238 12811 7272
rect 12845 7238 13123 7272
rect 13157 7255 13387 7272
rect 13421 7255 13427 7289
rect 13157 7238 13427 7255
rect 10826 7237 13427 7238
rect 10786 7225 13427 7237
rect 10458 7187 10648 7224
tri 13338 7213 13350 7225 ne
rect 13350 7213 13427 7225
rect 10458 7185 10608 7187
rect 10458 7151 10464 7185
rect 10498 7151 10536 7185
rect 10570 7153 10608 7185
rect 10642 7153 10648 7187
tri 13350 7182 13381 7213 ne
rect 13381 7179 13387 7213
rect 13421 7179 13427 7213
rect 10570 7151 10648 7153
rect 10458 7113 10648 7151
rect 10458 7112 10608 7113
rect 10458 7078 10464 7112
rect 10498 7078 10536 7112
rect 10570 7079 10608 7112
rect 10642 7079 10648 7113
rect 10570 7078 10648 7079
rect 10458 7039 10648 7078
rect 10458 7005 10464 7039
rect 10498 7005 10536 7039
rect 10570 7005 10608 7039
rect 10642 7005 10648 7039
rect 10458 6965 10648 7005
rect 10458 6931 10464 6965
rect 10498 6931 10536 6965
rect 10570 6931 10608 6965
rect 10642 6931 10648 6965
rect 10458 6891 10648 6931
rect 10458 6857 10464 6891
rect 10498 6857 10536 6891
rect 10570 6857 10608 6891
rect 10642 6857 10648 6891
rect 10458 6817 10648 6857
rect 10458 6783 10464 6817
rect 10498 6783 10536 6817
rect 10570 6783 10608 6817
rect 10642 6783 10648 6817
rect 10458 6743 10648 6783
rect 10458 6709 10464 6743
rect 10498 6709 10536 6743
rect 10570 6709 10608 6743
rect 10642 6709 10648 6743
rect 10458 6669 10648 6709
rect 10458 6635 10464 6669
rect 10498 6635 10536 6669
rect 10570 6635 10608 6669
rect 10642 6635 10648 6669
rect 10458 6595 10648 6635
rect 10458 6561 10464 6595
rect 10498 6561 10536 6595
rect 10570 6561 10608 6595
rect 10642 6561 10648 6595
rect 10458 6521 10648 6561
rect 10458 6487 10464 6521
rect 10498 6487 10536 6521
rect 10570 6487 10608 6521
rect 10642 6487 10648 6521
rect 10985 7160 13317 7166
rect 11037 7154 11111 7160
rect 11163 7154 13317 7160
rect 11037 7120 11093 7154
rect 11163 7120 11405 7154
rect 11439 7120 11717 7154
rect 11751 7120 12029 7154
rect 12063 7120 12341 7154
rect 12375 7120 12653 7154
rect 12687 7120 12965 7154
rect 12999 7120 13277 7154
rect 13311 7120 13317 7154
rect 11037 7108 11111 7120
rect 11163 7108 13317 7120
rect 10985 7095 13317 7108
rect 11037 7080 11111 7095
rect 11163 7080 13317 7095
rect 11037 7046 11093 7080
rect 11163 7046 11405 7080
rect 11439 7046 11717 7080
rect 11751 7046 12029 7080
rect 12063 7046 12341 7080
rect 12375 7046 12653 7080
rect 12687 7046 12965 7080
rect 12999 7046 13277 7080
rect 13311 7046 13317 7080
rect 11037 7043 11111 7046
rect 11163 7043 13317 7046
rect 10985 7030 13317 7043
rect 11037 7006 11111 7030
rect 11163 7006 13317 7030
rect 11037 6978 11093 7006
rect 11163 6978 11405 7006
rect 10985 6972 11093 6978
rect 11127 6972 11405 6978
rect 11439 6972 11717 7006
rect 11751 6972 12029 7006
rect 12063 6972 12341 7006
rect 12375 6972 12653 7006
rect 12687 6972 12965 7006
rect 12999 6972 13277 7006
rect 13311 6972 13317 7006
rect 10985 6965 13317 6972
rect 11037 6932 11111 6965
rect 11163 6932 13317 6965
rect 11037 6913 11093 6932
rect 11163 6913 11405 6932
rect 10985 6899 11093 6913
rect 11127 6899 11405 6913
rect 11037 6898 11093 6899
rect 11163 6898 11405 6899
rect 11439 6898 11717 6932
rect 11751 6898 12029 6932
rect 12063 6898 12341 6932
rect 12375 6898 12653 6932
rect 12687 6898 12965 6932
rect 12999 6898 13277 6932
rect 13311 6898 13317 6932
rect 11037 6858 11111 6898
rect 11163 6858 13317 6898
rect 11037 6847 11093 6858
rect 11163 6847 11405 6858
rect 10985 6833 11093 6847
rect 11127 6833 11405 6847
rect 11037 6824 11093 6833
rect 11163 6824 11405 6833
rect 11439 6824 11717 6858
rect 11751 6824 12029 6858
rect 12063 6824 12341 6858
rect 12375 6824 12653 6858
rect 12687 6824 12965 6858
rect 12999 6824 13277 6858
rect 13311 6824 13317 6858
rect 11037 6783 11111 6824
rect 11163 6783 13317 6824
rect 11037 6781 11093 6783
rect 11163 6781 11405 6783
rect 10985 6767 11093 6781
rect 11127 6767 11405 6781
rect 11037 6749 11093 6767
rect 11163 6749 11405 6767
rect 11439 6749 11717 6783
rect 11751 6749 12029 6783
rect 12063 6749 12341 6783
rect 12375 6749 12653 6783
rect 12687 6749 12965 6783
rect 12999 6749 13277 6783
rect 13311 6749 13317 6783
rect 11037 6715 11111 6749
rect 11163 6715 13317 6749
rect 10985 6708 13317 6715
rect 10985 6701 11093 6708
rect 11127 6701 11405 6708
rect 11037 6674 11093 6701
rect 11163 6674 11405 6701
rect 11439 6674 11717 6708
rect 11751 6674 12029 6708
rect 12063 6674 12341 6708
rect 12375 6674 12653 6708
rect 12687 6674 12965 6708
rect 12999 6674 13277 6708
rect 13311 6674 13317 6708
rect 11037 6649 11111 6674
rect 11163 6649 13317 6674
rect 10985 6635 13317 6649
rect 11037 6633 11111 6635
rect 11163 6633 13317 6635
rect 11037 6599 11093 6633
rect 11163 6599 11405 6633
rect 11439 6599 11717 6633
rect 11751 6599 12029 6633
rect 12063 6599 12341 6633
rect 12375 6599 12653 6633
rect 12687 6599 12965 6633
rect 12999 6599 13277 6633
rect 13311 6599 13317 6633
rect 11037 6583 11111 6599
rect 11163 6583 13317 6599
rect 10985 6569 13317 6583
rect 11037 6558 11111 6569
rect 11163 6558 13317 6569
rect 11037 6524 11093 6558
rect 11163 6524 11405 6558
rect 11439 6524 11717 6558
rect 11751 6524 12029 6558
rect 12063 6524 12341 6558
rect 12375 6524 12653 6558
rect 12687 6524 12965 6558
rect 12999 6524 13277 6558
rect 13311 6524 13317 6558
rect 11037 6517 11111 6524
rect 11163 6517 13317 6524
rect 10985 6511 13317 6517
rect 13381 7139 13427 7179
rect 13381 7105 13387 7139
rect 13421 7105 13427 7139
rect 13381 7065 13427 7105
rect 13381 7031 13387 7065
rect 13421 7031 13427 7065
rect 13381 6991 13427 7031
rect 13381 6957 13387 6991
rect 13421 6957 13427 6991
rect 13381 6917 13427 6957
rect 13381 6883 13387 6917
rect 13421 6883 13427 6917
rect 13381 6843 13427 6883
rect 13381 6809 13387 6843
rect 13421 6809 13427 6843
rect 13381 6769 13427 6809
rect 13381 6735 13387 6769
rect 13421 6735 13427 6769
rect 13381 6695 13427 6735
rect 13381 6661 13387 6695
rect 13421 6661 13427 6695
rect 13381 6621 13427 6661
rect 13381 6587 13387 6621
rect 13421 6587 13427 6621
rect 13381 6547 13427 6587
rect 13381 6513 13387 6547
rect 13421 6513 13427 6547
rect 10458 6428 10648 6487
rect 13381 6473 13427 6513
tri 13353 6440 13381 6468 se
rect 13381 6440 13387 6473
rect 10458 6394 10464 6428
rect 10498 6394 10536 6428
rect 10570 6394 10608 6428
rect 10642 6394 10648 6428
rect 10458 6350 10648 6394
rect 10786 6439 10832 6440
tri 10832 6439 10833 6440 sw
tri 13352 6439 13353 6440 se
rect 13353 6439 13387 6440
rect 13421 6439 13427 6473
rect 10786 6409 10833 6439
tri 10833 6409 10863 6439 sw
tri 13322 6409 13352 6439 se
rect 13352 6409 13427 6439
rect 10786 6407 10863 6409
tri 10863 6407 10865 6409 sw
tri 13320 6407 13322 6409 se
rect 13322 6407 13427 6409
rect 10786 6401 13427 6407
rect 10786 6367 10864 6401
rect 10898 6367 10937 6401
rect 10971 6367 11010 6401
rect 11044 6367 11083 6401
rect 11117 6367 11155 6401
rect 11189 6367 11227 6401
rect 11261 6367 11299 6401
rect 11333 6367 11371 6401
rect 11405 6367 11443 6401
rect 11477 6367 11515 6401
rect 11549 6367 11587 6401
rect 11621 6367 11659 6401
rect 11693 6367 11731 6401
rect 11765 6367 11803 6401
rect 11837 6367 11875 6401
rect 11909 6367 11947 6401
rect 11981 6367 12019 6401
rect 12053 6367 12091 6401
rect 12125 6367 12163 6401
rect 12197 6367 12235 6401
rect 12269 6367 12307 6401
rect 12341 6367 12379 6401
rect 12413 6367 12451 6401
rect 12485 6367 12523 6401
rect 12557 6367 12595 6401
rect 12629 6367 12667 6401
rect 12701 6367 12739 6401
rect 12773 6367 12811 6401
rect 12845 6367 12883 6401
rect 12917 6367 12955 6401
rect 12989 6367 13027 6401
rect 13061 6367 13099 6401
rect 13133 6367 13171 6401
rect 13205 6367 13243 6401
rect 13277 6367 13315 6401
rect 13349 6367 13427 6401
rect 10786 6361 13427 6367
rect 13589 8096 13779 8108
rect 13589 8062 13595 8096
rect 13629 8062 13667 8096
rect 13701 8062 13739 8096
rect 13773 8062 13779 8096
rect 13589 8022 13779 8062
rect 13589 7988 13595 8022
rect 13629 7988 13667 8022
rect 13701 7988 13739 8022
rect 13773 7988 13779 8022
rect 13589 7948 13779 7988
rect 13589 7914 13595 7948
rect 13629 7914 13667 7948
rect 13701 7914 13739 7948
rect 13773 7914 13779 7948
rect 13589 7874 13779 7914
rect 13589 7840 13595 7874
rect 13629 7840 13667 7874
rect 13701 7840 13739 7874
rect 13773 7840 13779 7874
rect 13589 7800 13779 7840
rect 13589 7766 13595 7800
rect 13629 7766 13667 7800
rect 13701 7766 13739 7800
rect 13773 7766 13779 7800
rect 13589 7726 13779 7766
rect 13589 7692 13595 7726
rect 13629 7692 13667 7726
rect 13701 7692 13739 7726
rect 13773 7692 13779 7726
rect 13589 7652 13779 7692
rect 13589 7618 13595 7652
rect 13629 7618 13667 7652
rect 13701 7618 13739 7652
rect 13773 7618 13779 7652
rect 13589 7578 13779 7618
rect 13589 7544 13595 7578
rect 13629 7544 13667 7578
rect 13701 7544 13739 7578
rect 13773 7544 13779 7578
rect 13589 7504 13779 7544
rect 13589 7470 13595 7504
rect 13629 7470 13667 7504
rect 13701 7470 13739 7504
rect 13773 7470 13779 7504
rect 13589 7431 13779 7470
rect 13589 7430 13667 7431
rect 13589 7396 13595 7430
rect 13629 7397 13667 7430
rect 13701 7397 13739 7431
rect 13773 7397 13779 7431
rect 13629 7396 13779 7397
rect 13589 7358 13779 7396
rect 13589 7356 13667 7358
rect 13589 7322 13595 7356
rect 13629 7324 13667 7356
rect 13701 7324 13739 7358
rect 13773 7324 13779 7358
rect 13629 7322 13779 7324
rect 13589 7285 13779 7322
rect 13589 7283 13667 7285
rect 13589 7249 13595 7283
rect 13629 7251 13667 7283
rect 13701 7251 13739 7285
rect 13773 7251 13779 7285
rect 13629 7249 13779 7251
rect 13589 7212 13779 7249
rect 13589 7210 13667 7212
rect 13589 7176 13595 7210
rect 13629 7178 13667 7210
rect 13701 7178 13739 7212
rect 13773 7178 13779 7212
rect 13629 7176 13779 7178
rect 13589 7139 13779 7176
rect 13589 7137 13667 7139
rect 13589 7103 13595 7137
rect 13629 7105 13667 7137
rect 13701 7105 13739 7139
rect 13773 7105 13779 7139
rect 13629 7103 13779 7105
rect 13589 7066 13779 7103
rect 13589 7064 13667 7066
rect 13589 7030 13595 7064
rect 13629 7032 13667 7064
rect 13701 7032 13739 7066
rect 13773 7032 13779 7066
rect 13629 7030 13779 7032
rect 13589 6993 13779 7030
rect 13589 6991 13667 6993
rect 13589 6957 13595 6991
rect 13629 6959 13667 6991
rect 13701 6959 13739 6993
rect 13773 6959 13779 6993
rect 13629 6957 13779 6959
rect 13589 6920 13779 6957
rect 13589 6918 13667 6920
rect 13589 6884 13595 6918
rect 13629 6886 13667 6918
rect 13701 6886 13739 6920
rect 13773 6886 13779 6920
rect 13629 6884 13779 6886
rect 13589 6847 13779 6884
rect 13589 6845 13667 6847
rect 13589 6811 13595 6845
rect 13629 6813 13667 6845
rect 13701 6813 13739 6847
rect 13773 6813 13779 6847
rect 13629 6811 13779 6813
rect 13589 6774 13779 6811
rect 13589 6772 13667 6774
rect 13589 6738 13595 6772
rect 13629 6740 13667 6772
rect 13701 6740 13739 6774
rect 13773 6740 13779 6774
rect 13629 6738 13779 6740
rect 13589 6701 13779 6738
rect 13589 6699 13667 6701
rect 13589 6665 13595 6699
rect 13629 6667 13667 6699
rect 13701 6667 13739 6701
rect 13773 6667 13779 6701
rect 13629 6665 13779 6667
rect 13589 6628 13779 6665
rect 13589 6626 13667 6628
rect 13589 6592 13595 6626
rect 13629 6594 13667 6626
rect 13701 6594 13739 6628
rect 13773 6594 13779 6628
rect 13629 6592 13779 6594
rect 13589 6555 13779 6592
rect 13589 6553 13667 6555
rect 13589 6519 13595 6553
rect 13629 6521 13667 6553
rect 13701 6521 13739 6555
rect 13773 6521 13779 6555
rect 13629 6519 13779 6521
rect 13589 6482 13779 6519
rect 13589 6480 13667 6482
rect 13589 6446 13595 6480
rect 13629 6448 13667 6480
rect 13701 6448 13739 6482
rect 13773 6448 13779 6482
rect 13629 6446 13779 6448
rect 13589 6409 13779 6446
rect 13589 6407 13667 6409
rect 13589 6373 13595 6407
rect 13629 6375 13667 6407
rect 13701 6375 13739 6409
rect 13773 6375 13779 6409
rect 13629 6373 13779 6375
rect 10458 6316 10464 6350
rect 10498 6316 10536 6350
rect 10570 6348 10648 6350
rect 10570 6316 10608 6348
rect 10458 6314 10608 6316
rect 10642 6314 10648 6348
rect 10458 6272 10648 6314
rect 10458 6238 10464 6272
rect 10498 6238 10536 6272
rect 10570 6268 10648 6272
rect 10570 6238 10608 6268
rect 10458 6234 10608 6238
rect 10642 6234 10648 6268
rect 13589 6336 13779 6373
rect 13589 6334 13667 6336
rect 13589 6300 13595 6334
rect 13629 6302 13667 6334
rect 13701 6302 13739 6336
rect 13773 6302 13779 6336
rect 13629 6300 13779 6302
rect 13589 6263 13779 6300
rect 13589 6261 13667 6263
tri 13572 6238 13589 6255 se
rect 13589 6238 13595 6261
rect 10458 6227 10648 6234
tri 10648 6227 10659 6238 sw
tri 13561 6227 13572 6238 se
rect 13572 6227 13595 6238
rect 13629 6229 13667 6261
rect 13701 6229 13739 6263
rect 13773 6229 13779 6263
rect 13629 6227 13779 6229
rect 10458 6194 10659 6227
tri 10659 6194 10692 6227 sw
tri 13528 6194 13561 6227 se
rect 13561 6194 13779 6227
rect 10458 6160 10464 6194
rect 10498 6160 10536 6194
rect 10570 6190 13779 6194
rect 10570 6188 13667 6190
rect 10570 6160 10608 6188
rect 10458 6116 10608 6160
rect 11074 6154 11113 6188
rect 11147 6154 11186 6188
rect 11220 6154 11259 6188
rect 11293 6154 11332 6188
rect 11366 6154 11405 6188
rect 11439 6154 11478 6188
rect 11512 6154 11551 6188
rect 11585 6154 11624 6188
rect 11658 6154 11697 6188
rect 11731 6154 11770 6188
rect 11804 6154 11843 6188
rect 11877 6154 11916 6188
rect 11950 6154 11989 6188
rect 12023 6154 12062 6188
rect 12096 6154 12135 6188
rect 12169 6154 12208 6188
rect 12242 6154 12281 6188
rect 12315 6154 12354 6188
rect 12388 6154 12427 6188
rect 12461 6154 12500 6188
rect 12534 6154 12573 6188
rect 12607 6154 12646 6188
rect 12680 6154 12719 6188
rect 12753 6154 12792 6188
rect 12826 6154 12865 6188
rect 12899 6154 12938 6188
rect 12972 6154 13011 6188
rect 13045 6154 13084 6188
rect 13118 6154 13157 6188
rect 13191 6154 13230 6188
rect 13264 6154 13303 6188
rect 13337 6154 13376 6188
rect 13410 6154 13449 6188
rect 13483 6154 13522 6188
rect 13556 6154 13595 6188
rect 13629 6156 13667 6188
rect 13701 6156 13739 6190
rect 13773 6156 13779 6190
rect 13629 6154 13779 6156
rect 11074 6117 13779 6154
rect 11074 6116 13739 6117
rect 10458 6082 10464 6116
rect 10498 6082 10536 6116
rect 10458 6010 10536 6082
rect 11146 6082 11185 6116
rect 11219 6082 11258 6116
rect 11292 6082 11331 6116
rect 11365 6082 11404 6116
rect 11438 6082 11477 6116
rect 11511 6082 11550 6116
rect 11584 6082 11623 6116
rect 11657 6082 11696 6116
rect 11730 6082 11769 6116
rect 11803 6082 11842 6116
rect 11876 6082 11915 6116
rect 11949 6082 11988 6116
rect 12022 6082 12061 6116
rect 12095 6082 12134 6116
rect 12168 6082 12207 6116
rect 12241 6082 12280 6116
rect 12314 6082 12353 6116
rect 12387 6082 12426 6116
rect 12460 6082 12499 6116
rect 12533 6082 12572 6116
rect 12606 6082 12645 6116
rect 12679 6082 12718 6116
rect 12752 6082 12791 6116
rect 12825 6082 12864 6116
rect 12898 6082 12937 6116
rect 12971 6082 13010 6116
rect 13044 6082 13083 6116
rect 13117 6082 13156 6116
rect 13190 6082 13229 6116
rect 13263 6082 13302 6116
rect 13336 6082 13375 6116
rect 13409 6082 13448 6116
rect 13482 6082 13521 6116
rect 13555 6082 13594 6116
rect 13628 6082 13667 6116
rect 13701 6083 13739 6116
rect 13773 6083 13779 6117
rect 13701 6082 13779 6083
rect 11146 6044 13779 6082
rect 11146 6010 11185 6044
rect 11219 6010 11258 6044
rect 11292 6010 11331 6044
rect 11365 6010 11404 6044
rect 11438 6010 11477 6044
rect 11511 6010 11550 6044
rect 11584 6010 11623 6044
rect 11657 6010 11696 6044
rect 11730 6010 11769 6044
rect 11803 6010 11842 6044
rect 11876 6010 11915 6044
rect 11949 6010 11988 6044
rect 12022 6010 12061 6044
rect 12095 6010 12134 6044
rect 12168 6010 12207 6044
rect 12241 6010 12280 6044
rect 12314 6010 12353 6044
rect 12387 6010 12426 6044
rect 12460 6010 12499 6044
rect 12533 6010 12572 6044
rect 12606 6010 12645 6044
rect 12679 6010 12718 6044
rect 12752 6010 12791 6044
rect 12825 6010 12864 6044
rect 12898 6010 12937 6044
rect 12971 6010 13010 6044
rect 13044 6010 13083 6044
rect 13117 6010 13156 6044
rect 13190 6010 13229 6044
rect 13263 6010 13302 6044
rect 13336 6010 13375 6044
rect 13409 6010 13448 6044
rect 13482 6010 13521 6044
rect 13555 6010 13594 6044
rect 13628 6010 13667 6044
rect 13701 6010 13779 6044
rect 10458 6004 13779 6010
tri 13779 6004 13809 6034 sw
rect 10458 5950 13809 6004
rect 10458 5916 10473 5950
rect 10507 5916 10546 5950
rect 10580 5916 10619 5950
rect 10653 5916 10692 5950
rect 10726 5916 10765 5950
rect 10799 5916 10838 5950
rect 10872 5916 10911 5950
rect 10945 5916 10984 5950
rect 11018 5916 11057 5950
rect 11091 5916 11130 5950
rect 11164 5916 11203 5950
rect 11237 5916 11276 5950
rect 11310 5916 11349 5950
rect 11383 5916 11422 5950
rect 11456 5916 11495 5950
rect 11529 5916 11568 5950
rect 11602 5916 11641 5950
rect 11675 5916 11714 5950
rect 11748 5916 11787 5950
rect 11821 5916 11860 5950
rect 11894 5916 11933 5950
rect 11967 5916 12005 5950
rect 12039 5916 12077 5950
rect 12111 5916 12149 5950
rect 12183 5916 12221 5950
rect 12255 5916 12293 5950
rect 12327 5916 12365 5950
rect 12399 5916 12437 5950
rect 12471 5916 12509 5950
rect 12543 5916 12581 5950
rect 12615 5916 12653 5950
rect 12687 5916 12725 5950
rect 12759 5916 12797 5950
rect 12831 5916 12869 5950
rect 12903 5916 12941 5950
rect 12975 5916 13013 5950
rect 13047 5916 13085 5950
rect 13119 5916 13157 5950
rect 13191 5916 13229 5950
rect 13263 5916 13301 5950
rect 13335 5916 13373 5950
rect 13407 5916 13445 5950
rect 13479 5916 13517 5950
rect 13551 5916 13589 5950
rect 13623 5916 13661 5950
rect 13695 5916 13733 5950
rect 13767 5916 13809 5950
rect 10458 5853 13809 5916
tri 13809 5853 13960 6004 sw
rect 10458 5847 14132 5853
rect 10458 5819 10904 5847
tri 10458 5775 10502 5819 ne
rect 10502 5775 10904 5819
rect 9456 5764 9534 5766
rect 9456 5730 9462 5764
rect 9496 5732 9534 5764
rect 9568 5732 9606 5766
rect 9640 5732 9646 5766
tri 10502 5741 10536 5775 ne
rect 10536 5741 10832 5775
rect 10866 5741 10904 5775
rect 12594 5813 12633 5847
rect 12667 5813 12706 5847
rect 12740 5813 12779 5847
rect 12813 5813 12852 5847
rect 12886 5813 12925 5847
rect 12959 5813 12998 5847
rect 13032 5813 13071 5847
rect 13105 5813 13144 5847
rect 13178 5813 13217 5847
rect 13251 5813 13290 5847
rect 13324 5813 13363 5847
rect 13397 5813 13436 5847
rect 13470 5813 13509 5847
rect 13543 5813 13582 5847
rect 13616 5813 13655 5847
rect 13689 5813 13728 5847
rect 13762 5813 13801 5847
rect 13835 5813 13874 5847
rect 13908 5813 13947 5847
rect 13981 5813 14020 5847
rect 14054 5813 14132 5847
rect 12594 5775 14132 5813
rect 12594 5741 12633 5775
rect 12667 5741 12706 5775
rect 12740 5741 12779 5775
rect 12813 5741 12852 5775
rect 12886 5741 12925 5775
rect 12959 5741 12998 5775
rect 13032 5741 13071 5775
rect 13105 5741 13144 5775
rect 13178 5741 13217 5775
rect 13251 5741 13290 5775
rect 13324 5741 13363 5775
rect 13397 5741 13436 5775
rect 13470 5741 13509 5775
rect 13543 5741 13582 5775
rect 13616 5741 13655 5775
rect 13689 5741 13728 5775
rect 13762 5741 13801 5775
rect 13835 5741 13874 5775
rect 13908 5741 13947 5775
rect 13981 5741 14020 5775
rect 9496 5730 9646 5732
rect 9456 5690 9646 5730
tri 10536 5700 10577 5741 ne
rect 10577 5700 10976 5741
tri 10577 5699 10578 5700 ne
rect 10578 5699 10904 5700
rect 9456 5685 9534 5690
tri 810 5651 833 5674 sw
tri 9446 5651 9456 5661 se
rect 9456 5651 9462 5685
rect 9496 5656 9534 5685
rect 9568 5656 9606 5690
rect 9640 5656 9646 5690
tri 10578 5665 10612 5699 ne
rect 10612 5665 10832 5699
rect 10866 5666 10904 5699
rect 10938 5669 10976 5700
rect 12522 5703 14020 5741
rect 12522 5669 12561 5703
rect 12595 5669 12634 5703
rect 12668 5669 12707 5703
rect 12741 5669 12780 5703
rect 12814 5669 12853 5703
rect 12887 5669 12926 5703
rect 12960 5669 12999 5703
rect 13033 5669 13072 5703
rect 13106 5669 13145 5703
rect 13179 5669 13218 5703
rect 13252 5669 13291 5703
rect 13325 5669 13364 5703
rect 13398 5669 13437 5703
rect 13471 5669 13510 5703
rect 13544 5669 13583 5703
rect 13617 5669 13656 5703
rect 13690 5669 13729 5703
rect 13763 5669 13802 5703
rect 13836 5669 13875 5703
rect 13909 5669 13948 5703
rect 10938 5666 13948 5669
rect 10866 5665 13948 5666
rect 9496 5651 9646 5656
rect 804 5645 833 5651
rect 620 5607 749 5617
rect 620 5573 626 5607
rect 660 5604 698 5607
rect 683 5573 698 5604
rect 732 5606 749 5607
rect 801 5628 833 5645
tri 833 5628 856 5651 sw
tri 9423 5628 9446 5651 se
rect 9446 5628 9646 5651
tri 10612 5628 10649 5665 ne
rect 10649 5663 13948 5665
rect 10649 5628 11053 5663
rect 801 5625 856 5628
tri 856 5625 859 5628 sw
tri 9420 5625 9423 5628 se
rect 9423 5625 9646 5628
tri 10649 5625 10652 5628 ne
rect 10652 5625 10976 5628
rect 801 5623 859 5625
tri 859 5623 861 5625 sw
tri 9418 5623 9420 5625 se
rect 9420 5623 9646 5625
tri 10652 5623 10654 5625 ne
rect 10654 5623 10904 5625
rect 801 5614 861 5623
tri 861 5614 870 5623 sw
tri 9409 5614 9418 5623 se
rect 9418 5614 9646 5623
rect 801 5612 870 5614
tri 870 5612 872 5614 sw
tri 9407 5612 9409 5614 se
rect 9409 5612 9534 5614
rect 801 5606 9534 5612
rect 732 5593 770 5606
rect 732 5573 749 5593
rect 620 5552 631 5573
rect 683 5552 749 5573
rect 620 5541 749 5552
rect 5700 5572 5739 5606
rect 5773 5572 5812 5606
rect 5846 5572 5885 5606
rect 5919 5572 5958 5606
rect 5992 5572 6031 5606
rect 6065 5572 6104 5606
rect 6138 5572 6177 5606
rect 6211 5572 6250 5606
rect 6284 5572 6323 5606
rect 6357 5572 6396 5606
rect 6430 5572 6469 5606
rect 6503 5572 6542 5606
rect 6576 5572 6615 5606
rect 6649 5572 6688 5606
rect 6722 5572 6761 5606
rect 6795 5572 6834 5606
rect 6868 5572 6907 5606
rect 6941 5572 6980 5606
rect 7014 5572 7053 5606
rect 7087 5572 7126 5606
rect 7160 5572 7199 5606
rect 7233 5572 7272 5606
rect 7306 5572 7345 5606
rect 7379 5572 7418 5606
rect 7452 5572 7491 5606
rect 7525 5572 7564 5606
rect 7598 5572 7637 5606
rect 7671 5572 7710 5606
rect 7744 5572 7783 5606
rect 7817 5572 7856 5606
rect 7890 5572 7929 5606
rect 7963 5572 8002 5606
rect 8036 5572 8075 5606
rect 8109 5572 8148 5606
rect 8182 5572 8221 5606
rect 8255 5572 8294 5606
rect 8328 5572 8367 5606
rect 8401 5572 8440 5606
rect 8474 5572 8513 5606
rect 8547 5572 8586 5606
rect 8620 5572 8659 5606
rect 8693 5572 8732 5606
rect 8766 5572 8805 5606
rect 8839 5572 8878 5606
rect 8912 5572 8951 5606
rect 8985 5572 9024 5606
rect 9058 5572 9097 5606
rect 9131 5572 9170 5606
rect 9204 5572 9243 5606
rect 9277 5572 9316 5606
rect 9350 5572 9389 5606
rect 9423 5572 9462 5606
rect 9496 5580 9534 5606
rect 9568 5580 9606 5614
rect 9640 5580 9646 5614
tri 10654 5589 10688 5623 ne
rect 10688 5589 10832 5623
rect 10866 5591 10904 5623
rect 10938 5594 10976 5625
rect 11010 5594 11053 5628
rect 10938 5591 11053 5594
rect 10866 5589 11053 5591
rect 9496 5572 9646 5580
rect 620 5539 770 5541
rect 620 5534 631 5539
rect 683 5534 770 5539
rect 5700 5538 9646 5572
tri 10688 5553 10724 5589 ne
rect 10724 5553 11053 5589
tri 10724 5550 10727 5553 ne
rect 10727 5550 10976 5553
tri 10727 5548 10729 5550 ne
rect 10729 5548 10904 5550
rect 5700 5534 9606 5538
rect 620 5500 626 5534
rect 620 5487 631 5500
rect 683 5487 698 5534
rect 620 5475 698 5487
rect 5772 5500 5811 5534
rect 5845 5500 5884 5534
rect 5918 5500 5957 5534
rect 5991 5500 6030 5534
rect 6064 5500 6103 5534
rect 6137 5500 6176 5534
rect 6210 5500 6249 5534
rect 6283 5500 6322 5534
rect 6356 5500 6395 5534
rect 6429 5500 6468 5534
rect 6502 5500 6541 5534
rect 6575 5500 6614 5534
rect 6648 5500 6687 5534
rect 6721 5500 6760 5534
rect 6794 5500 6833 5534
rect 6867 5500 6906 5534
rect 6940 5500 6979 5534
rect 7013 5500 7052 5534
rect 7086 5500 7125 5534
rect 7159 5500 7198 5534
rect 7232 5500 7271 5534
rect 7305 5500 7344 5534
rect 7378 5500 7417 5534
rect 7451 5500 7490 5534
rect 7524 5500 7563 5534
rect 7597 5500 7636 5534
rect 7670 5500 7709 5534
rect 7743 5500 7782 5534
rect 7816 5500 7855 5534
rect 7889 5500 7928 5534
rect 7962 5500 8001 5534
rect 8035 5500 8074 5534
rect 8108 5500 8147 5534
rect 8181 5500 8220 5534
rect 8254 5500 8293 5534
rect 8327 5500 8366 5534
rect 8400 5500 8439 5534
rect 8473 5500 8512 5534
rect 8546 5500 8585 5534
rect 8619 5500 8658 5534
rect 8692 5500 8731 5534
rect 8765 5500 8804 5534
rect 8838 5500 8877 5534
rect 8911 5500 8950 5534
rect 8984 5500 9023 5534
rect 9057 5500 9096 5534
rect 9130 5500 9169 5534
rect 9203 5500 9242 5534
rect 9276 5500 9315 5534
rect 9349 5500 9388 5534
rect 9422 5500 9461 5534
rect 9495 5500 9534 5534
rect 9568 5504 9606 5534
rect 9640 5504 9646 5538
tri 10729 5514 10763 5548 ne
rect 10763 5514 10832 5548
rect 10866 5516 10904 5548
rect 10938 5519 10976 5550
rect 11010 5537 11053 5553
tri 11053 5537 11179 5663 nw
tri 13881 5602 13942 5663 ne
rect 11364 5537 12562 5543
rect 11010 5519 11019 5537
rect 10938 5516 11019 5519
rect 10866 5514 11019 5516
rect 9568 5500 9646 5504
tri 10763 5503 10774 5514 ne
rect 10774 5503 11019 5514
tri 11019 5503 11053 5537 nw
rect 11364 5503 11468 5537
rect 11502 5503 11540 5537
rect 11574 5503 11612 5537
rect 11646 5503 11684 5537
rect 11718 5503 11756 5537
rect 11790 5503 11828 5537
rect 11862 5503 11900 5537
rect 11934 5503 11972 5537
rect 12006 5503 12044 5537
rect 12078 5503 12116 5537
rect 12150 5503 12188 5537
rect 12222 5503 12260 5537
rect 12294 5503 12332 5537
rect 12366 5503 12404 5537
rect 12438 5503 12476 5537
rect 12510 5503 12562 5537
rect 620 5423 697 5475
rect 5772 5462 9646 5500
tri 10774 5478 10799 5503 ne
rect 10799 5478 11016 5503
tri 11016 5500 11019 5503 nw
tri 10799 5475 10802 5478 ne
rect 10802 5475 10976 5478
tri 10802 5473 10804 5475 ne
rect 10804 5473 10904 5475
rect 5772 5428 5811 5462
rect 5845 5428 5884 5462
rect 5918 5428 5957 5462
rect 5991 5428 6030 5462
rect 6064 5428 6103 5462
rect 6137 5428 6176 5462
rect 6210 5428 6249 5462
rect 6283 5428 6322 5462
rect 6356 5428 6395 5462
rect 6429 5428 6468 5462
rect 6502 5428 6541 5462
rect 6575 5428 6614 5462
rect 6648 5428 6687 5462
rect 6721 5428 6760 5462
rect 6794 5428 6833 5462
rect 6867 5428 6906 5462
rect 6940 5428 6979 5462
rect 7013 5428 7052 5462
rect 7086 5428 7125 5462
rect 7159 5428 7198 5462
rect 7232 5428 7271 5462
rect 7305 5428 7344 5462
rect 7378 5428 7417 5462
rect 7451 5428 7490 5462
rect 7524 5428 7563 5462
rect 7597 5428 7636 5462
rect 7670 5428 7709 5462
rect 7743 5428 7782 5462
rect 7816 5428 7855 5462
rect 7889 5428 7928 5462
rect 7962 5428 8001 5462
rect 8035 5428 8074 5462
rect 8108 5428 8147 5462
rect 8181 5428 8220 5462
rect 8254 5428 8293 5462
rect 8327 5428 8366 5462
rect 8400 5428 8439 5462
rect 8473 5428 8512 5462
rect 8546 5428 8585 5462
rect 8619 5428 8658 5462
rect 8692 5428 8731 5462
rect 8765 5428 8804 5462
rect 8838 5428 8877 5462
rect 8911 5428 8950 5462
rect 8984 5428 9023 5462
rect 9057 5428 9096 5462
rect 9130 5428 9169 5462
rect 9203 5428 9242 5462
rect 9276 5428 9315 5462
rect 9349 5428 9388 5462
rect 9422 5428 9461 5462
rect 9495 5428 9534 5462
rect 9568 5428 9646 5462
tri 10804 5451 10826 5473 ne
rect 749 5423 763 5428
rect 815 5423 829 5428
rect 881 5423 895 5428
rect 947 5423 961 5428
rect 1013 5423 1027 5428
rect 1079 5423 1094 5428
rect 1146 5423 1161 5428
rect 1213 5423 1228 5428
rect 1280 5423 1295 5428
rect 1347 5423 1362 5428
rect 1414 5423 1429 5428
rect 1481 5423 1496 5428
rect 1548 5423 1563 5428
rect 1615 5423 1630 5428
rect 1682 5423 1697 5428
rect 1749 5423 1764 5428
rect 1816 5423 1831 5428
rect 1883 5423 1898 5428
rect 1950 5423 1965 5428
rect 2017 5423 2032 5428
rect 2084 5423 2099 5428
rect 2151 5423 2166 5428
rect 2218 5423 9646 5428
rect 620 5422 9646 5423
rect 10826 5439 10832 5473
rect 10866 5441 10904 5473
rect 10938 5444 10976 5475
rect 11010 5444 11016 5478
rect 10938 5441 11016 5444
rect 10866 5439 11016 5441
tri 437 5403 447 5413 sw
rect 10826 5403 11016 5439
rect 357 5400 447 5403
tri 447 5400 450 5403 sw
rect 10826 5400 10976 5403
rect 357 5398 450 5400
tri 450 5398 452 5400 sw
rect 10826 5398 10904 5400
rect 357 5379 452 5398
tri 452 5379 471 5398 sw
rect 357 5365 4040 5379
rect 357 5313 3854 5365
rect 3906 5313 3918 5365
rect 3970 5313 3982 5365
rect 4034 5313 4040 5365
rect 357 5299 4040 5313
rect 10826 5364 10832 5398
rect 10866 5366 10904 5398
rect 10938 5369 10976 5400
rect 11010 5369 11016 5403
rect 10938 5366 11016 5369
rect 10866 5364 11016 5366
rect 10826 5328 11016 5364
rect 10826 5325 10976 5328
rect 10826 5323 10904 5325
rect 10826 5289 10832 5323
rect 10866 5291 10904 5323
rect 10938 5294 10976 5325
rect 11010 5294 11016 5328
rect 10938 5291 11016 5294
rect 10866 5289 11016 5291
rect 10826 5253 11016 5289
rect 10826 5250 10976 5253
rect 10826 5248 10904 5250
rect 10826 5214 10832 5248
rect 10866 5216 10904 5248
rect 10938 5219 10976 5250
rect 11010 5219 11016 5253
rect 10938 5216 11016 5219
rect 10866 5214 11016 5216
rect 10826 5178 11016 5214
rect 10826 5175 10976 5178
rect 10826 5173 10904 5175
rect 10826 5139 10832 5173
rect 10866 5141 10904 5173
rect 10938 5144 10976 5175
rect 11010 5144 11016 5178
rect 10938 5141 11016 5144
rect 10866 5139 11016 5141
rect 10826 5103 11016 5139
rect 10826 5100 10976 5103
rect 10826 5098 10904 5100
rect 10826 5064 10832 5098
rect 10866 5066 10904 5098
rect 10938 5069 10976 5100
rect 11010 5069 11016 5103
rect 10938 5066 11016 5069
rect 10866 5064 11016 5066
rect 10826 5028 11016 5064
rect 10826 5025 10976 5028
rect 10826 5023 10904 5025
rect 10826 4989 10832 5023
rect 10866 4991 10904 5023
rect 10938 4994 10976 5025
rect 11010 4994 11016 5028
rect 10938 4991 11016 4994
rect 10866 4989 11016 4991
rect 10826 4953 11016 4989
rect 10826 4950 10976 4953
rect 10826 4948 10904 4950
rect 10826 4914 10832 4948
rect 10866 4916 10904 4948
rect 10938 4919 10976 4950
rect 11010 4919 11016 4953
rect 10938 4916 11016 4919
rect 10866 4914 11016 4916
rect 10826 4878 11016 4914
rect 10826 4875 10976 4878
rect 10826 4873 10904 4875
tri 10805 4839 10826 4860 se
rect 10826 4839 10832 4873
rect 10866 4841 10904 4873
rect 10938 4844 10976 4875
rect 11010 4844 11016 4878
rect 10938 4841 11016 4844
rect 10866 4839 11016 4841
tri 10796 4830 10805 4839 se
rect 10805 4830 11016 4839
tri 10780 4814 10796 4830 se
rect 10796 4814 11016 4830
tri 10769 4803 10780 4814 se
rect 10780 4803 11016 4814
rect 11364 5497 12562 5503
rect 11364 5462 11410 5497
tri 11410 5463 11444 5497 nw
tri 12482 5463 12516 5497 ne
rect 11364 5428 11370 5462
rect 11404 5428 11410 5462
rect 11364 5390 11410 5428
rect 11364 5356 11370 5390
rect 11404 5356 11410 5390
rect 11364 5318 11410 5356
rect 12516 5462 12562 5497
rect 12516 5428 12522 5462
rect 12556 5428 12562 5462
rect 12516 5390 12562 5428
rect 12516 5356 12522 5390
rect 12556 5356 12562 5390
tri 11410 5318 11412 5320 sw
tri 12514 5318 12516 5320 se
rect 12516 5318 12562 5356
rect 11364 5284 11370 5318
rect 11404 5286 11412 5318
tri 11412 5286 11444 5318 sw
tri 12482 5286 12514 5318 se
rect 12514 5286 12522 5318
rect 11404 5284 12522 5286
rect 12556 5284 12562 5318
rect 11364 5246 12562 5284
rect 11364 5212 11370 5246
rect 11404 5212 11517 5246
rect 11551 5212 12376 5246
rect 12410 5212 12522 5246
rect 12556 5212 12562 5246
rect 11364 5174 12562 5212
rect 11364 5140 11370 5174
rect 11404 5140 11517 5174
rect 11551 5140 12376 5174
rect 12410 5140 12522 5174
rect 12556 5140 12562 5174
rect 11364 5102 12562 5140
rect 11364 5068 11370 5102
rect 11404 5068 11517 5102
rect 11551 5068 12376 5102
rect 12410 5068 12522 5102
rect 12556 5068 12562 5102
rect 11364 5030 12562 5068
rect 11364 4996 11370 5030
rect 11404 4996 11517 5030
rect 11551 4996 12376 5030
rect 12410 4996 12522 5030
rect 12556 4996 12562 5030
rect 11364 4958 12562 4996
rect 11364 4924 11370 4958
rect 11404 4924 11517 4958
rect 11551 4924 12376 4958
rect 12410 4924 12522 4958
rect 12556 4924 12562 4958
rect 11364 4886 12562 4924
rect 11364 4852 11370 4886
rect 11404 4852 11517 4886
rect 11551 4852 12376 4886
rect 12410 4852 12522 4886
rect 12556 4852 12562 4886
rect 11364 4814 12562 4852
tri 10766 4800 10769 4803 se
rect 10769 4800 10976 4803
tri 10764 4798 10766 4800 se
rect 10766 4798 10904 4800
tri 10730 4764 10764 4798 se
rect 10764 4764 10832 4798
rect 10866 4766 10904 4798
rect 10938 4769 10976 4800
rect 11010 4769 11016 4803
tri 11340 4780 11364 4804 se
rect 11364 4780 11370 4814
rect 11404 4780 11517 4814
rect 11551 4780 12376 4814
rect 12410 4780 12522 4814
rect 12556 4780 12562 4814
rect 10938 4766 11016 4769
rect 10866 4764 11016 4766
tri 10723 4757 10730 4764 se
rect 10730 4757 11016 4764
tri 11317 4757 11340 4780 se
rect 11340 4757 12562 4780
tri 10708 4742 10723 4757 se
rect 10723 4742 11016 4757
tri 11302 4742 11317 4757 se
rect 11317 4742 12562 4757
tri 10694 4728 10708 4742 se
rect 10708 4728 11016 4742
tri 10692 4726 10694 4728 se
rect 10694 4726 10976 4728
tri 10689 4723 10692 4726 se
rect 10692 4723 10904 4726
tri 10655 4689 10689 4723 se
rect 10689 4689 10832 4723
rect 10866 4692 10904 4723
rect 10938 4694 10976 4726
rect 11010 4694 11016 4728
rect 10938 4692 11016 4694
rect 10866 4689 11016 4692
tri 10650 4684 10655 4689 se
rect 10655 4684 11016 4689
tri 10620 4654 10650 4684 se
rect 10650 4654 11016 4684
rect 2324 4653 11016 4654
rect 2324 4652 10976 4653
rect 2324 4648 10904 4652
rect 2324 4576 2402 4648
rect 10428 4614 10467 4648
rect 10501 4614 10540 4648
rect 10574 4614 10613 4648
rect 10647 4614 10686 4648
rect 10720 4614 10759 4648
rect 10793 4614 10832 4648
rect 10866 4618 10904 4648
rect 10938 4619 10976 4652
rect 11010 4619 11016 4653
rect 10938 4618 11016 4619
rect 10866 4614 11016 4618
rect 10428 4578 11016 4614
rect 10428 4576 10976 4578
rect 2324 4542 2330 4576
rect 2364 4542 2402 4576
rect 10500 4542 10539 4576
rect 10573 4542 10612 4576
rect 10646 4542 10685 4576
rect 10719 4542 10758 4576
rect 10792 4542 10831 4576
rect 10865 4542 10904 4576
rect 10938 4544 10976 4576
rect 11010 4544 11016 4578
rect 10938 4542 11016 4544
rect 2324 4503 2474 4542
rect 2324 4469 2330 4503
rect 2364 4469 2402 4503
rect 2436 4470 2474 4503
rect 10500 4504 11016 4542
rect 10500 4470 10539 4504
rect 10573 4470 10612 4504
rect 10646 4470 10685 4504
rect 10719 4470 10758 4504
rect 10792 4470 10831 4504
rect 10865 4470 10904 4504
rect 10938 4470 11016 4504
rect 2436 4469 11016 4470
rect 2324 4464 11016 4469
tri 11284 4724 11302 4742 se
rect 11302 4724 11370 4742
rect 11284 4708 11370 4724
rect 11404 4708 11517 4742
rect 11551 4708 12376 4742
rect 12410 4708 12522 4742
rect 12556 4708 12562 4742
rect 11284 4696 12562 4708
rect 13942 5453 13948 5663
rect 14126 5453 14132 5775
rect 13942 5414 14132 5453
rect 13942 5380 13948 5414
rect 13982 5380 14020 5414
rect 14054 5380 14092 5414
rect 14126 5380 14132 5414
rect 13942 5341 14132 5380
rect 13942 5307 13948 5341
rect 13982 5307 14020 5341
rect 14054 5307 14092 5341
rect 14126 5307 14132 5341
rect 13942 5268 14132 5307
rect 13942 5234 13948 5268
rect 13982 5234 14020 5268
rect 14054 5234 14092 5268
rect 14126 5234 14132 5268
rect 13942 5195 14132 5234
rect 13942 5161 13948 5195
rect 13982 5161 14020 5195
rect 14054 5161 14092 5195
rect 14126 5161 14132 5195
rect 13942 5122 14132 5161
rect 13942 5088 13948 5122
rect 13982 5088 14020 5122
rect 14054 5088 14092 5122
rect 14126 5088 14132 5122
rect 13942 5049 14132 5088
rect 13942 5015 13948 5049
rect 13982 5015 14020 5049
rect 14054 5015 14092 5049
rect 14126 5015 14132 5049
rect 13942 4976 14132 5015
rect 13942 4942 13948 4976
rect 13982 4942 14020 4976
rect 14054 4942 14092 4976
rect 14126 4942 14132 4976
rect 13942 4903 14132 4942
rect 13942 4869 13948 4903
rect 13982 4869 14020 4903
rect 14054 4869 14092 4903
rect 14126 4869 14132 4903
rect 13942 4830 14132 4869
rect 13942 4796 13948 4830
rect 13982 4796 14020 4830
rect 14054 4796 14092 4830
rect 14126 4796 14132 4830
rect 13942 4757 14132 4796
rect 13942 4723 13948 4757
rect 13982 4723 14020 4757
rect 14054 4723 14092 4757
rect 14126 4723 14132 4757
rect 11284 4684 11352 4696
tri 11352 4684 11364 4696 nw
rect 13942 4684 14132 4723
rect 11284 4650 11318 4684
tri 11318 4650 11352 4684 nw
rect 13942 4650 13948 4684
rect 13982 4650 14020 4684
rect 14054 4650 14092 4684
rect 14126 4650 14132 4684
rect 2324 4431 2514 4464
rect 2324 4430 2474 4431
rect 2324 4396 2330 4430
rect 2364 4396 2402 4430
rect 2436 4397 2474 4430
rect 2508 4397 2514 4431
tri 2514 4400 2578 4464 nw
rect 2436 4396 2514 4397
rect 2324 4358 2514 4396
rect 2324 4357 2474 4358
rect 2324 4323 2330 4357
rect 2364 4323 2402 4357
rect 2436 4324 2474 4357
rect 2508 4324 2514 4358
rect 2436 4323 2514 4324
rect 2324 4285 2514 4323
tri 11250 4299 11284 4333 se
rect 11284 4298 11312 4650
tri 11312 4644 11318 4650 nw
rect 13942 4611 14132 4650
rect 13942 4577 13948 4611
rect 13982 4577 14020 4611
rect 14054 4577 14092 4611
rect 14126 4577 14132 4611
rect 13942 4538 14132 4577
rect 13942 4504 13948 4538
rect 13982 4504 14020 4538
rect 14054 4504 14092 4538
rect 14126 4504 14132 4538
rect 13942 4492 14132 4504
tri 14642 4396 14676 4430 se
rect 14676 4396 14724 8162
rect 11362 4387 12564 4396
rect 11362 4353 11597 4387
rect 11631 4353 11669 4387
rect 11703 4353 11741 4387
rect 11775 4353 11813 4387
rect 11847 4353 11885 4387
rect 11919 4353 11957 4387
rect 11991 4353 12029 4387
rect 12063 4353 12101 4387
rect 12135 4353 12173 4387
rect 12207 4353 12245 4387
rect 12279 4353 12317 4387
rect 12351 4353 12564 4387
rect 11362 4344 12564 4353
rect 13716 4344 14724 4396
tri 14642 4333 14653 4344 ne
rect 14653 4333 14724 4344
tri 11312 4299 11346 4333 sw
tri 14653 4310 14676 4333 ne
rect 2324 4284 2474 4285
rect 2324 4250 2330 4284
rect 2364 4250 2402 4284
rect 2436 4251 2474 4284
rect 2508 4251 2514 4285
rect 11370 4253 12556 4299
rect 2436 4250 2514 4251
rect 2324 4212 2514 4250
rect 2324 4211 2474 4212
rect 2324 4177 2330 4211
rect 2364 4177 2402 4211
rect 2436 4178 2474 4211
rect 2508 4178 2514 4212
rect 2436 4177 2514 4178
rect 2324 4139 2514 4177
rect 2324 4138 2474 4139
rect 2324 4104 2330 4138
rect 2364 4104 2402 4138
rect 2436 4105 2474 4138
rect 2508 4105 2514 4139
rect 2436 4104 2514 4105
rect 2324 4066 2514 4104
rect 2324 4065 2474 4066
rect 2324 4031 2330 4065
rect 2364 4031 2402 4065
rect 2436 4032 2474 4065
rect 2508 4032 2514 4066
rect 2436 4031 2514 4032
rect 2324 3993 2514 4031
rect 13947 4247 14131 4259
rect 13947 4213 13953 4247
rect 13987 4213 14091 4247
rect 14125 4213 14131 4247
rect 13947 4172 14131 4213
rect 13947 4138 13953 4172
rect 13987 4138 14091 4172
rect 14125 4138 14131 4172
rect 13947 4097 14131 4138
rect 13947 4063 13953 4097
rect 13987 4063 14091 4097
rect 14125 4063 14131 4097
rect 13947 4022 14131 4063
rect 2324 3992 2474 3993
rect 2324 3958 2330 3992
rect 2364 3958 2402 3992
rect 2436 3959 2474 3992
rect 2508 3959 2514 3993
rect 2436 3958 2514 3959
rect 2324 3920 2514 3958
rect 2324 3919 2474 3920
rect 2324 3885 2330 3919
rect 2364 3885 2402 3919
rect 2436 3886 2474 3919
rect 2508 3886 2514 3920
rect 2436 3885 2514 3886
rect 2324 3847 2514 3885
rect 2324 3846 2474 3847
rect 2324 3812 2330 3846
rect 2364 3812 2402 3846
rect 2436 3813 2474 3846
rect 2508 3813 2514 3847
rect 2436 3812 2514 3813
rect 2324 3774 2514 3812
rect 2324 3773 2474 3774
rect 2324 3739 2330 3773
rect 2364 3739 2402 3773
rect 2436 3740 2474 3773
rect 2508 3740 2514 3774
rect 2436 3739 2514 3740
rect 2324 3701 2514 3739
rect 2324 3700 2474 3701
rect 2324 3666 2330 3700
rect 2364 3666 2402 3700
rect 2436 3667 2474 3700
rect 2508 3667 2514 3701
rect 2436 3666 2514 3667
rect 2324 3628 2514 3666
rect 2324 3627 2474 3628
rect 2324 3593 2330 3627
rect 2364 3593 2402 3627
rect 2436 3594 2474 3627
rect 2508 3594 2514 3628
rect 2436 3593 2514 3594
rect 2324 3555 2514 3593
rect 2324 3554 2474 3555
rect 2324 3520 2330 3554
rect 2364 3520 2402 3554
rect 2436 3521 2474 3554
rect 2508 3521 2514 3555
rect 2436 3520 2514 3521
rect 2324 3482 2514 3520
rect 2324 3481 2474 3482
rect 2324 3447 2330 3481
rect 2364 3447 2402 3481
rect 2436 3448 2474 3481
rect 2508 3448 2514 3482
rect 2765 4004 3832 4010
rect 2765 3952 2771 4004
rect 2823 3952 2838 4004
rect 2890 3952 2905 4004
rect 2957 3952 2972 4004
rect 3024 3952 3039 4004
rect 3091 3952 3106 4004
rect 3158 3952 3173 4004
rect 3225 3952 3240 4004
rect 3292 3952 3307 4004
rect 3359 3952 3374 4004
rect 3426 3952 3441 4004
rect 3493 3952 3508 4004
rect 3560 3952 3575 4004
rect 3627 3952 3642 4004
rect 3694 3952 3708 4004
rect 3760 3952 3774 4004
rect 3826 3952 3832 4004
rect 2765 3936 3832 3952
rect 2765 3884 2771 3936
rect 2823 3884 2838 3936
rect 2890 3884 2905 3936
rect 2957 3884 2972 3936
rect 3024 3884 3039 3936
rect 3091 3884 3106 3936
rect 3158 3884 3173 3936
rect 3225 3884 3240 3936
rect 3292 3884 3307 3936
rect 3359 3884 3374 3936
rect 3426 3884 3441 3936
rect 3493 3884 3508 3936
rect 3560 3884 3575 3936
rect 3627 3884 3642 3936
rect 3694 3884 3708 3936
rect 3760 3884 3774 3936
rect 3826 3884 3832 3936
rect 2765 3868 3832 3884
rect 2765 3816 2771 3868
rect 2823 3816 2838 3868
rect 2890 3816 2905 3868
rect 2957 3816 2972 3868
rect 3024 3816 3039 3868
rect 3091 3816 3106 3868
rect 3158 3816 3173 3868
rect 3225 3816 3240 3868
rect 3292 3816 3307 3868
rect 3359 3816 3374 3868
rect 3426 3816 3441 3868
rect 3493 3816 3508 3868
rect 3560 3816 3575 3868
rect 3627 3816 3642 3868
rect 3694 3816 3708 3868
rect 3760 3816 3774 3868
rect 3826 3816 3832 3868
rect 2765 3800 3832 3816
rect 2765 3748 2771 3800
rect 2823 3748 2838 3800
rect 2890 3748 2905 3800
rect 2957 3748 2972 3800
rect 3024 3748 3039 3800
rect 3091 3748 3106 3800
rect 3158 3748 3173 3800
rect 3225 3748 3240 3800
rect 3292 3748 3307 3800
rect 3359 3748 3374 3800
rect 3426 3748 3441 3800
rect 3493 3748 3508 3800
rect 3560 3748 3575 3800
rect 3627 3748 3642 3800
rect 3694 3748 3708 3800
rect 3760 3748 3774 3800
rect 3826 3748 3832 3800
rect 2765 3732 3832 3748
rect 2765 3680 2771 3732
rect 2823 3680 2838 3732
rect 2890 3680 2905 3732
rect 2957 3680 2972 3732
rect 3024 3680 3039 3732
rect 3091 3680 3106 3732
rect 3158 3680 3173 3732
rect 3225 3680 3240 3732
rect 3292 3680 3307 3732
rect 3359 3680 3374 3732
rect 3426 3680 3441 3732
rect 3493 3680 3508 3732
rect 3560 3680 3575 3732
rect 3627 3680 3642 3732
rect 3694 3680 3708 3732
rect 3760 3680 3774 3732
rect 3826 3680 3832 3732
rect 2765 3664 3832 3680
rect 2765 3612 2771 3664
rect 2823 3612 2838 3664
rect 2890 3612 2905 3664
rect 2957 3612 2972 3664
rect 3024 3612 3039 3664
rect 3091 3612 3106 3664
rect 3158 3612 3173 3664
rect 3225 3612 3240 3664
rect 3292 3612 3307 3664
rect 3359 3612 3374 3664
rect 3426 3612 3441 3664
rect 3493 3612 3508 3664
rect 3560 3612 3575 3664
rect 3627 3612 3642 3664
rect 3694 3612 3708 3664
rect 3760 3612 3774 3664
rect 3826 3612 3832 3664
rect 2765 3596 3832 3612
rect 2765 3544 2771 3596
rect 2823 3544 2838 3596
rect 2890 3544 2905 3596
rect 2957 3544 2972 3596
rect 3024 3544 3039 3596
rect 3091 3544 3106 3596
rect 3158 3544 3173 3596
rect 3225 3544 3240 3596
rect 3292 3544 3307 3596
rect 3359 3544 3374 3596
rect 3426 3544 3441 3596
rect 3493 3544 3508 3596
rect 3560 3544 3575 3596
rect 3627 3544 3642 3596
rect 3694 3544 3708 3596
rect 3760 3544 3774 3596
rect 3826 3544 3832 3596
rect 2765 3528 3832 3544
rect 2765 3476 2771 3528
rect 2823 3476 2838 3528
rect 2890 3476 2905 3528
rect 2957 3476 2972 3528
rect 3024 3476 3039 3528
rect 3091 3476 3106 3528
rect 3158 3476 3173 3528
rect 3225 3476 3240 3528
rect 3292 3476 3307 3528
rect 3359 3476 3374 3528
rect 3426 3476 3441 3528
rect 3493 3476 3508 3528
rect 3560 3476 3575 3528
rect 3627 3476 3642 3528
rect 3694 3476 3708 3528
rect 3760 3476 3774 3528
rect 3826 3476 3832 3528
rect 2765 3470 3832 3476
rect 13947 3988 13953 4022
rect 13987 3988 14091 4022
rect 14125 3988 14131 4022
rect 13947 3947 14131 3988
rect 13947 3913 13953 3947
rect 13987 3913 14091 3947
rect 14125 3913 14131 3947
rect 13947 3872 14131 3913
rect 13947 3838 13953 3872
rect 13987 3838 14091 3872
rect 14125 3838 14131 3872
rect 13947 3797 14131 3838
rect 13947 3763 13953 3797
rect 13987 3763 14091 3797
rect 14125 3763 14131 3797
rect 13947 3722 14131 3763
rect 13947 3688 13953 3722
rect 13987 3688 14091 3722
rect 14125 3688 14131 3722
rect 13947 3647 14131 3688
rect 13947 3613 13953 3647
rect 13987 3613 14091 3647
rect 14125 3613 14131 3647
rect 13947 3571 14131 3613
rect 13947 3537 13953 3571
rect 13987 3537 14091 3571
rect 14125 3537 14131 3571
rect 13947 3495 14131 3537
rect 2436 3447 2514 3448
rect 2324 3409 2514 3447
rect 2324 3408 2474 3409
rect 2324 3374 2330 3408
rect 2364 3374 2402 3408
rect 2436 3375 2474 3408
rect 2508 3375 2514 3409
rect 2436 3374 2514 3375
rect 2324 3336 2514 3374
rect 2324 3335 2474 3336
rect 2324 3301 2330 3335
rect 2364 3301 2402 3335
rect 2436 3302 2474 3335
rect 2508 3302 2514 3336
rect 2436 3301 2514 3302
rect 2324 3263 2514 3301
rect 2324 3262 2474 3263
rect 2324 3228 2330 3262
rect 2364 3228 2402 3262
rect 2436 3229 2474 3262
rect 2508 3229 2514 3263
rect 2436 3228 2514 3229
rect 2324 3190 2514 3228
rect 13947 3461 13953 3495
rect 13987 3461 14091 3495
rect 14125 3461 14131 3495
rect 13947 3419 14131 3461
rect 13947 3385 13953 3419
rect 13987 3385 14091 3419
rect 14125 3385 14131 3419
rect 13947 3343 14131 3385
rect 13947 3309 13953 3343
rect 13987 3309 14091 3343
rect 14125 3309 14131 3343
rect 13947 3267 14131 3309
rect 13947 3233 13953 3267
rect 13987 3233 14091 3267
rect 14125 3233 14131 3267
rect 13947 3221 14131 3233
rect 2324 3189 2474 3190
rect 2324 3155 2330 3189
rect 2364 3155 2402 3189
rect 2436 3156 2474 3189
rect 2508 3156 2514 3190
rect 2436 3155 2514 3156
rect 2324 3117 2514 3155
tri 14642 3152 14676 3186 se
rect 14676 3152 14724 4333
rect 2324 3116 2474 3117
rect 2324 3082 2330 3116
rect 2364 3082 2402 3116
rect 2436 3083 2474 3116
rect 2508 3083 2514 3117
rect 13716 3100 14724 3152
rect 2436 3082 2514 3083
rect 2324 3044 2514 3082
tri 14642 3066 14676 3100 ne
rect 2324 3043 2474 3044
rect 2324 3009 2330 3043
rect 2364 3009 2402 3043
rect 2436 3010 2474 3043
rect 2508 3010 2514 3044
rect 2436 3009 2514 3010
rect 2324 2971 2514 3009
rect 2324 2970 2474 2971
rect 2324 272 2330 2970
rect 2436 2937 2474 2970
rect 2508 2937 2514 2971
rect 2436 2898 2514 2937
rect 2508 472 2514 2898
rect 13947 2983 14131 2995
rect 13947 2949 13953 2983
rect 13987 2949 14091 2983
rect 14125 2949 14131 2983
rect 13947 2908 14131 2949
rect 13947 2874 13953 2908
rect 13987 2874 14091 2908
rect 14125 2874 14131 2908
rect 13947 2833 14131 2874
rect 13947 2799 13953 2833
rect 13987 2799 14091 2833
rect 14125 2799 14131 2833
rect 2760 2792 4879 2793
rect 2760 2740 2766 2792
rect 2818 2740 2831 2792
rect 2883 2740 2896 2792
rect 2948 2740 2961 2792
rect 3013 2740 3026 2792
rect 3078 2740 3091 2792
rect 3143 2740 3156 2792
rect 3208 2740 3221 2792
rect 3273 2740 3285 2792
rect 3337 2740 3349 2792
rect 3401 2740 3413 2792
rect 3465 2740 3477 2792
rect 3529 2740 3541 2792
rect 3593 2740 3605 2792
rect 3657 2740 3669 2792
rect 3721 2740 3733 2792
rect 3785 2740 3797 2792
rect 3849 2740 3861 2792
rect 3913 2740 3925 2792
rect 3977 2740 3989 2792
rect 4041 2740 4053 2792
rect 4105 2740 4117 2792
rect 4169 2740 4181 2792
rect 4233 2740 4245 2792
rect 4297 2740 4309 2792
rect 4361 2740 4373 2792
rect 4425 2740 4437 2792
rect 4489 2740 4501 2792
rect 4553 2740 4565 2792
rect 4617 2740 4629 2792
rect 4681 2740 4693 2792
rect 4745 2740 4757 2792
rect 4809 2740 4821 2792
rect 4873 2740 4879 2792
rect 2760 2726 4879 2740
rect 2760 2674 2766 2726
rect 2818 2674 2831 2726
rect 2883 2674 2896 2726
rect 2948 2674 2961 2726
rect 3013 2674 3026 2726
rect 3078 2674 3091 2726
rect 3143 2674 3156 2726
rect 3208 2674 3221 2726
rect 3273 2674 3285 2726
rect 3337 2674 3349 2726
rect 3401 2674 3413 2726
rect 3465 2674 3477 2726
rect 3529 2674 3541 2726
rect 3593 2674 3605 2726
rect 3657 2674 3669 2726
rect 3721 2674 3733 2726
rect 3785 2674 3797 2726
rect 3849 2674 3861 2726
rect 3913 2674 3925 2726
rect 3977 2674 3989 2726
rect 4041 2674 4053 2726
rect 4105 2674 4117 2726
rect 4169 2674 4181 2726
rect 4233 2674 4245 2726
rect 4297 2674 4309 2726
rect 4361 2674 4373 2726
rect 4425 2674 4437 2726
rect 4489 2674 4501 2726
rect 4553 2674 4565 2726
rect 4617 2674 4629 2726
rect 4681 2674 4693 2726
rect 4745 2674 4757 2726
rect 4809 2674 4821 2726
rect 4873 2674 4879 2726
rect 2760 2660 4879 2674
rect 2760 2608 2766 2660
rect 2818 2608 2831 2660
rect 2883 2608 2896 2660
rect 2948 2608 2961 2660
rect 3013 2608 3026 2660
rect 3078 2608 3091 2660
rect 3143 2608 3156 2660
rect 3208 2608 3221 2660
rect 3273 2608 3285 2660
rect 3337 2608 3349 2660
rect 3401 2608 3413 2660
rect 3465 2608 3477 2660
rect 3529 2608 3541 2660
rect 3593 2608 3605 2660
rect 3657 2608 3669 2660
rect 3721 2608 3733 2660
rect 3785 2608 3797 2660
rect 3849 2608 3861 2660
rect 3913 2608 3925 2660
rect 3977 2608 3989 2660
rect 4041 2608 4053 2660
rect 4105 2608 4117 2660
rect 4169 2608 4181 2660
rect 4233 2608 4245 2660
rect 4297 2608 4309 2660
rect 4361 2608 4373 2660
rect 4425 2608 4437 2660
rect 4489 2608 4501 2660
rect 4553 2608 4565 2660
rect 4617 2608 4629 2660
rect 4681 2608 4693 2660
rect 4745 2608 4757 2660
rect 4809 2608 4821 2660
rect 4873 2608 4879 2660
rect 2760 2594 4879 2608
rect 2760 2542 2766 2594
rect 2818 2542 2831 2594
rect 2883 2542 2896 2594
rect 2948 2542 2961 2594
rect 3013 2542 3026 2594
rect 3078 2542 3091 2594
rect 3143 2542 3156 2594
rect 3208 2542 3221 2594
rect 3273 2542 3285 2594
rect 3337 2542 3349 2594
rect 3401 2542 3413 2594
rect 3465 2542 3477 2594
rect 3529 2542 3541 2594
rect 3593 2542 3605 2594
rect 3657 2542 3669 2594
rect 3721 2542 3733 2594
rect 3785 2542 3797 2594
rect 3849 2542 3861 2594
rect 3913 2542 3925 2594
rect 3977 2542 3989 2594
rect 4041 2542 4053 2594
rect 4105 2542 4117 2594
rect 4169 2542 4181 2594
rect 4233 2542 4245 2594
rect 4297 2542 4309 2594
rect 4361 2542 4373 2594
rect 4425 2542 4437 2594
rect 4489 2542 4501 2594
rect 4553 2542 4565 2594
rect 4617 2542 4629 2594
rect 4681 2542 4693 2594
rect 4745 2542 4757 2594
rect 4809 2542 4821 2594
rect 4873 2542 4879 2594
rect 2760 2528 4879 2542
rect 2760 2476 2766 2528
rect 2818 2476 2831 2528
rect 2883 2476 2896 2528
rect 2948 2476 2961 2528
rect 3013 2476 3026 2528
rect 3078 2476 3091 2528
rect 3143 2476 3156 2528
rect 3208 2476 3221 2528
rect 3273 2476 3285 2528
rect 3337 2476 3349 2528
rect 3401 2476 3413 2528
rect 3465 2476 3477 2528
rect 3529 2476 3541 2528
rect 3593 2476 3605 2528
rect 3657 2476 3669 2528
rect 3721 2476 3733 2528
rect 3785 2476 3797 2528
rect 3849 2476 3861 2528
rect 3913 2476 3925 2528
rect 3977 2476 3989 2528
rect 4041 2476 4053 2528
rect 4105 2476 4117 2528
rect 4169 2476 4181 2528
rect 4233 2476 4245 2528
rect 4297 2476 4309 2528
rect 4361 2476 4373 2528
rect 4425 2476 4437 2528
rect 4489 2476 4501 2528
rect 4553 2476 4565 2528
rect 4617 2476 4629 2528
rect 4681 2476 4693 2528
rect 4745 2476 4757 2528
rect 4809 2476 4821 2528
rect 4873 2476 4879 2528
rect 2760 2462 4879 2476
rect 2760 2410 2766 2462
rect 2818 2410 2831 2462
rect 2883 2410 2896 2462
rect 2948 2410 2961 2462
rect 3013 2410 3026 2462
rect 3078 2410 3091 2462
rect 3143 2410 3156 2462
rect 3208 2410 3221 2462
rect 3273 2410 3285 2462
rect 3337 2410 3349 2462
rect 3401 2410 3413 2462
rect 3465 2410 3477 2462
rect 3529 2410 3541 2462
rect 3593 2410 3605 2462
rect 3657 2410 3669 2462
rect 3721 2410 3733 2462
rect 3785 2410 3797 2462
rect 3849 2410 3861 2462
rect 3913 2410 3925 2462
rect 3977 2410 3989 2462
rect 4041 2410 4053 2462
rect 4105 2410 4117 2462
rect 4169 2410 4181 2462
rect 4233 2410 4245 2462
rect 4297 2410 4309 2462
rect 4361 2410 4373 2462
rect 4425 2410 4437 2462
rect 4489 2410 4501 2462
rect 4553 2410 4565 2462
rect 4617 2410 4629 2462
rect 4681 2410 4693 2462
rect 4745 2410 4757 2462
rect 4809 2410 4821 2462
rect 4873 2410 4879 2462
rect 2760 2396 4879 2410
rect 2760 2344 2766 2396
rect 2818 2344 2831 2396
rect 2883 2344 2896 2396
rect 2948 2344 2961 2396
rect 3013 2344 3026 2396
rect 3078 2344 3091 2396
rect 3143 2344 3156 2396
rect 3208 2344 3221 2396
rect 3273 2344 3285 2396
rect 3337 2344 3349 2396
rect 3401 2344 3413 2396
rect 3465 2344 3477 2396
rect 3529 2344 3541 2396
rect 3593 2344 3605 2396
rect 3657 2344 3669 2396
rect 3721 2344 3733 2396
rect 3785 2344 3797 2396
rect 3849 2344 3861 2396
rect 3913 2344 3925 2396
rect 3977 2344 3989 2396
rect 4041 2344 4053 2396
rect 4105 2344 4117 2396
rect 4169 2344 4181 2396
rect 4233 2344 4245 2396
rect 4297 2344 4309 2396
rect 4361 2344 4373 2396
rect 4425 2344 4437 2396
rect 4489 2344 4501 2396
rect 4553 2344 4565 2396
rect 4617 2344 4629 2396
rect 4681 2344 4693 2396
rect 4745 2344 4757 2396
rect 4809 2344 4821 2396
rect 4873 2344 4879 2396
rect 2760 2330 4879 2344
rect 2760 2278 2766 2330
rect 2818 2278 2831 2330
rect 2883 2278 2896 2330
rect 2948 2278 2961 2330
rect 3013 2278 3026 2330
rect 3078 2278 3091 2330
rect 3143 2278 3156 2330
rect 3208 2278 3221 2330
rect 3273 2278 3285 2330
rect 3337 2278 3349 2330
rect 3401 2278 3413 2330
rect 3465 2278 3477 2330
rect 3529 2278 3541 2330
rect 3593 2278 3605 2330
rect 3657 2278 3669 2330
rect 3721 2278 3733 2330
rect 3785 2278 3797 2330
rect 3849 2278 3861 2330
rect 3913 2278 3925 2330
rect 3977 2278 3989 2330
rect 4041 2278 4053 2330
rect 4105 2278 4117 2330
rect 4169 2278 4181 2330
rect 4233 2278 4245 2330
rect 4297 2278 4309 2330
rect 4361 2278 4373 2330
rect 4425 2278 4437 2330
rect 4489 2278 4501 2330
rect 4553 2278 4565 2330
rect 4617 2278 4629 2330
rect 4681 2278 4693 2330
rect 4745 2278 4757 2330
rect 4809 2278 4821 2330
rect 4873 2278 4879 2330
rect 2760 2264 4879 2278
rect 2760 2212 2766 2264
rect 2818 2212 2831 2264
rect 2883 2212 2896 2264
rect 2948 2212 2961 2264
rect 3013 2212 3026 2264
rect 3078 2212 3091 2264
rect 3143 2212 3156 2264
rect 3208 2212 3221 2264
rect 3273 2212 3285 2264
rect 3337 2212 3349 2264
rect 3401 2212 3413 2264
rect 3465 2212 3477 2264
rect 3529 2212 3541 2264
rect 3593 2212 3605 2264
rect 3657 2212 3669 2264
rect 3721 2212 3733 2264
rect 3785 2212 3797 2264
rect 3849 2212 3861 2264
rect 3913 2212 3925 2264
rect 3977 2212 3989 2264
rect 4041 2212 4053 2264
rect 4105 2212 4117 2264
rect 4169 2212 4181 2264
rect 4233 2212 4245 2264
rect 4297 2212 4309 2264
rect 4361 2212 4373 2264
rect 4425 2212 4437 2264
rect 4489 2212 4501 2264
rect 4553 2212 4565 2264
rect 4617 2212 4629 2264
rect 4681 2212 4693 2264
rect 4745 2212 4757 2264
rect 4809 2212 4821 2264
rect 4873 2212 4879 2264
rect 2760 2211 4879 2212
rect 13947 2758 14131 2799
rect 13947 2724 13953 2758
rect 13987 2724 14091 2758
rect 14125 2724 14131 2758
rect 13947 2683 14131 2724
rect 13947 2649 13953 2683
rect 13987 2649 14091 2683
rect 14125 2649 14131 2683
rect 13947 2608 14131 2649
rect 13947 2574 13953 2608
rect 13987 2574 14091 2608
rect 14125 2574 14131 2608
rect 13947 2533 14131 2574
rect 13947 2499 13953 2533
rect 13987 2499 14091 2533
rect 14125 2499 14131 2533
rect 13947 2458 14131 2499
rect 13947 2424 13953 2458
rect 13987 2424 14091 2458
rect 14125 2424 14131 2458
rect 13947 2383 14131 2424
rect 13947 2349 13953 2383
rect 13987 2349 14091 2383
rect 14125 2349 14131 2383
rect 13947 2307 14131 2349
rect 13947 2273 13953 2307
rect 13987 2273 14091 2307
rect 14125 2273 14131 2307
rect 13947 2231 14131 2273
rect 13947 2197 13953 2231
rect 13987 2197 14091 2231
rect 14125 2197 14131 2231
rect 13947 2155 14131 2197
rect 13947 2121 13953 2155
rect 13987 2121 14091 2155
rect 14125 2121 14131 2155
rect 13947 2079 14131 2121
rect 13947 2045 13953 2079
rect 13987 2045 14091 2079
rect 14125 2045 14131 2079
rect 13947 2003 14131 2045
rect 13947 1969 13953 2003
rect 13987 1969 14091 2003
rect 14125 1969 14131 2003
rect 13947 1957 14131 1969
tri 14642 1908 14676 1942 se
rect 14676 1908 14724 3100
rect 13716 1856 14724 1908
tri 14642 1822 14676 1856 ne
rect 13947 1783 14131 1795
rect 13947 1749 13953 1783
rect 13987 1749 14091 1783
rect 14125 1749 14131 1783
rect 13947 1708 14131 1749
rect 13947 1674 13953 1708
rect 13987 1674 14091 1708
rect 14125 1674 14131 1708
rect 13947 1633 14131 1674
rect 13947 1599 13953 1633
rect 13987 1599 14091 1633
rect 14125 1599 14131 1633
rect 13947 1558 14131 1599
rect 13947 1524 13953 1558
rect 13987 1524 14091 1558
rect 14125 1524 14131 1558
rect 2770 1513 4879 1519
rect 2770 1461 2776 1513
rect 2828 1461 2842 1513
rect 2894 1461 2908 1513
rect 2960 1461 2974 1513
rect 3026 1461 3040 1513
rect 3092 1461 3106 1513
rect 3158 1461 3172 1513
rect 3224 1461 3238 1513
rect 3290 1461 3304 1513
rect 3356 1461 3370 1513
rect 3422 1461 3436 1513
rect 3488 1461 3502 1513
rect 3554 1461 3568 1513
rect 3620 1461 3634 1513
rect 3686 1461 3700 1513
rect 3752 1461 3766 1513
rect 3818 1461 3832 1513
rect 3884 1461 3898 1513
rect 3950 1461 3964 1513
rect 4016 1461 4030 1513
rect 4082 1461 4096 1513
rect 4148 1461 4162 1513
rect 4214 1461 4228 1513
rect 4280 1461 4294 1513
rect 4346 1461 4360 1513
rect 4412 1461 4426 1513
rect 4478 1461 4492 1513
rect 4544 1461 4558 1513
rect 4610 1461 4624 1513
rect 4676 1461 4690 1513
rect 4742 1461 4756 1513
rect 4808 1461 4821 1513
rect 4873 1461 4879 1513
rect 2770 1445 4879 1461
rect 2770 1393 2776 1445
rect 2828 1393 2842 1445
rect 2894 1393 2908 1445
rect 2960 1393 2974 1445
rect 3026 1393 3040 1445
rect 3092 1393 3106 1445
rect 3158 1393 3172 1445
rect 3224 1393 3238 1445
rect 3290 1393 3304 1445
rect 3356 1393 3370 1445
rect 3422 1393 3436 1445
rect 3488 1393 3502 1445
rect 3554 1393 3568 1445
rect 3620 1393 3634 1445
rect 3686 1393 3700 1445
rect 3752 1393 3766 1445
rect 3818 1393 3832 1445
rect 3884 1393 3898 1445
rect 3950 1393 3964 1445
rect 4016 1393 4030 1445
rect 4082 1393 4096 1445
rect 4148 1393 4162 1445
rect 4214 1393 4228 1445
rect 4280 1393 4294 1445
rect 4346 1393 4360 1445
rect 4412 1393 4426 1445
rect 4478 1393 4492 1445
rect 4544 1393 4558 1445
rect 4610 1393 4624 1445
rect 4676 1393 4690 1445
rect 4742 1393 4756 1445
rect 4808 1393 4821 1445
rect 4873 1393 4879 1445
rect 2770 1377 4879 1393
rect 2770 1325 2776 1377
rect 2828 1325 2842 1377
rect 2894 1325 2908 1377
rect 2960 1325 2974 1377
rect 3026 1325 3040 1377
rect 3092 1325 3106 1377
rect 3158 1325 3172 1377
rect 3224 1325 3238 1377
rect 3290 1325 3304 1377
rect 3356 1325 3370 1377
rect 3422 1325 3436 1377
rect 3488 1325 3502 1377
rect 3554 1325 3568 1377
rect 3620 1325 3634 1377
rect 3686 1325 3700 1377
rect 3752 1325 3766 1377
rect 3818 1325 3832 1377
rect 3884 1325 3898 1377
rect 3950 1325 3964 1377
rect 4016 1325 4030 1377
rect 4082 1325 4096 1377
rect 4148 1325 4162 1377
rect 4214 1325 4228 1377
rect 4280 1325 4294 1377
rect 4346 1325 4360 1377
rect 4412 1325 4426 1377
rect 4478 1325 4492 1377
rect 4544 1325 4558 1377
rect 4610 1325 4624 1377
rect 4676 1325 4690 1377
rect 4742 1325 4756 1377
rect 4808 1325 4821 1377
rect 4873 1325 4879 1377
rect 2770 1309 4879 1325
rect 2770 1257 2776 1309
rect 2828 1257 2842 1309
rect 2894 1257 2908 1309
rect 2960 1257 2974 1309
rect 3026 1257 3040 1309
rect 3092 1257 3106 1309
rect 3158 1257 3172 1309
rect 3224 1257 3238 1309
rect 3290 1257 3304 1309
rect 3356 1257 3370 1309
rect 3422 1257 3436 1309
rect 3488 1257 3502 1309
rect 3554 1257 3568 1309
rect 3620 1257 3634 1309
rect 3686 1257 3700 1309
rect 3752 1257 3766 1309
rect 3818 1257 3832 1309
rect 3884 1257 3898 1309
rect 3950 1257 3964 1309
rect 4016 1257 4030 1309
rect 4082 1257 4096 1309
rect 4148 1257 4162 1309
rect 4214 1257 4228 1309
rect 4280 1257 4294 1309
rect 4346 1257 4360 1309
rect 4412 1257 4426 1309
rect 4478 1257 4492 1309
rect 4544 1257 4558 1309
rect 4610 1257 4624 1309
rect 4676 1257 4690 1309
rect 4742 1257 4756 1309
rect 4808 1257 4821 1309
rect 4873 1257 4879 1309
rect 2770 1241 4879 1257
rect 2770 1189 2776 1241
rect 2828 1189 2842 1241
rect 2894 1189 2908 1241
rect 2960 1189 2974 1241
rect 3026 1189 3040 1241
rect 3092 1189 3106 1241
rect 3158 1189 3172 1241
rect 3224 1189 3238 1241
rect 3290 1189 3304 1241
rect 3356 1189 3370 1241
rect 3422 1189 3436 1241
rect 3488 1189 3502 1241
rect 3554 1189 3568 1241
rect 3620 1189 3634 1241
rect 3686 1189 3700 1241
rect 3752 1189 3766 1241
rect 3818 1189 3832 1241
rect 3884 1189 3898 1241
rect 3950 1189 3964 1241
rect 4016 1189 4030 1241
rect 4082 1189 4096 1241
rect 4148 1189 4162 1241
rect 4214 1189 4228 1241
rect 4280 1189 4294 1241
rect 4346 1189 4360 1241
rect 4412 1189 4426 1241
rect 4478 1189 4492 1241
rect 4544 1189 4558 1241
rect 4610 1189 4624 1241
rect 4676 1189 4690 1241
rect 4742 1189 4756 1241
rect 4808 1189 4821 1241
rect 4873 1189 4879 1241
rect 2770 1173 4879 1189
rect 2770 1121 2776 1173
rect 2828 1121 2842 1173
rect 2894 1121 2908 1173
rect 2960 1121 2974 1173
rect 3026 1121 3040 1173
rect 3092 1121 3106 1173
rect 3158 1121 3172 1173
rect 3224 1121 3238 1173
rect 3290 1121 3304 1173
rect 3356 1121 3370 1173
rect 3422 1121 3436 1173
rect 3488 1121 3502 1173
rect 3554 1121 3568 1173
rect 3620 1121 3634 1173
rect 3686 1121 3700 1173
rect 3752 1121 3766 1173
rect 3818 1121 3832 1173
rect 3884 1121 3898 1173
rect 3950 1121 3964 1173
rect 4016 1121 4030 1173
rect 4082 1121 4096 1173
rect 4148 1121 4162 1173
rect 4214 1121 4228 1173
rect 4280 1121 4294 1173
rect 4346 1121 4360 1173
rect 4412 1121 4426 1173
rect 4478 1121 4492 1173
rect 4544 1121 4558 1173
rect 4610 1121 4624 1173
rect 4676 1121 4690 1173
rect 4742 1121 4756 1173
rect 4808 1121 4821 1173
rect 4873 1121 4879 1173
rect 2770 1105 4879 1121
rect 13947 1483 14131 1524
rect 13947 1449 13953 1483
rect 13987 1449 14091 1483
rect 14125 1449 14131 1483
rect 13947 1408 14131 1449
rect 13947 1374 13953 1408
rect 13987 1374 14091 1408
rect 14125 1374 14131 1408
rect 13947 1333 14131 1374
rect 13947 1299 13953 1333
rect 13987 1299 14091 1333
rect 14125 1299 14131 1333
rect 13947 1258 14131 1299
rect 13947 1224 13953 1258
rect 13987 1224 14091 1258
rect 14125 1224 14131 1258
rect 13947 1183 14131 1224
rect 13947 1149 13953 1183
rect 13987 1149 14091 1183
rect 14125 1149 14131 1183
rect 2770 1053 2776 1105
rect 2828 1053 2842 1105
rect 2894 1053 2908 1105
rect 2960 1053 2974 1105
rect 3026 1053 3040 1105
rect 3092 1053 3106 1105
rect 3158 1053 3172 1105
rect 3224 1053 3238 1105
rect 3290 1053 3304 1105
rect 3356 1053 3370 1105
rect 3422 1053 3436 1105
rect 3488 1053 3502 1105
rect 3554 1053 3568 1105
rect 3620 1053 3634 1105
rect 3686 1053 3700 1105
rect 3752 1053 3766 1105
rect 3818 1053 3832 1105
rect 3884 1053 3898 1105
rect 3950 1053 3964 1105
rect 4016 1053 4030 1105
rect 4082 1053 4096 1105
rect 4148 1053 4162 1105
rect 4214 1053 4228 1105
rect 4280 1053 4294 1105
rect 4346 1053 4360 1105
rect 4412 1053 4426 1105
rect 4478 1053 4492 1105
rect 4544 1053 4558 1105
rect 4610 1053 4624 1105
rect 4676 1053 4690 1105
rect 4742 1053 4756 1105
rect 4808 1053 4821 1105
rect 4873 1053 4879 1105
rect 2770 1037 4879 1053
rect 2770 985 2776 1037
rect 2828 985 2842 1037
rect 2894 985 2908 1037
rect 2960 985 2974 1037
rect 3026 985 3040 1037
rect 3092 985 3106 1037
rect 3158 985 3172 1037
rect 3224 985 3238 1037
rect 3290 985 3304 1037
rect 3356 985 3370 1037
rect 3422 985 3436 1037
rect 3488 985 3502 1037
rect 3554 985 3568 1037
rect 3620 985 3634 1037
rect 3686 985 3700 1037
rect 3752 985 3766 1037
rect 3818 985 3832 1037
rect 3884 985 3898 1037
rect 3950 985 3964 1037
rect 4016 985 4030 1037
rect 4082 985 4096 1037
rect 4148 985 4162 1037
rect 4214 985 4228 1037
rect 4280 985 4294 1037
rect 4346 985 4360 1037
rect 4412 985 4426 1037
rect 4478 985 4492 1037
rect 4544 985 4558 1037
rect 4610 985 4624 1037
rect 4676 985 4690 1037
rect 4742 985 4756 1037
rect 4808 985 4821 1037
rect 4873 985 4879 1037
rect 2770 979 4879 985
rect 6749 1106 6801 1112
rect 6749 1022 6801 1054
rect 6749 964 6801 970
rect 8703 1106 8755 1112
rect 8703 1022 8755 1054
rect 8703 964 8755 970
rect 13947 1107 14131 1149
rect 13947 1073 13953 1107
rect 13987 1073 14091 1107
rect 14125 1073 14131 1107
rect 13947 1031 14131 1073
rect 13947 997 13953 1031
rect 13987 997 14091 1031
rect 14125 997 14131 1031
rect 13947 955 14131 997
rect 13947 921 13953 955
rect 13987 921 14091 955
rect 14125 921 14131 955
rect 13947 879 14131 921
rect 13947 845 13953 879
rect 13987 845 14091 879
rect 14125 845 14131 879
rect 13947 803 14131 845
rect 13947 769 13953 803
rect 13987 769 14091 803
rect 14125 769 14131 803
rect 13947 757 14131 769
tri 14642 664 14676 698 se
rect 14676 664 14724 1856
rect 13716 612 14724 664
tri 14642 578 14676 612 ne
rect 14676 578 14724 612
rect 6701 521 6707 567
tri 6695 520 6696 521 ne
rect 6696 520 6707 521
tri 6696 515 6701 520 ne
rect 6701 515 6707 520
rect 6759 515 6791 567
rect 6843 521 6849 567
rect 8655 521 8661 567
rect 6843 520 6854 521
tri 6854 520 6855 521 nw
tri 8649 520 8650 521 ne
rect 8650 520 8661 521
rect 6843 515 6849 520
tri 6849 515 6854 520 nw
tri 8650 515 8655 520 ne
rect 8655 515 8661 520
rect 8713 515 8745 567
rect 8797 521 8803 567
rect 13946 554 14136 566
rect 8797 520 8808 521
tri 8808 520 8809 521 nw
rect 13946 520 13952 554
rect 13986 520 14024 554
rect 14058 520 14096 554
rect 14130 520 14136 554
rect 8797 515 8803 520
tri 8803 515 8808 520 nw
tri 2514 472 2522 480 sw
rect 13946 472 14136 520
rect 2508 466 2522 472
tri 2522 466 2528 472 sw
rect 13946 466 14024 472
rect 2508 432 2528 466
tri 2528 432 2562 466 sw
tri 13933 432 13946 445 se
rect 13946 432 13952 466
rect 13986 438 14024 466
rect 14058 438 14096 472
rect 14130 438 14136 472
rect 13986 432 14136 438
rect 2508 389 2562 432
tri 2562 389 2605 432 sw
tri 13890 389 13933 432 se
rect 13933 389 14136 432
rect 2508 384 2605 389
tri 2605 384 2610 389 sw
tri 13885 384 13890 389 se
rect 13890 384 14024 389
rect 2508 378 14024 384
rect 2508 344 2547 378
rect 2581 344 2620 378
rect 2654 344 2693 378
rect 2727 344 2766 378
rect 2800 344 2839 378
rect 2873 344 2912 378
rect 2946 344 2985 378
rect 3019 344 3058 378
rect 3092 344 3131 378
rect 3165 344 3204 378
rect 3238 344 3277 378
rect 3311 344 3350 378
rect 3384 344 3423 378
rect 3457 344 3496 378
rect 3530 344 3569 378
rect 3603 344 3642 378
rect 3676 344 3715 378
rect 3749 344 3788 378
rect 3822 344 3861 378
rect 3895 344 3934 378
rect 3968 344 4007 378
rect 4041 344 4080 378
rect 4114 344 4153 378
rect 4187 344 4226 378
rect 4260 344 4299 378
rect 4333 344 4372 378
rect 4406 344 4445 378
rect 4479 344 4518 378
rect 4552 344 4591 378
rect 4625 344 4664 378
rect 2436 306 4664 344
rect 13986 355 14024 378
rect 14058 355 14096 389
rect 14130 355 14136 389
rect 2436 272 2475 306
rect 2509 272 2548 306
rect 2582 272 2621 306
rect 2655 272 2694 306
rect 2728 272 2767 306
rect 2801 272 2840 306
rect 2874 272 2913 306
rect 2947 272 2986 306
rect 3020 272 3059 306
rect 3093 272 3132 306
rect 3166 272 3205 306
rect 3239 272 3278 306
rect 3312 272 3351 306
rect 3385 272 3424 306
rect 3458 272 3497 306
rect 3531 272 3570 306
rect 3604 272 3643 306
rect 3677 272 3716 306
rect 3750 272 3789 306
rect 3823 272 3862 306
rect 3896 272 3935 306
rect 3969 272 4008 306
rect 4042 272 4081 306
rect 4115 272 4154 306
rect 4188 272 4227 306
rect 4261 272 4300 306
rect 4334 272 4373 306
rect 4407 272 4446 306
rect 4480 272 4519 306
rect 4553 272 4592 306
rect 2324 234 4592 272
rect 13986 306 14136 355
rect 14058 272 14096 306
rect 14130 272 14136 306
rect 2324 200 2402 234
rect 2436 200 2475 234
rect 2509 200 2548 234
rect 2582 200 2621 234
rect 2655 200 2694 234
rect 2728 200 2767 234
rect 2801 200 2840 234
rect 2874 200 2913 234
rect 2947 200 2986 234
rect 3020 200 3059 234
rect 3093 200 3132 234
rect 3166 200 3205 234
rect 3239 200 3278 234
rect 3312 200 3351 234
rect 3385 200 3424 234
rect 3458 200 3497 234
rect 3531 200 3570 234
rect 3604 200 3643 234
rect 3677 200 3716 234
rect 3750 200 3789 234
rect 3823 200 3862 234
rect 3896 200 3935 234
rect 3969 200 4008 234
rect 4042 200 4081 234
rect 4115 200 4154 234
rect 4188 200 4227 234
rect 4261 200 4300 234
rect 4334 200 4373 234
rect 4407 200 4446 234
rect 4480 200 4519 234
rect 4553 200 4592 234
rect 14058 200 14136 272
rect 2324 197 5190 200
rect 5242 197 5256 200
rect 5308 197 5322 200
rect 5374 197 5388 200
rect 5440 197 5453 200
rect 5505 197 5518 200
rect 5570 197 14136 200
rect 2324 194 14136 197
<< via1 >>
rect 2231 37941 2283 37993
rect 2335 37941 2387 37993
rect 2231 37877 2283 37929
rect 2335 37877 2387 37929
rect 2231 37855 2283 37865
rect 2335 37855 2387 37865
rect 2231 37816 2283 37855
rect 2335 37816 2387 37855
rect 2231 37813 2254 37816
rect 2254 37813 2283 37816
rect 2231 37782 2254 37801
rect 2254 37782 2283 37801
rect 2335 37813 2364 37816
rect 2364 37813 2387 37816
rect 2335 37782 2364 37801
rect 2364 37782 2387 37801
rect 2231 37749 2283 37782
rect 2335 37749 2387 37782
rect 2231 37709 2254 37737
rect 2254 37709 2283 37737
rect 2335 37709 2364 37737
rect 2364 37709 2387 37737
rect 2231 37685 2283 37709
rect 2335 37685 2387 37709
rect 2231 37670 2283 37673
rect 2335 37670 2387 37673
rect 2231 37636 2254 37670
rect 2254 37636 2283 37670
rect 2335 37636 2364 37670
rect 2364 37636 2387 37670
rect 2231 37621 2283 37636
rect 2335 37621 2387 37636
rect 2231 37597 2283 37609
rect 2335 37597 2387 37609
rect 2231 37563 2254 37597
rect 2254 37563 2283 37597
rect 2335 37563 2364 37597
rect 2364 37563 2387 37597
rect 2231 37557 2283 37563
rect 2335 37557 2387 37563
rect 2231 37524 2283 37545
rect 2335 37524 2387 37545
rect 2231 37493 2254 37524
rect 2254 37493 2283 37524
rect 2335 37493 2364 37524
rect 2364 37493 2387 37524
rect 2231 37451 2283 37481
rect 2335 37451 2387 37481
rect 2231 37429 2254 37451
rect 2254 37429 2283 37451
rect 2335 37429 2364 37451
rect 2364 37429 2387 37451
rect 2231 37378 2283 37417
rect 2335 37378 2387 37417
rect 2231 37365 2254 37378
rect 2254 37365 2283 37378
rect 2231 37344 2254 37353
rect 2254 37344 2283 37353
rect 2335 37365 2364 37378
rect 2364 37365 2387 37378
rect 2335 37344 2364 37353
rect 2364 37344 2387 37353
rect 2231 37305 2283 37344
rect 2335 37305 2387 37344
rect 2231 37301 2254 37305
rect 2254 37301 2283 37305
rect 2231 37271 2254 37289
rect 2254 37271 2283 37289
rect 2335 37301 2364 37305
rect 2364 37301 2387 37305
rect 2335 37271 2364 37289
rect 2364 37271 2387 37289
rect 2231 37237 2283 37271
rect 2335 37237 2387 37271
rect 2231 37198 2254 37225
rect 2254 37198 2283 37225
rect 2335 37198 2364 37225
rect 2364 37198 2387 37225
rect 2231 37173 2283 37198
rect 2335 37173 2387 37198
rect 2231 37159 2283 37161
rect 2335 37159 2387 37161
rect 2231 37125 2254 37159
rect 2254 37125 2283 37159
rect 2335 37125 2364 37159
rect 2364 37125 2387 37159
rect 2231 37109 2283 37125
rect 2335 37109 2387 37125
rect 2231 37086 2283 37097
rect 2335 37086 2387 37097
rect 2231 37052 2254 37086
rect 2254 37052 2283 37086
rect 2335 37052 2364 37086
rect 2364 37052 2387 37086
rect 2231 37045 2283 37052
rect 2335 37045 2387 37052
rect 2231 37013 2283 37033
rect 2335 37013 2387 37033
rect 2231 36981 2254 37013
rect 2254 36981 2283 37013
rect 2335 36981 2364 37013
rect 2364 36981 2387 37013
rect 2231 36940 2283 36969
rect 2335 36940 2387 36969
rect 2231 36917 2254 36940
rect 2254 36917 2283 36940
rect 2335 36917 2364 36940
rect 2364 36917 2387 36940
rect 2231 36867 2283 36905
rect 2335 36867 2387 36905
rect 2231 36853 2254 36867
rect 2254 36853 2283 36867
rect 2231 36833 2254 36841
rect 2254 36833 2283 36841
rect 2335 36853 2364 36867
rect 2364 36853 2387 36867
rect 2335 36833 2364 36841
rect 2364 36833 2387 36841
rect 2231 36794 2283 36833
rect 2335 36794 2387 36833
rect 2231 36789 2254 36794
rect 2254 36789 2283 36794
rect 2231 36760 2254 36777
rect 2254 36760 2283 36777
rect 2335 36789 2364 36794
rect 2364 36789 2387 36794
rect 2335 36760 2364 36777
rect 2364 36760 2387 36777
rect 2231 36725 2283 36760
rect 2335 36725 2387 36760
rect 2231 36687 2254 36713
rect 2254 36687 2283 36713
rect 2335 36687 2364 36713
rect 2364 36687 2387 36713
rect 2231 36661 2283 36687
rect 2335 36661 2387 36687
rect 2231 36648 2283 36649
rect 2335 36648 2387 36649
rect 2231 36614 2254 36648
rect 2254 36614 2283 36648
rect 2335 36614 2364 36648
rect 2364 36614 2387 36648
rect 2231 36597 2283 36614
rect 2335 36597 2387 36614
rect 2231 36575 2283 36585
rect 2335 36575 2387 36585
rect 2231 36541 2254 36575
rect 2254 36541 2283 36575
rect 2335 36541 2364 36575
rect 2364 36541 2387 36575
rect 2231 36533 2283 36541
rect 2335 36533 2387 36541
rect 2231 36502 2283 36521
rect 2335 36502 2387 36521
rect 2231 36469 2254 36502
rect 2254 36469 2283 36502
rect 2335 36469 2364 36502
rect 2364 36469 2387 36502
rect 2231 36429 2283 36457
rect 2335 36429 2387 36457
rect 2231 36405 2254 36429
rect 2254 36405 2283 36429
rect 2335 36405 2364 36429
rect 2364 36405 2387 36429
rect 2231 36356 2283 36393
rect 2335 36356 2387 36393
rect 2231 36341 2254 36356
rect 2254 36341 2283 36356
rect 2231 36322 2254 36329
rect 2254 36322 2283 36329
rect 2335 36341 2364 36356
rect 2364 36341 2387 36356
rect 2335 36322 2364 36329
rect 2364 36322 2387 36329
rect 2231 36283 2283 36322
rect 2335 36283 2387 36322
rect 2231 36277 2254 36283
rect 2254 36277 2283 36283
rect 2231 36249 2254 36265
rect 2254 36249 2283 36265
rect 2335 36277 2364 36283
rect 2364 36277 2387 36283
rect 2335 36249 2364 36265
rect 2364 36249 2387 36265
rect 2231 36213 2283 36249
rect 2335 36213 2387 36249
rect 2231 36176 2254 36201
rect 2254 36176 2283 36201
rect 2335 36176 2364 36201
rect 2364 36176 2387 36201
rect 2231 36149 2283 36176
rect 2335 36149 2387 36176
rect 2231 36103 2254 36137
rect 2254 36103 2283 36137
rect 2335 36103 2364 36137
rect 2364 36103 2387 36137
rect 2231 36085 2283 36103
rect 2335 36085 2387 36103
rect 2231 36064 2283 36073
rect 2335 36064 2387 36073
rect 2231 36030 2254 36064
rect 2254 36030 2283 36064
rect 2335 36030 2364 36064
rect 2364 36030 2387 36064
rect 2231 36021 2283 36030
rect 2335 36021 2387 36030
rect 2231 35991 2283 36009
rect 2335 35991 2387 36009
rect 2231 35957 2254 35991
rect 2254 35957 2283 35991
rect 2335 35957 2364 35991
rect 2364 35957 2387 35991
rect 2231 35918 2283 35945
rect 2335 35918 2387 35945
rect 2231 35893 2254 35918
rect 2254 35893 2283 35918
rect 2335 35893 2364 35918
rect 2364 35893 2387 35918
rect 2231 35845 2283 35881
rect 2335 35845 2387 35881
rect 2231 35829 2254 35845
rect 2254 35829 2283 35845
rect 2231 35811 2254 35817
rect 2254 35811 2283 35817
rect 2335 35829 2364 35845
rect 2364 35829 2387 35845
rect 2335 35811 2364 35817
rect 2364 35811 2387 35817
rect 2231 35772 2283 35811
rect 2335 35772 2387 35811
rect 2231 35765 2254 35772
rect 2254 35765 2283 35772
rect 2231 35738 2254 35753
rect 2254 35738 2283 35753
rect 2335 35765 2364 35772
rect 2364 35765 2387 35772
rect 2335 35738 2364 35753
rect 2364 35738 2387 35753
rect 2231 35701 2283 35738
rect 2335 35701 2387 35738
rect 2231 35665 2254 35689
rect 2254 35665 2283 35689
rect 2335 35665 2364 35689
rect 2364 35665 2387 35689
rect 2231 35637 2283 35665
rect 2335 35637 2387 35665
rect 2231 35592 2254 35625
rect 2254 35592 2283 35625
rect 2335 35592 2364 35625
rect 2364 35592 2387 35625
rect 2231 35573 2283 35592
rect 2335 35573 2387 35592
rect 2231 35553 2283 35561
rect 2335 35553 2387 35561
rect 2231 35519 2254 35553
rect 2254 35519 2283 35553
rect 2335 35519 2364 35553
rect 2364 35519 2387 35553
rect 2231 35509 2283 35519
rect 2335 35509 2387 35519
rect 2231 35480 2283 35497
rect 2335 35480 2387 35497
rect 2231 35446 2254 35480
rect 2254 35446 2283 35480
rect 2335 35446 2364 35480
rect 2364 35446 2387 35480
rect 2231 35445 2283 35446
rect 2335 35445 2387 35446
rect 2231 35407 2283 35433
rect 2335 35407 2387 35433
rect 2231 35381 2254 35407
rect 2254 35381 2283 35407
rect 2335 35381 2364 35407
rect 2364 35381 2387 35407
rect 2231 35334 2283 35369
rect 2335 35334 2387 35369
rect 2231 35317 2254 35334
rect 2254 35317 2283 35334
rect 2231 35300 2254 35305
rect 2254 35300 2283 35305
rect 2335 35317 2364 35334
rect 2364 35317 2387 35334
rect 2335 35300 2364 35305
rect 2364 35300 2387 35305
rect 2231 35261 2283 35300
rect 2335 35261 2387 35300
rect 2231 35253 2254 35261
rect 2254 35253 2283 35261
rect 2231 35227 2254 35241
rect 2254 35227 2283 35241
rect 2335 35253 2364 35261
rect 2364 35253 2387 35261
rect 2335 35227 2364 35241
rect 2364 35227 2387 35241
rect 2231 35189 2283 35227
rect 2335 35189 2387 35227
rect 2231 35154 2254 35176
rect 2254 35154 2283 35176
rect 2335 35154 2364 35176
rect 2364 35154 2387 35176
rect 2231 35124 2283 35154
rect 2335 35124 2387 35154
rect 2231 35081 2254 35111
rect 2254 35081 2283 35111
rect 2335 35081 2364 35111
rect 2364 35081 2387 35111
rect 2231 35059 2283 35081
rect 2335 35059 2387 35081
rect 2231 35042 2283 35046
rect 2335 35042 2387 35046
rect 2231 35008 2254 35042
rect 2254 35008 2283 35042
rect 2335 35008 2364 35042
rect 2364 35008 2387 35042
rect 2231 34994 2283 35008
rect 2335 34994 2387 35008
rect 2231 34969 2283 34981
rect 2335 34969 2387 34981
rect 2231 34935 2254 34969
rect 2254 34935 2283 34969
rect 2335 34935 2364 34969
rect 2364 34935 2387 34969
rect 2231 34929 2283 34935
rect 2335 34929 2387 34935
rect 2231 34896 2283 34916
rect 2335 34896 2387 34916
rect 2231 34864 2254 34896
rect 2254 34864 2283 34896
rect 2335 34864 2364 34896
rect 2364 34864 2387 34896
rect 2231 34823 2283 34851
rect 2335 34823 2387 34851
rect 2231 34799 2254 34823
rect 2254 34799 2283 34823
rect 2335 34799 2364 34823
rect 2364 34799 2387 34823
rect 2231 34750 2283 34786
rect 2335 34750 2387 34786
rect 2231 34734 2254 34750
rect 2254 34734 2283 34750
rect 2231 34716 2254 34721
rect 2254 34716 2283 34721
rect 2335 34734 2364 34750
rect 2364 34734 2387 34750
rect 2335 34716 2364 34721
rect 2364 34716 2387 34721
rect 2231 34677 2283 34716
rect 2335 34677 2387 34716
rect 2231 34669 2254 34677
rect 2254 34669 2283 34677
rect 2231 34643 2254 34656
rect 2254 34643 2283 34656
rect 2335 34669 2364 34677
rect 2364 34669 2387 34677
rect 2335 34643 2364 34656
rect 2364 34643 2387 34656
rect 2231 34604 2283 34643
rect 2335 34604 2387 34643
rect 2231 34570 2254 34591
rect 2254 34570 2283 34591
rect 2335 34570 2364 34591
rect 2364 34570 2387 34591
rect 2231 34539 2283 34570
rect 2335 34539 2387 34570
rect 2231 34497 2254 34526
rect 2254 34497 2283 34526
rect 2335 34497 2364 34526
rect 2364 34497 2387 34526
rect 2231 34474 2283 34497
rect 2335 34474 2387 34497
rect 2231 34458 2283 34461
rect 2335 34458 2387 34461
rect 2231 34424 2254 34458
rect 2254 34424 2283 34458
rect 2335 34424 2364 34458
rect 2364 34424 2387 34458
rect 2231 34409 2283 34424
rect 2335 34409 2387 34424
rect 2231 34385 2283 34396
rect 2335 34385 2387 34396
rect 2231 34351 2254 34385
rect 2254 34351 2283 34385
rect 2335 34351 2364 34385
rect 2364 34351 2387 34385
rect 2231 34344 2283 34351
rect 2335 34344 2387 34351
rect 2231 34312 2283 34331
rect 2335 34312 2387 34331
rect 2231 34279 2254 34312
rect 2254 34279 2283 34312
rect 2335 34279 2364 34312
rect 2364 34279 2387 34312
rect 2231 34239 2283 34266
rect 2335 34239 2387 34266
rect 2231 34214 2254 34239
rect 2254 34214 2283 34239
rect 2335 34214 2364 34239
rect 2364 34214 2387 34239
rect 2872 38957 2877 39009
rect 2877 38957 2924 39009
rect 2940 38957 2992 39009
rect 3008 38957 3055 39009
rect 3055 38957 3060 39009
rect 2872 38892 2877 38944
rect 2877 38892 2924 38944
rect 2940 38892 2992 38944
rect 3008 38892 3055 38944
rect 3055 38892 3060 38944
rect 2872 38827 2877 38879
rect 2877 38827 2924 38879
rect 2940 38827 2992 38879
rect 3008 38827 3055 38879
rect 3055 38827 3060 38879
rect 2872 38762 2877 38814
rect 2877 38762 2924 38814
rect 2940 38762 2992 38814
rect 3008 38762 3055 38814
rect 3055 38762 3060 38814
rect 2872 38697 2877 38749
rect 2877 38697 2924 38749
rect 2940 38697 2992 38749
rect 3008 38697 3055 38749
rect 3055 38697 3060 38749
rect 2872 38632 2877 38684
rect 2877 38632 2924 38684
rect 2940 38632 2992 38684
rect 3008 38632 3055 38684
rect 3055 38632 3060 38684
rect 2872 38567 2877 38619
rect 2877 38567 2924 38619
rect 2940 38567 2992 38619
rect 3008 38567 3055 38619
rect 3055 38567 3060 38619
rect 2872 38502 2877 38554
rect 2877 38502 2924 38554
rect 2940 38502 2992 38554
rect 3008 38502 3055 38554
rect 3055 38502 3060 38554
rect 2872 38438 2877 38490
rect 2877 38438 2924 38490
rect 2940 38438 2992 38490
rect 3008 38438 3055 38490
rect 3055 38438 3060 38490
rect 2872 38374 2877 38426
rect 2877 38374 2924 38426
rect 2940 38374 2992 38426
rect 3008 38374 3055 38426
rect 3055 38374 3060 38426
rect 2872 38310 2877 38362
rect 2877 38310 2924 38362
rect 2940 38310 2992 38362
rect 3008 38310 3055 38362
rect 3055 38310 3060 38362
rect 2872 38246 2877 38298
rect 2877 38246 2924 38298
rect 2940 38246 2992 38298
rect 3008 38246 3055 38298
rect 3055 38246 3060 38298
rect 2872 38182 2877 38234
rect 2877 38182 2924 38234
rect 2940 38182 2992 38234
rect 3008 38182 3055 38234
rect 3055 38182 3060 38234
rect 2872 38118 2877 38170
rect 2877 38118 2924 38170
rect 2940 38118 2992 38170
rect 3008 38118 3055 38170
rect 3055 38118 3060 38170
rect 3792 38957 3797 39009
rect 3797 38957 3844 39009
rect 3860 38957 3912 39009
rect 3928 38957 3975 39009
rect 3975 38957 3980 39009
rect 3792 38892 3797 38944
rect 3797 38892 3844 38944
rect 3860 38892 3912 38944
rect 3928 38892 3975 38944
rect 3975 38892 3980 38944
rect 3792 38827 3797 38879
rect 3797 38827 3844 38879
rect 3860 38827 3912 38879
rect 3928 38827 3975 38879
rect 3975 38827 3980 38879
rect 3792 38762 3797 38814
rect 3797 38762 3844 38814
rect 3860 38762 3912 38814
rect 3928 38762 3975 38814
rect 3975 38762 3980 38814
rect 3792 38697 3797 38749
rect 3797 38697 3844 38749
rect 3860 38697 3912 38749
rect 3928 38697 3975 38749
rect 3975 38697 3980 38749
rect 3792 38632 3797 38684
rect 3797 38632 3844 38684
rect 3860 38632 3912 38684
rect 3928 38632 3975 38684
rect 3975 38632 3980 38684
rect 3792 38567 3797 38619
rect 3797 38567 3844 38619
rect 3860 38567 3912 38619
rect 3928 38567 3975 38619
rect 3975 38567 3980 38619
rect 3792 38502 3797 38554
rect 3797 38502 3844 38554
rect 3860 38502 3912 38554
rect 3928 38502 3975 38554
rect 3975 38502 3980 38554
rect 3792 38438 3797 38490
rect 3797 38438 3844 38490
rect 3860 38438 3912 38490
rect 3928 38438 3975 38490
rect 3975 38438 3980 38490
rect 3792 38374 3797 38426
rect 3797 38374 3844 38426
rect 3860 38374 3912 38426
rect 3928 38374 3975 38426
rect 3975 38374 3980 38426
rect 3792 38310 3797 38362
rect 3797 38310 3844 38362
rect 3860 38310 3912 38362
rect 3928 38310 3975 38362
rect 3975 38310 3980 38362
rect 3792 38246 3797 38298
rect 3797 38246 3844 38298
rect 3860 38246 3912 38298
rect 3928 38246 3975 38298
rect 3975 38246 3980 38298
rect 3792 38182 3797 38234
rect 3797 38182 3844 38234
rect 3860 38182 3912 38234
rect 3928 38182 3975 38234
rect 3975 38182 3980 38234
rect 3792 38118 3797 38170
rect 3797 38118 3844 38170
rect 3860 38118 3912 38170
rect 3928 38118 3975 38170
rect 3975 38118 3980 38170
rect 2872 36316 2924 36368
rect 2940 36362 2992 36368
rect 2940 36328 2943 36362
rect 2943 36328 2977 36362
rect 2977 36328 2992 36362
rect 2940 36316 2992 36328
rect 3008 36362 3060 36368
rect 3008 36328 3021 36362
rect 3021 36328 3055 36362
rect 3055 36328 3060 36362
rect 3008 36316 3060 36328
rect 2872 36252 2924 36304
rect 2940 36290 2992 36304
rect 2940 36256 2943 36290
rect 2943 36256 2977 36290
rect 2977 36256 2992 36290
rect 2940 36252 2992 36256
rect 3008 36290 3060 36304
rect 3008 36256 3021 36290
rect 3021 36256 3055 36290
rect 3055 36256 3060 36290
rect 3008 36252 3060 36256
rect 2872 36187 2924 36239
rect 2940 36218 2992 36239
rect 2940 36187 2943 36218
rect 2943 36187 2977 36218
rect 2977 36187 2992 36218
rect 3008 36218 3060 36239
rect 3008 36187 3021 36218
rect 3021 36187 3055 36218
rect 3055 36187 3060 36218
rect 2872 36122 2924 36174
rect 2940 36146 2992 36174
rect 2940 36122 2943 36146
rect 2943 36122 2977 36146
rect 2977 36122 2992 36146
rect 3008 36146 3060 36174
rect 3008 36122 3021 36146
rect 3021 36122 3055 36146
rect 3055 36122 3060 36146
rect 2872 36057 2924 36109
rect 2940 36074 2992 36109
rect 2940 36057 2943 36074
rect 2943 36057 2977 36074
rect 2977 36057 2992 36074
rect 3008 36074 3060 36109
rect 3008 36057 3021 36074
rect 3021 36057 3055 36074
rect 3055 36057 3060 36074
rect 2872 35992 2924 36044
rect 2940 36040 2943 36044
rect 2943 36040 2977 36044
rect 2977 36040 2992 36044
rect 2940 36002 2992 36040
rect 2940 35992 2943 36002
rect 2943 35992 2977 36002
rect 2977 35992 2992 36002
rect 3008 36040 3021 36044
rect 3021 36040 3055 36044
rect 3055 36040 3060 36044
rect 3008 36002 3060 36040
rect 3008 35992 3021 36002
rect 3021 35992 3055 36002
rect 3055 35992 3060 36002
rect 2872 35927 2924 35979
rect 2940 35968 2943 35979
rect 2943 35968 2977 35979
rect 2977 35968 2992 35979
rect 2940 35930 2992 35968
rect 2940 35927 2943 35930
rect 2943 35927 2977 35930
rect 2977 35927 2992 35930
rect 3008 35968 3021 35979
rect 3021 35968 3055 35979
rect 3055 35968 3060 35979
rect 3008 35930 3060 35968
rect 3008 35927 3021 35930
rect 3021 35927 3055 35930
rect 3055 35927 3060 35930
rect 2872 35862 2924 35914
rect 2940 35896 2943 35914
rect 2943 35896 2977 35914
rect 2977 35896 2992 35914
rect 2940 35862 2992 35896
rect 3008 35896 3021 35914
rect 3021 35896 3055 35914
rect 3055 35896 3060 35914
rect 3008 35862 3060 35896
rect 2872 35797 2924 35849
rect 2940 35824 2943 35849
rect 2943 35824 2977 35849
rect 2977 35824 2992 35849
rect 2940 35797 2992 35824
rect 3008 35824 3021 35849
rect 3021 35824 3055 35849
rect 3055 35824 3060 35849
rect 3008 35797 3060 35824
rect 2872 35732 2924 35784
rect 2940 35752 2943 35784
rect 2943 35752 2977 35784
rect 2977 35752 2992 35784
rect 2940 35732 2992 35752
rect 3008 35752 3021 35784
rect 3021 35752 3055 35784
rect 3055 35752 3060 35784
rect 3008 35732 3060 35752
rect 2872 35667 2924 35719
rect 2940 35714 2992 35719
rect 2940 35680 2943 35714
rect 2943 35680 2977 35714
rect 2977 35680 2992 35714
rect 2940 35667 2992 35680
rect 3008 35714 3060 35719
rect 3008 35680 3021 35714
rect 3021 35680 3055 35714
rect 3055 35680 3060 35714
rect 3008 35667 3060 35680
rect 2872 35602 2924 35654
rect 2940 35642 2992 35654
rect 2940 35608 2943 35642
rect 2943 35608 2977 35642
rect 2977 35608 2992 35642
rect 2940 35602 2992 35608
rect 3008 35642 3060 35654
rect 3008 35608 3021 35642
rect 3021 35608 3055 35642
rect 3055 35608 3060 35642
rect 3008 35602 3060 35608
rect 2872 35537 2924 35589
rect 2940 35570 2992 35589
rect 2940 35537 2943 35570
rect 2943 35537 2977 35570
rect 2977 35537 2992 35570
rect 3008 35570 3060 35589
rect 3008 35537 3021 35570
rect 3021 35537 3055 35570
rect 3055 35537 3060 35570
rect 2872 35472 2924 35524
rect 2940 35498 2992 35524
rect 2940 35472 2943 35498
rect 2943 35472 2977 35498
rect 2977 35472 2992 35498
rect 3008 35498 3060 35524
rect 3008 35472 3021 35498
rect 3021 35472 3055 35498
rect 3055 35472 3060 35498
rect 2872 35407 2924 35459
rect 2940 35426 2992 35459
rect 2940 35407 2943 35426
rect 2943 35407 2977 35426
rect 2977 35407 2992 35426
rect 3008 35426 3060 35459
rect 3008 35407 3021 35426
rect 3021 35407 3055 35426
rect 3055 35407 3060 35426
rect 2872 35342 2924 35394
rect 2940 35392 2943 35394
rect 2943 35392 2977 35394
rect 2977 35392 2992 35394
rect 2940 35354 2992 35392
rect 2940 35342 2943 35354
rect 2943 35342 2977 35354
rect 2977 35342 2992 35354
rect 3008 35392 3021 35394
rect 3021 35392 3055 35394
rect 3055 35392 3060 35394
rect 3008 35354 3060 35392
rect 3008 35342 3021 35354
rect 3021 35342 3055 35354
rect 3055 35342 3060 35354
rect 2872 35277 2924 35329
rect 2940 35320 2943 35329
rect 2943 35320 2977 35329
rect 2977 35320 2992 35329
rect 2940 35282 2992 35320
rect 2940 35277 2943 35282
rect 2943 35277 2977 35282
rect 2977 35277 2992 35282
rect 3008 35320 3021 35329
rect 3021 35320 3055 35329
rect 3055 35320 3060 35329
rect 3008 35282 3060 35320
rect 3008 35277 3021 35282
rect 3021 35277 3055 35282
rect 3055 35277 3060 35282
rect 2872 35212 2924 35264
rect 2940 35248 2943 35264
rect 2943 35248 2977 35264
rect 2977 35248 2992 35264
rect 2940 35212 2992 35248
rect 3008 35248 3021 35264
rect 3021 35248 3055 35264
rect 3055 35248 3060 35264
rect 3008 35212 3060 35248
rect 2872 35147 2924 35199
rect 2940 35176 2943 35199
rect 2943 35176 2977 35199
rect 2977 35176 2992 35199
rect 2940 35147 2992 35176
rect 3008 35176 3021 35199
rect 3021 35176 3055 35199
rect 3055 35176 3060 35199
rect 3008 35147 3060 35176
rect 2872 35082 2924 35134
rect 2940 35104 2943 35134
rect 2943 35104 2977 35134
rect 2977 35104 2992 35134
rect 2940 35082 2992 35104
rect 3008 35104 3021 35134
rect 3021 35104 3055 35134
rect 3055 35104 3060 35134
rect 3008 35082 3060 35104
rect 2872 35017 2924 35069
rect 2940 35066 2992 35069
rect 2940 35032 2943 35066
rect 2943 35032 2977 35066
rect 2977 35032 2992 35066
rect 2940 35017 2992 35032
rect 3008 35066 3060 35069
rect 3008 35032 3021 35066
rect 3021 35032 3055 35066
rect 3055 35032 3060 35066
rect 3008 35017 3060 35032
rect 2872 34952 2924 35004
rect 2940 34994 2992 35004
rect 2940 34960 2943 34994
rect 2943 34960 2977 34994
rect 2977 34960 2992 34994
rect 2940 34952 2992 34960
rect 3008 34994 3060 35004
rect 3008 34960 3021 34994
rect 3021 34960 3055 34994
rect 3055 34960 3060 34994
rect 3008 34952 3060 34960
rect 2872 34887 2924 34939
rect 2940 34922 2992 34939
rect 2940 34888 2943 34922
rect 2943 34888 2977 34922
rect 2977 34888 2992 34922
rect 2940 34887 2992 34888
rect 3008 34922 3060 34939
rect 3008 34888 3021 34922
rect 3021 34888 3055 34922
rect 3055 34888 3060 34922
rect 3008 34887 3060 34888
rect 2872 34822 2924 34874
rect 2940 34850 2992 34874
rect 2940 34822 2943 34850
rect 2943 34822 2977 34850
rect 2977 34822 2992 34850
rect 3008 34850 3060 34874
rect 3008 34822 3021 34850
rect 3021 34822 3055 34850
rect 3055 34822 3060 34850
rect 2872 34757 2924 34809
rect 2940 34778 2992 34809
rect 2940 34757 2943 34778
rect 2943 34757 2977 34778
rect 2977 34757 2992 34778
rect 3008 34778 3060 34809
rect 3008 34757 3021 34778
rect 3021 34757 3055 34778
rect 3055 34757 3060 34778
rect 2872 34692 2924 34744
rect 2940 34706 2992 34744
rect 2940 34692 2943 34706
rect 2943 34692 2977 34706
rect 2977 34692 2992 34706
rect 3008 34706 3060 34744
rect 3008 34692 3021 34706
rect 3021 34692 3055 34706
rect 3055 34692 3060 34706
rect 2872 34627 2924 34679
rect 2940 34672 2943 34679
rect 2943 34672 2977 34679
rect 2977 34672 2992 34679
rect 2940 34634 2992 34672
rect 2940 34627 2943 34634
rect 2943 34627 2977 34634
rect 2977 34627 2992 34634
rect 3008 34672 3021 34679
rect 3021 34672 3055 34679
rect 3055 34672 3060 34679
rect 3008 34634 3060 34672
rect 3008 34627 3021 34634
rect 3021 34627 3055 34634
rect 3055 34627 3060 34634
rect 2872 34562 2924 34614
rect 2940 34600 2943 34614
rect 2943 34600 2977 34614
rect 2977 34600 2992 34614
rect 2940 34562 2992 34600
rect 3008 34600 3021 34614
rect 3021 34600 3055 34614
rect 3055 34600 3060 34614
rect 3008 34562 3060 34600
rect 3361 37945 3413 37997
rect 3439 37945 3491 37997
rect 3361 37877 3413 37929
rect 3439 37877 3491 37929
rect 3361 37809 3413 37861
rect 3439 37809 3491 37861
rect 3361 37741 3413 37793
rect 3439 37741 3491 37793
rect 3361 37673 3413 37725
rect 3439 37673 3491 37725
rect 3361 37605 3413 37657
rect 3439 37605 3491 37657
rect 3361 37537 3413 37589
rect 3439 37537 3491 37589
rect 3361 37469 3413 37521
rect 3439 37469 3491 37521
rect 3361 37401 3413 37453
rect 3439 37401 3491 37453
rect 3361 37333 3413 37385
rect 3439 37333 3491 37385
rect 3361 37266 3413 37318
rect 3439 37266 3491 37318
rect 3361 37199 3413 37251
rect 3439 37199 3491 37251
rect 3361 37132 3413 37184
rect 3439 37132 3491 37184
rect 3361 37065 3413 37117
rect 3439 37065 3491 37117
rect 3361 34173 3413 34225
rect 3439 34173 3491 34225
rect 3361 34109 3413 34161
rect 3439 34109 3491 34161
rect 3361 34045 3413 34097
rect 3439 34045 3491 34097
rect 3361 33981 3413 34033
rect 3439 33981 3491 34033
rect 3361 33917 3413 33969
rect 3439 33917 3491 33969
rect 3361 33853 3413 33905
rect 3439 33853 3491 33905
rect 3361 33789 3413 33841
rect 3439 33789 3491 33841
rect 3361 33725 3413 33777
rect 3439 33725 3491 33777
rect 3361 33661 3413 33713
rect 3439 33661 3491 33713
rect 3361 33597 3413 33649
rect 3439 33597 3491 33649
rect 3361 33533 3413 33585
rect 3439 33533 3491 33585
rect 3361 33469 3413 33521
rect 3439 33469 3491 33521
rect 3361 33405 3413 33457
rect 3439 33405 3491 33457
rect 3361 33341 3413 33393
rect 3439 33341 3491 33393
rect 3361 33277 3413 33329
rect 3439 33277 3491 33329
rect 3361 33212 3413 33264
rect 3439 33212 3491 33264
rect 3361 33147 3413 33199
rect 3439 33147 3491 33199
rect 3361 33082 3413 33134
rect 3439 33082 3491 33134
rect 3361 33017 3413 33069
rect 3439 33017 3491 33069
rect 3361 32952 3413 33004
rect 3439 32952 3491 33004
rect 3361 32887 3413 32939
rect 3439 32887 3491 32939
rect 3361 32822 3413 32874
rect 3439 32822 3491 32874
rect 3361 32757 3413 32809
rect 3439 32757 3491 32809
rect 3361 32692 3413 32744
rect 3439 32692 3491 32744
rect 3361 32627 3413 32679
rect 3439 32627 3491 32679
rect 3361 32562 3413 32614
rect 3439 32562 3491 32614
rect 3361 32497 3413 32549
rect 3439 32497 3491 32549
rect 2872 31762 2924 31768
rect 2940 31762 2992 31768
rect 3008 31762 3060 31768
rect 2872 31716 2877 31762
rect 2877 31716 2924 31762
rect 2940 31716 2992 31762
rect 3008 31716 3055 31762
rect 3055 31716 3060 31762
rect 2872 31652 2877 31704
rect 2877 31652 2924 31704
rect 2940 31652 2992 31704
rect 3008 31652 3055 31704
rect 3055 31652 3060 31704
rect 2872 31587 2877 31639
rect 2877 31587 2924 31639
rect 2940 31587 2992 31639
rect 3008 31587 3055 31639
rect 3055 31587 3060 31639
rect 2872 31522 2877 31574
rect 2877 31522 2924 31574
rect 2940 31522 2992 31574
rect 3008 31522 3055 31574
rect 3055 31522 3060 31574
rect 2872 31457 2877 31509
rect 2877 31457 2924 31509
rect 2940 31457 2992 31509
rect 3008 31457 3055 31509
rect 3055 31457 3060 31509
rect 2872 31392 2877 31444
rect 2877 31392 2924 31444
rect 2940 31392 2992 31444
rect 3008 31392 3055 31444
rect 3055 31392 3060 31444
rect 2872 31327 2877 31379
rect 2877 31327 2924 31379
rect 2940 31327 2992 31379
rect 3008 31327 3055 31379
rect 3055 31327 3060 31379
rect 2872 31262 2877 31314
rect 2877 31262 2924 31314
rect 2940 31262 2992 31314
rect 3008 31262 3055 31314
rect 3055 31262 3060 31314
rect 2872 31197 2877 31249
rect 2877 31197 2924 31249
rect 2940 31197 2992 31249
rect 3008 31197 3055 31249
rect 3055 31197 3060 31249
rect 2872 31132 2877 31184
rect 2877 31132 2924 31184
rect 2940 31132 2992 31184
rect 3008 31132 3055 31184
rect 3055 31132 3060 31184
rect 2872 31067 2877 31119
rect 2877 31067 2924 31119
rect 2940 31067 2992 31119
rect 3008 31067 3055 31119
rect 3055 31067 3060 31119
rect 2872 31002 2877 31054
rect 2877 31002 2924 31054
rect 2940 31002 2992 31054
rect 3008 31002 3055 31054
rect 3055 31002 3060 31054
rect 2872 30937 2877 30989
rect 2877 30937 2924 30989
rect 2940 30937 2992 30989
rect 3008 30937 3055 30989
rect 3055 30937 3060 30989
rect 2872 30872 2877 30924
rect 2877 30872 2924 30924
rect 2940 30872 2992 30924
rect 3008 30872 3055 30924
rect 3055 30872 3060 30924
rect 2872 30807 2877 30859
rect 2877 30807 2924 30859
rect 2940 30807 2992 30859
rect 3008 30807 3055 30859
rect 3055 30807 3060 30859
rect 2872 30742 2877 30794
rect 2877 30742 2924 30794
rect 2940 30742 2992 30794
rect 3008 30742 3055 30794
rect 3055 30742 3060 30794
rect 2872 30677 2877 30729
rect 2877 30677 2924 30729
rect 2940 30677 2992 30729
rect 3008 30677 3055 30729
rect 3055 30677 3060 30729
rect 2872 30612 2877 30664
rect 2877 30612 2924 30664
rect 2940 30612 2992 30664
rect 3008 30612 3055 30664
rect 3055 30612 3060 30664
rect 2872 30547 2877 30599
rect 2877 30547 2924 30599
rect 2940 30547 2992 30599
rect 3008 30547 3055 30599
rect 3055 30547 3060 30599
rect 2872 30482 2877 30534
rect 2877 30482 2924 30534
rect 2940 30482 2992 30534
rect 3008 30482 3055 30534
rect 3055 30482 3060 30534
rect 2872 30417 2877 30469
rect 2877 30417 2924 30469
rect 2940 30417 2992 30469
rect 3008 30417 3055 30469
rect 3055 30417 3060 30469
rect 2872 30352 2877 30404
rect 2877 30352 2924 30404
rect 2940 30352 2992 30404
rect 3008 30352 3055 30404
rect 3055 30352 3060 30404
rect 2872 30287 2877 30339
rect 2877 30287 2924 30339
rect 2940 30287 2992 30339
rect 3008 30287 3055 30339
rect 3055 30287 3060 30339
rect 2872 30222 2877 30274
rect 2877 30222 2924 30274
rect 2940 30222 2992 30274
rect 3008 30222 3055 30274
rect 3055 30222 3060 30274
rect 2872 30157 2877 30209
rect 2877 30157 2924 30209
rect 2940 30157 2992 30209
rect 3008 30157 3055 30209
rect 3055 30157 3060 30209
rect 2872 30092 2877 30144
rect 2877 30092 2924 30144
rect 2940 30092 2992 30144
rect 3008 30092 3055 30144
rect 3055 30092 3060 30144
rect 2872 30027 2877 30079
rect 2877 30027 2924 30079
rect 2940 30027 2992 30079
rect 3008 30027 3055 30079
rect 3055 30027 3060 30079
rect 2872 29962 2877 30014
rect 2877 29962 2924 30014
rect 2940 29962 2992 30014
rect 3008 29962 3055 30014
rect 3055 29962 3060 30014
rect 3361 29284 3413 29336
rect 3439 29284 3491 29336
rect 3361 29218 3413 29270
rect 3439 29218 3491 29270
rect 3361 29152 3413 29204
rect 3439 29152 3491 29204
rect 3361 29086 3413 29138
rect 3439 29086 3491 29138
rect 3361 29020 3413 29072
rect 3439 29020 3491 29072
rect 3361 28954 3413 29006
rect 3439 28954 3491 29006
rect 3361 28888 3413 28940
rect 3439 28888 3491 28940
rect 3361 28822 3413 28874
rect 3439 28822 3491 28874
rect 3361 28756 3413 28808
rect 3439 28756 3491 28808
rect 3361 28690 3413 28742
rect 3439 28690 3491 28742
rect 3361 28624 3413 28676
rect 3439 28624 3491 28676
rect 3361 28558 3413 28610
rect 3439 28558 3491 28610
rect 3361 28492 3413 28544
rect 3439 28492 3491 28544
rect 3361 28426 3413 28478
rect 3439 28426 3491 28478
rect 3361 28360 3413 28412
rect 3439 28360 3491 28412
rect 3361 28294 3413 28346
rect 3439 28294 3491 28346
rect 3361 28228 3413 28280
rect 3439 28228 3491 28280
rect 3361 28162 3413 28214
rect 3439 28162 3491 28214
rect 3361 28096 3413 28148
rect 3439 28096 3491 28148
rect 3361 28030 3413 28082
rect 3439 28030 3491 28082
rect 3361 27964 3413 28016
rect 3439 27964 3491 28016
rect 3361 27897 3413 27949
rect 3439 27897 3491 27949
rect 4712 39006 4764 39009
rect 4712 38972 4717 39006
rect 4717 38972 4751 39006
rect 4751 38972 4764 39006
rect 4712 38957 4764 38972
rect 4780 39006 4832 39009
rect 4780 38972 4789 39006
rect 4789 38972 4823 39006
rect 4823 38972 4832 39006
rect 4780 38957 4832 38972
rect 4848 39006 4900 39009
rect 4848 38972 4861 39006
rect 4861 38972 4895 39006
rect 4895 38972 4900 39006
rect 4848 38957 4900 38972
rect 4712 38932 4764 38944
rect 4712 38898 4717 38932
rect 4717 38898 4751 38932
rect 4751 38898 4764 38932
rect 4712 38892 4764 38898
rect 4780 38932 4832 38944
rect 4780 38898 4789 38932
rect 4789 38898 4823 38932
rect 4823 38898 4832 38932
rect 4780 38892 4832 38898
rect 4848 38932 4900 38944
rect 4848 38898 4861 38932
rect 4861 38898 4895 38932
rect 4895 38898 4900 38932
rect 4848 38892 4900 38898
rect 4712 38858 4764 38879
rect 4712 38827 4717 38858
rect 4717 38827 4751 38858
rect 4751 38827 4764 38858
rect 4780 38858 4832 38879
rect 4780 38827 4789 38858
rect 4789 38827 4823 38858
rect 4823 38827 4832 38858
rect 4848 38858 4900 38879
rect 4848 38827 4861 38858
rect 4861 38827 4895 38858
rect 4895 38827 4900 38858
rect 4712 38784 4764 38814
rect 4712 38762 4717 38784
rect 4717 38762 4751 38784
rect 4751 38762 4764 38784
rect 4780 38784 4832 38814
rect 4780 38762 4789 38784
rect 4789 38762 4823 38784
rect 4823 38762 4832 38784
rect 4848 38784 4900 38814
rect 4848 38762 4861 38784
rect 4861 38762 4895 38784
rect 4895 38762 4900 38784
rect 4712 38710 4764 38749
rect 4712 38697 4717 38710
rect 4717 38697 4751 38710
rect 4751 38697 4764 38710
rect 4780 38710 4832 38749
rect 4780 38697 4789 38710
rect 4789 38697 4823 38710
rect 4823 38697 4832 38710
rect 4848 38710 4900 38749
rect 4848 38697 4861 38710
rect 4861 38697 4895 38710
rect 4895 38697 4900 38710
rect 4712 38676 4717 38684
rect 4717 38676 4751 38684
rect 4751 38676 4764 38684
rect 4712 38636 4764 38676
rect 4712 38632 4717 38636
rect 4717 38632 4751 38636
rect 4751 38632 4764 38636
rect 4780 38676 4789 38684
rect 4789 38676 4823 38684
rect 4823 38676 4832 38684
rect 4780 38636 4832 38676
rect 4780 38632 4789 38636
rect 4789 38632 4823 38636
rect 4823 38632 4832 38636
rect 4848 38676 4861 38684
rect 4861 38676 4895 38684
rect 4895 38676 4900 38684
rect 4848 38636 4900 38676
rect 4848 38632 4861 38636
rect 4861 38632 4895 38636
rect 4895 38632 4900 38636
rect 4712 38602 4717 38619
rect 4717 38602 4751 38619
rect 4751 38602 4764 38619
rect 4712 38567 4764 38602
rect 4780 38602 4789 38619
rect 4789 38602 4823 38619
rect 4823 38602 4832 38619
rect 4780 38567 4832 38602
rect 4848 38602 4861 38619
rect 4861 38602 4895 38619
rect 4895 38602 4900 38619
rect 4848 38567 4900 38602
rect 4712 38528 4717 38554
rect 4717 38528 4751 38554
rect 4751 38528 4764 38554
rect 4712 38502 4764 38528
rect 4780 38528 4789 38554
rect 4789 38528 4823 38554
rect 4823 38528 4832 38554
rect 4780 38502 4832 38528
rect 4848 38528 4861 38554
rect 4861 38528 4895 38554
rect 4895 38528 4900 38554
rect 4848 38502 4900 38528
rect 4712 38487 4764 38490
rect 4712 38453 4717 38487
rect 4717 38453 4751 38487
rect 4751 38453 4764 38487
rect 4712 38438 4764 38453
rect 4780 38487 4832 38490
rect 4780 38453 4789 38487
rect 4789 38453 4823 38487
rect 4823 38453 4832 38487
rect 4780 38438 4832 38453
rect 4848 38487 4900 38490
rect 4848 38453 4861 38487
rect 4861 38453 4895 38487
rect 4895 38453 4900 38487
rect 4848 38438 4900 38453
rect 4712 38412 4764 38426
rect 4712 38378 4717 38412
rect 4717 38378 4751 38412
rect 4751 38378 4764 38412
rect 4712 38374 4764 38378
rect 4780 38412 4832 38426
rect 4780 38378 4789 38412
rect 4789 38378 4823 38412
rect 4823 38378 4832 38412
rect 4780 38374 4832 38378
rect 4848 38412 4900 38426
rect 4848 38378 4861 38412
rect 4861 38378 4895 38412
rect 4895 38378 4900 38412
rect 4848 38374 4900 38378
rect 4712 38337 4764 38362
rect 4712 38310 4717 38337
rect 4717 38310 4751 38337
rect 4751 38310 4764 38337
rect 4780 38337 4832 38362
rect 4780 38310 4789 38337
rect 4789 38310 4823 38337
rect 4823 38310 4832 38337
rect 4848 38337 4900 38362
rect 4848 38310 4861 38337
rect 4861 38310 4895 38337
rect 4895 38310 4900 38337
rect 4712 38262 4764 38298
rect 4712 38246 4717 38262
rect 4717 38246 4751 38262
rect 4751 38246 4764 38262
rect 4780 38262 4832 38298
rect 4780 38246 4789 38262
rect 4789 38246 4823 38262
rect 4823 38246 4832 38262
rect 4848 38262 4900 38298
rect 4848 38246 4861 38262
rect 4861 38246 4895 38262
rect 4895 38246 4900 38262
rect 4712 38228 4717 38234
rect 4717 38228 4751 38234
rect 4751 38228 4764 38234
rect 4712 38187 4764 38228
rect 4712 38182 4717 38187
rect 4717 38182 4751 38187
rect 4751 38182 4764 38187
rect 4780 38228 4789 38234
rect 4789 38228 4823 38234
rect 4823 38228 4832 38234
rect 4780 38187 4832 38228
rect 4780 38182 4789 38187
rect 4789 38182 4823 38187
rect 4823 38182 4832 38187
rect 4848 38228 4861 38234
rect 4861 38228 4895 38234
rect 4895 38228 4900 38234
rect 4848 38187 4900 38228
rect 4848 38182 4861 38187
rect 4861 38182 4895 38187
rect 4895 38182 4900 38187
rect 4712 38153 4717 38170
rect 4717 38153 4751 38170
rect 4751 38153 4764 38170
rect 4712 38118 4764 38153
rect 4780 38153 4789 38170
rect 4789 38153 4823 38170
rect 4823 38153 4832 38170
rect 4780 38118 4832 38153
rect 4848 38153 4861 38170
rect 4861 38153 4895 38170
rect 4895 38153 4900 38170
rect 4848 38118 4900 38153
rect 5632 39006 5684 39009
rect 5632 38972 5637 39006
rect 5637 38972 5671 39006
rect 5671 38972 5684 39006
rect 5632 38957 5684 38972
rect 5700 39006 5752 39009
rect 5700 38972 5709 39006
rect 5709 38972 5743 39006
rect 5743 38972 5752 39006
rect 5700 38957 5752 38972
rect 5768 39006 5820 39009
rect 5768 38972 5781 39006
rect 5781 38972 5815 39006
rect 5815 38972 5820 39006
rect 5768 38957 5820 38972
rect 5632 38932 5684 38944
rect 5632 38898 5637 38932
rect 5637 38898 5671 38932
rect 5671 38898 5684 38932
rect 5632 38892 5684 38898
rect 5700 38932 5752 38944
rect 5700 38898 5709 38932
rect 5709 38898 5743 38932
rect 5743 38898 5752 38932
rect 5700 38892 5752 38898
rect 5768 38932 5820 38944
rect 5768 38898 5781 38932
rect 5781 38898 5815 38932
rect 5815 38898 5820 38932
rect 5768 38892 5820 38898
rect 5632 38858 5684 38879
rect 5632 38827 5637 38858
rect 5637 38827 5671 38858
rect 5671 38827 5684 38858
rect 5700 38858 5752 38879
rect 5700 38827 5709 38858
rect 5709 38827 5743 38858
rect 5743 38827 5752 38858
rect 5768 38858 5820 38879
rect 5768 38827 5781 38858
rect 5781 38827 5815 38858
rect 5815 38827 5820 38858
rect 5632 38784 5684 38814
rect 5632 38762 5637 38784
rect 5637 38762 5671 38784
rect 5671 38762 5684 38784
rect 5700 38784 5752 38814
rect 5700 38762 5709 38784
rect 5709 38762 5743 38784
rect 5743 38762 5752 38784
rect 5768 38784 5820 38814
rect 5768 38762 5781 38784
rect 5781 38762 5815 38784
rect 5815 38762 5820 38784
rect 5632 38710 5684 38749
rect 5632 38697 5637 38710
rect 5637 38697 5671 38710
rect 5671 38697 5684 38710
rect 5700 38710 5752 38749
rect 5700 38697 5709 38710
rect 5709 38697 5743 38710
rect 5743 38697 5752 38710
rect 5768 38710 5820 38749
rect 5768 38697 5781 38710
rect 5781 38697 5815 38710
rect 5815 38697 5820 38710
rect 5632 38676 5637 38684
rect 5637 38676 5671 38684
rect 5671 38676 5684 38684
rect 5632 38636 5684 38676
rect 5632 38632 5637 38636
rect 5637 38632 5671 38636
rect 5671 38632 5684 38636
rect 5700 38676 5709 38684
rect 5709 38676 5743 38684
rect 5743 38676 5752 38684
rect 5700 38636 5752 38676
rect 5700 38632 5709 38636
rect 5709 38632 5743 38636
rect 5743 38632 5752 38636
rect 5768 38676 5781 38684
rect 5781 38676 5815 38684
rect 5815 38676 5820 38684
rect 5768 38636 5820 38676
rect 5768 38632 5781 38636
rect 5781 38632 5815 38636
rect 5815 38632 5820 38636
rect 5632 38602 5637 38619
rect 5637 38602 5671 38619
rect 5671 38602 5684 38619
rect 5632 38567 5684 38602
rect 5700 38602 5709 38619
rect 5709 38602 5743 38619
rect 5743 38602 5752 38619
rect 5700 38567 5752 38602
rect 5768 38602 5781 38619
rect 5781 38602 5815 38619
rect 5815 38602 5820 38619
rect 5768 38567 5820 38602
rect 5632 38528 5637 38554
rect 5637 38528 5671 38554
rect 5671 38528 5684 38554
rect 5632 38502 5684 38528
rect 5700 38528 5709 38554
rect 5709 38528 5743 38554
rect 5743 38528 5752 38554
rect 5700 38502 5752 38528
rect 5768 38528 5781 38554
rect 5781 38528 5815 38554
rect 5815 38528 5820 38554
rect 5768 38502 5820 38528
rect 5632 38487 5684 38490
rect 5632 38453 5637 38487
rect 5637 38453 5671 38487
rect 5671 38453 5684 38487
rect 5632 38438 5684 38453
rect 5700 38487 5752 38490
rect 5700 38453 5709 38487
rect 5709 38453 5743 38487
rect 5743 38453 5752 38487
rect 5700 38438 5752 38453
rect 5768 38487 5820 38490
rect 5768 38453 5781 38487
rect 5781 38453 5815 38487
rect 5815 38453 5820 38487
rect 5768 38438 5820 38453
rect 5632 38412 5684 38426
rect 5632 38378 5637 38412
rect 5637 38378 5671 38412
rect 5671 38378 5684 38412
rect 5632 38374 5684 38378
rect 5700 38412 5752 38426
rect 5700 38378 5709 38412
rect 5709 38378 5743 38412
rect 5743 38378 5752 38412
rect 5700 38374 5752 38378
rect 5768 38412 5820 38426
rect 5768 38378 5781 38412
rect 5781 38378 5815 38412
rect 5815 38378 5820 38412
rect 5768 38374 5820 38378
rect 5632 38337 5684 38362
rect 5632 38310 5637 38337
rect 5637 38310 5671 38337
rect 5671 38310 5684 38337
rect 5700 38337 5752 38362
rect 5700 38310 5709 38337
rect 5709 38310 5743 38337
rect 5743 38310 5752 38337
rect 5768 38337 5820 38362
rect 5768 38310 5781 38337
rect 5781 38310 5815 38337
rect 5815 38310 5820 38337
rect 5632 38262 5684 38298
rect 5632 38246 5637 38262
rect 5637 38246 5671 38262
rect 5671 38246 5684 38262
rect 5700 38262 5752 38298
rect 5700 38246 5709 38262
rect 5709 38246 5743 38262
rect 5743 38246 5752 38262
rect 5768 38262 5820 38298
rect 5768 38246 5781 38262
rect 5781 38246 5815 38262
rect 5815 38246 5820 38262
rect 5632 38228 5637 38234
rect 5637 38228 5671 38234
rect 5671 38228 5684 38234
rect 5632 38187 5684 38228
rect 5632 38182 5637 38187
rect 5637 38182 5671 38187
rect 5671 38182 5684 38187
rect 5700 38228 5709 38234
rect 5709 38228 5743 38234
rect 5743 38228 5752 38234
rect 5700 38187 5752 38228
rect 5700 38182 5709 38187
rect 5709 38182 5743 38187
rect 5743 38182 5752 38187
rect 5768 38228 5781 38234
rect 5781 38228 5815 38234
rect 5815 38228 5820 38234
rect 5768 38187 5820 38228
rect 5768 38182 5781 38187
rect 5781 38182 5815 38187
rect 5815 38182 5820 38187
rect 5632 38153 5637 38170
rect 5637 38153 5671 38170
rect 5671 38153 5684 38170
rect 5632 38118 5684 38153
rect 5700 38153 5709 38170
rect 5709 38153 5743 38170
rect 5743 38153 5752 38170
rect 5700 38118 5752 38153
rect 5768 38153 5781 38170
rect 5781 38153 5815 38170
rect 5815 38153 5820 38170
rect 5768 38118 5820 38153
rect 6552 39006 6604 39009
rect 6552 38972 6557 39006
rect 6557 38972 6591 39006
rect 6591 38972 6604 39006
rect 6552 38957 6604 38972
rect 6620 39006 6672 39009
rect 6620 38972 6629 39006
rect 6629 38972 6663 39006
rect 6663 38972 6672 39006
rect 6620 38957 6672 38972
rect 6688 39006 6740 39009
rect 6688 38972 6701 39006
rect 6701 38972 6735 39006
rect 6735 38972 6740 39006
rect 6688 38957 6740 38972
rect 6552 38932 6604 38944
rect 6552 38898 6557 38932
rect 6557 38898 6591 38932
rect 6591 38898 6604 38932
rect 6552 38892 6604 38898
rect 6620 38932 6672 38944
rect 6620 38898 6629 38932
rect 6629 38898 6663 38932
rect 6663 38898 6672 38932
rect 6620 38892 6672 38898
rect 6688 38932 6740 38944
rect 6688 38898 6701 38932
rect 6701 38898 6735 38932
rect 6735 38898 6740 38932
rect 6688 38892 6740 38898
rect 6552 38858 6604 38879
rect 6552 38827 6557 38858
rect 6557 38827 6591 38858
rect 6591 38827 6604 38858
rect 6620 38858 6672 38879
rect 6620 38827 6629 38858
rect 6629 38827 6663 38858
rect 6663 38827 6672 38858
rect 6688 38858 6740 38879
rect 6688 38827 6701 38858
rect 6701 38827 6735 38858
rect 6735 38827 6740 38858
rect 6552 38784 6604 38814
rect 6552 38762 6557 38784
rect 6557 38762 6591 38784
rect 6591 38762 6604 38784
rect 6620 38784 6672 38814
rect 6620 38762 6629 38784
rect 6629 38762 6663 38784
rect 6663 38762 6672 38784
rect 6688 38784 6740 38814
rect 6688 38762 6701 38784
rect 6701 38762 6735 38784
rect 6735 38762 6740 38784
rect 6552 38710 6604 38749
rect 6552 38697 6557 38710
rect 6557 38697 6591 38710
rect 6591 38697 6604 38710
rect 6620 38710 6672 38749
rect 6620 38697 6629 38710
rect 6629 38697 6663 38710
rect 6663 38697 6672 38710
rect 6688 38710 6740 38749
rect 6688 38697 6701 38710
rect 6701 38697 6735 38710
rect 6735 38697 6740 38710
rect 6552 38676 6557 38684
rect 6557 38676 6591 38684
rect 6591 38676 6604 38684
rect 6552 38636 6604 38676
rect 6552 38632 6557 38636
rect 6557 38632 6591 38636
rect 6591 38632 6604 38636
rect 6620 38676 6629 38684
rect 6629 38676 6663 38684
rect 6663 38676 6672 38684
rect 6620 38636 6672 38676
rect 6620 38632 6629 38636
rect 6629 38632 6663 38636
rect 6663 38632 6672 38636
rect 6688 38676 6701 38684
rect 6701 38676 6735 38684
rect 6735 38676 6740 38684
rect 6688 38636 6740 38676
rect 6688 38632 6701 38636
rect 6701 38632 6735 38636
rect 6735 38632 6740 38636
rect 6552 38602 6557 38619
rect 6557 38602 6591 38619
rect 6591 38602 6604 38619
rect 6552 38567 6604 38602
rect 6620 38602 6629 38619
rect 6629 38602 6663 38619
rect 6663 38602 6672 38619
rect 6620 38567 6672 38602
rect 6688 38602 6701 38619
rect 6701 38602 6735 38619
rect 6735 38602 6740 38619
rect 6688 38567 6740 38602
rect 6552 38528 6557 38554
rect 6557 38528 6591 38554
rect 6591 38528 6604 38554
rect 6552 38502 6604 38528
rect 6620 38528 6629 38554
rect 6629 38528 6663 38554
rect 6663 38528 6672 38554
rect 6620 38502 6672 38528
rect 6688 38528 6701 38554
rect 6701 38528 6735 38554
rect 6735 38528 6740 38554
rect 6688 38502 6740 38528
rect 6552 38487 6604 38490
rect 6552 38453 6557 38487
rect 6557 38453 6591 38487
rect 6591 38453 6604 38487
rect 6552 38438 6604 38453
rect 6620 38487 6672 38490
rect 6620 38453 6629 38487
rect 6629 38453 6663 38487
rect 6663 38453 6672 38487
rect 6620 38438 6672 38453
rect 6688 38487 6740 38490
rect 6688 38453 6701 38487
rect 6701 38453 6735 38487
rect 6735 38453 6740 38487
rect 6688 38438 6740 38453
rect 6552 38412 6604 38426
rect 6552 38378 6557 38412
rect 6557 38378 6591 38412
rect 6591 38378 6604 38412
rect 6552 38374 6604 38378
rect 6620 38412 6672 38426
rect 6620 38378 6629 38412
rect 6629 38378 6663 38412
rect 6663 38378 6672 38412
rect 6620 38374 6672 38378
rect 6688 38412 6740 38426
rect 6688 38378 6701 38412
rect 6701 38378 6735 38412
rect 6735 38378 6740 38412
rect 6688 38374 6740 38378
rect 6552 38337 6604 38362
rect 6552 38310 6557 38337
rect 6557 38310 6591 38337
rect 6591 38310 6604 38337
rect 6620 38337 6672 38362
rect 6620 38310 6629 38337
rect 6629 38310 6663 38337
rect 6663 38310 6672 38337
rect 6688 38337 6740 38362
rect 6688 38310 6701 38337
rect 6701 38310 6735 38337
rect 6735 38310 6740 38337
rect 6552 38262 6604 38298
rect 6552 38246 6557 38262
rect 6557 38246 6591 38262
rect 6591 38246 6604 38262
rect 6620 38262 6672 38298
rect 6620 38246 6629 38262
rect 6629 38246 6663 38262
rect 6663 38246 6672 38262
rect 6688 38262 6740 38298
rect 6688 38246 6701 38262
rect 6701 38246 6735 38262
rect 6735 38246 6740 38262
rect 6552 38228 6557 38234
rect 6557 38228 6591 38234
rect 6591 38228 6604 38234
rect 6552 38187 6604 38228
rect 6552 38182 6557 38187
rect 6557 38182 6591 38187
rect 6591 38182 6604 38187
rect 6620 38228 6629 38234
rect 6629 38228 6663 38234
rect 6663 38228 6672 38234
rect 6620 38187 6672 38228
rect 6620 38182 6629 38187
rect 6629 38182 6663 38187
rect 6663 38182 6672 38187
rect 6688 38228 6701 38234
rect 6701 38228 6735 38234
rect 6735 38228 6740 38234
rect 6688 38187 6740 38228
rect 6688 38182 6701 38187
rect 6701 38182 6735 38187
rect 6735 38182 6740 38187
rect 6552 38153 6557 38170
rect 6557 38153 6591 38170
rect 6591 38153 6604 38170
rect 6552 38118 6604 38153
rect 6620 38153 6629 38170
rect 6629 38153 6663 38170
rect 6663 38153 6672 38170
rect 6620 38118 6672 38153
rect 6688 38153 6701 38170
rect 6701 38153 6735 38170
rect 6735 38153 6740 38170
rect 6688 38118 6740 38153
rect 7472 39006 7524 39009
rect 7472 38972 7477 39006
rect 7477 38972 7511 39006
rect 7511 38972 7524 39006
rect 7472 38957 7524 38972
rect 7540 39006 7592 39009
rect 7540 38972 7549 39006
rect 7549 38972 7583 39006
rect 7583 38972 7592 39006
rect 7540 38957 7592 38972
rect 7608 39006 7660 39009
rect 7608 38972 7621 39006
rect 7621 38972 7655 39006
rect 7655 38972 7660 39006
rect 7608 38957 7660 38972
rect 7472 38932 7524 38944
rect 7472 38898 7477 38932
rect 7477 38898 7511 38932
rect 7511 38898 7524 38932
rect 7472 38892 7524 38898
rect 7540 38932 7592 38944
rect 7540 38898 7549 38932
rect 7549 38898 7583 38932
rect 7583 38898 7592 38932
rect 7540 38892 7592 38898
rect 7608 38932 7660 38944
rect 7608 38898 7621 38932
rect 7621 38898 7655 38932
rect 7655 38898 7660 38932
rect 7608 38892 7660 38898
rect 7472 38858 7524 38879
rect 7472 38827 7477 38858
rect 7477 38827 7511 38858
rect 7511 38827 7524 38858
rect 7540 38858 7592 38879
rect 7540 38827 7549 38858
rect 7549 38827 7583 38858
rect 7583 38827 7592 38858
rect 7608 38858 7660 38879
rect 7608 38827 7621 38858
rect 7621 38827 7655 38858
rect 7655 38827 7660 38858
rect 7472 38784 7524 38814
rect 7472 38762 7477 38784
rect 7477 38762 7511 38784
rect 7511 38762 7524 38784
rect 7540 38784 7592 38814
rect 7540 38762 7549 38784
rect 7549 38762 7583 38784
rect 7583 38762 7592 38784
rect 7608 38784 7660 38814
rect 7608 38762 7621 38784
rect 7621 38762 7655 38784
rect 7655 38762 7660 38784
rect 7472 38710 7524 38749
rect 7472 38697 7477 38710
rect 7477 38697 7511 38710
rect 7511 38697 7524 38710
rect 7540 38710 7592 38749
rect 7540 38697 7549 38710
rect 7549 38697 7583 38710
rect 7583 38697 7592 38710
rect 7608 38710 7660 38749
rect 7608 38697 7621 38710
rect 7621 38697 7655 38710
rect 7655 38697 7660 38710
rect 7472 38676 7477 38684
rect 7477 38676 7511 38684
rect 7511 38676 7524 38684
rect 7472 38636 7524 38676
rect 7472 38632 7477 38636
rect 7477 38632 7511 38636
rect 7511 38632 7524 38636
rect 7540 38676 7549 38684
rect 7549 38676 7583 38684
rect 7583 38676 7592 38684
rect 7540 38636 7592 38676
rect 7540 38632 7549 38636
rect 7549 38632 7583 38636
rect 7583 38632 7592 38636
rect 7608 38676 7621 38684
rect 7621 38676 7655 38684
rect 7655 38676 7660 38684
rect 7608 38636 7660 38676
rect 7608 38632 7621 38636
rect 7621 38632 7655 38636
rect 7655 38632 7660 38636
rect 7472 38602 7477 38619
rect 7477 38602 7511 38619
rect 7511 38602 7524 38619
rect 7472 38567 7524 38602
rect 7540 38602 7549 38619
rect 7549 38602 7583 38619
rect 7583 38602 7592 38619
rect 7540 38567 7592 38602
rect 7608 38602 7621 38619
rect 7621 38602 7655 38619
rect 7655 38602 7660 38619
rect 7608 38567 7660 38602
rect 7472 38528 7477 38554
rect 7477 38528 7511 38554
rect 7511 38528 7524 38554
rect 7472 38502 7524 38528
rect 7540 38528 7549 38554
rect 7549 38528 7583 38554
rect 7583 38528 7592 38554
rect 7540 38502 7592 38528
rect 7608 38528 7621 38554
rect 7621 38528 7655 38554
rect 7655 38528 7660 38554
rect 7608 38502 7660 38528
rect 7472 38487 7524 38490
rect 7472 38453 7477 38487
rect 7477 38453 7511 38487
rect 7511 38453 7524 38487
rect 7472 38438 7524 38453
rect 7540 38487 7592 38490
rect 7540 38453 7549 38487
rect 7549 38453 7583 38487
rect 7583 38453 7592 38487
rect 7540 38438 7592 38453
rect 7608 38487 7660 38490
rect 7608 38453 7621 38487
rect 7621 38453 7655 38487
rect 7655 38453 7660 38487
rect 7608 38438 7660 38453
rect 7472 38412 7524 38426
rect 7472 38378 7477 38412
rect 7477 38378 7511 38412
rect 7511 38378 7524 38412
rect 7472 38374 7524 38378
rect 7540 38412 7592 38426
rect 7540 38378 7549 38412
rect 7549 38378 7583 38412
rect 7583 38378 7592 38412
rect 7540 38374 7592 38378
rect 7608 38412 7660 38426
rect 7608 38378 7621 38412
rect 7621 38378 7655 38412
rect 7655 38378 7660 38412
rect 7608 38374 7660 38378
rect 7472 38337 7524 38362
rect 7472 38310 7477 38337
rect 7477 38310 7511 38337
rect 7511 38310 7524 38337
rect 7540 38337 7592 38362
rect 7540 38310 7549 38337
rect 7549 38310 7583 38337
rect 7583 38310 7592 38337
rect 7608 38337 7660 38362
rect 7608 38310 7621 38337
rect 7621 38310 7655 38337
rect 7655 38310 7660 38337
rect 7472 38262 7524 38298
rect 7472 38246 7477 38262
rect 7477 38246 7511 38262
rect 7511 38246 7524 38262
rect 7540 38262 7592 38298
rect 7540 38246 7549 38262
rect 7549 38246 7583 38262
rect 7583 38246 7592 38262
rect 7608 38262 7660 38298
rect 7608 38246 7621 38262
rect 7621 38246 7655 38262
rect 7655 38246 7660 38262
rect 7472 38228 7477 38234
rect 7477 38228 7511 38234
rect 7511 38228 7524 38234
rect 7472 38187 7524 38228
rect 7472 38182 7477 38187
rect 7477 38182 7511 38187
rect 7511 38182 7524 38187
rect 7540 38228 7549 38234
rect 7549 38228 7583 38234
rect 7583 38228 7592 38234
rect 7540 38187 7592 38228
rect 7540 38182 7549 38187
rect 7549 38182 7583 38187
rect 7583 38182 7592 38187
rect 7608 38228 7621 38234
rect 7621 38228 7655 38234
rect 7655 38228 7660 38234
rect 7608 38187 7660 38228
rect 7608 38182 7621 38187
rect 7621 38182 7655 38187
rect 7655 38182 7660 38187
rect 7472 38153 7477 38170
rect 7477 38153 7511 38170
rect 7511 38153 7524 38170
rect 7472 38118 7524 38153
rect 7540 38153 7549 38170
rect 7549 38153 7583 38170
rect 7583 38153 7592 38170
rect 7540 38118 7592 38153
rect 7608 38153 7621 38170
rect 7621 38153 7655 38170
rect 7655 38153 7660 38170
rect 7608 38118 7660 38153
rect 8392 39006 8444 39009
rect 8392 38972 8397 39006
rect 8397 38972 8431 39006
rect 8431 38972 8444 39006
rect 8392 38957 8444 38972
rect 8460 39006 8512 39009
rect 8460 38972 8469 39006
rect 8469 38972 8503 39006
rect 8503 38972 8512 39006
rect 8460 38957 8512 38972
rect 8528 39006 8580 39009
rect 8528 38972 8541 39006
rect 8541 38972 8575 39006
rect 8575 38972 8580 39006
rect 8528 38957 8580 38972
rect 8392 38932 8444 38944
rect 8392 38898 8397 38932
rect 8397 38898 8431 38932
rect 8431 38898 8444 38932
rect 8392 38892 8444 38898
rect 8460 38932 8512 38944
rect 8460 38898 8469 38932
rect 8469 38898 8503 38932
rect 8503 38898 8512 38932
rect 8460 38892 8512 38898
rect 8528 38932 8580 38944
rect 8528 38898 8541 38932
rect 8541 38898 8575 38932
rect 8575 38898 8580 38932
rect 8528 38892 8580 38898
rect 8392 38858 8444 38879
rect 8392 38827 8397 38858
rect 8397 38827 8431 38858
rect 8431 38827 8444 38858
rect 8460 38858 8512 38879
rect 8460 38827 8469 38858
rect 8469 38827 8503 38858
rect 8503 38827 8512 38858
rect 8528 38858 8580 38879
rect 8528 38827 8541 38858
rect 8541 38827 8575 38858
rect 8575 38827 8580 38858
rect 8392 38784 8444 38814
rect 8392 38762 8397 38784
rect 8397 38762 8431 38784
rect 8431 38762 8444 38784
rect 8460 38784 8512 38814
rect 8460 38762 8469 38784
rect 8469 38762 8503 38784
rect 8503 38762 8512 38784
rect 8528 38784 8580 38814
rect 8528 38762 8541 38784
rect 8541 38762 8575 38784
rect 8575 38762 8580 38784
rect 8392 38710 8444 38749
rect 8392 38697 8397 38710
rect 8397 38697 8431 38710
rect 8431 38697 8444 38710
rect 8460 38710 8512 38749
rect 8460 38697 8469 38710
rect 8469 38697 8503 38710
rect 8503 38697 8512 38710
rect 8528 38710 8580 38749
rect 8528 38697 8541 38710
rect 8541 38697 8575 38710
rect 8575 38697 8580 38710
rect 8392 38676 8397 38684
rect 8397 38676 8431 38684
rect 8431 38676 8444 38684
rect 8392 38636 8444 38676
rect 8392 38632 8397 38636
rect 8397 38632 8431 38636
rect 8431 38632 8444 38636
rect 8460 38676 8469 38684
rect 8469 38676 8503 38684
rect 8503 38676 8512 38684
rect 8460 38636 8512 38676
rect 8460 38632 8469 38636
rect 8469 38632 8503 38636
rect 8503 38632 8512 38636
rect 8528 38676 8541 38684
rect 8541 38676 8575 38684
rect 8575 38676 8580 38684
rect 8528 38636 8580 38676
rect 8528 38632 8541 38636
rect 8541 38632 8575 38636
rect 8575 38632 8580 38636
rect 8392 38602 8397 38619
rect 8397 38602 8431 38619
rect 8431 38602 8444 38619
rect 8392 38567 8444 38602
rect 8460 38602 8469 38619
rect 8469 38602 8503 38619
rect 8503 38602 8512 38619
rect 8460 38567 8512 38602
rect 8528 38602 8541 38619
rect 8541 38602 8575 38619
rect 8575 38602 8580 38619
rect 8528 38567 8580 38602
rect 8392 38528 8397 38554
rect 8397 38528 8431 38554
rect 8431 38528 8444 38554
rect 8392 38502 8444 38528
rect 8460 38528 8469 38554
rect 8469 38528 8503 38554
rect 8503 38528 8512 38554
rect 8460 38502 8512 38528
rect 8528 38528 8541 38554
rect 8541 38528 8575 38554
rect 8575 38528 8580 38554
rect 8528 38502 8580 38528
rect 8392 38487 8444 38490
rect 8392 38453 8397 38487
rect 8397 38453 8431 38487
rect 8431 38453 8444 38487
rect 8392 38438 8444 38453
rect 8460 38487 8512 38490
rect 8460 38453 8469 38487
rect 8469 38453 8503 38487
rect 8503 38453 8512 38487
rect 8460 38438 8512 38453
rect 8528 38487 8580 38490
rect 8528 38453 8541 38487
rect 8541 38453 8575 38487
rect 8575 38453 8580 38487
rect 8528 38438 8580 38453
rect 8392 38412 8444 38426
rect 8392 38378 8397 38412
rect 8397 38378 8431 38412
rect 8431 38378 8444 38412
rect 8392 38374 8444 38378
rect 8460 38412 8512 38426
rect 8460 38378 8469 38412
rect 8469 38378 8503 38412
rect 8503 38378 8512 38412
rect 8460 38374 8512 38378
rect 8528 38412 8580 38426
rect 8528 38378 8541 38412
rect 8541 38378 8575 38412
rect 8575 38378 8580 38412
rect 8528 38374 8580 38378
rect 8392 38337 8444 38362
rect 8392 38310 8397 38337
rect 8397 38310 8431 38337
rect 8431 38310 8444 38337
rect 8460 38337 8512 38362
rect 8460 38310 8469 38337
rect 8469 38310 8503 38337
rect 8503 38310 8512 38337
rect 8528 38337 8580 38362
rect 8528 38310 8541 38337
rect 8541 38310 8575 38337
rect 8575 38310 8580 38337
rect 8392 38262 8444 38298
rect 8392 38246 8397 38262
rect 8397 38246 8431 38262
rect 8431 38246 8444 38262
rect 8460 38262 8512 38298
rect 8460 38246 8469 38262
rect 8469 38246 8503 38262
rect 8503 38246 8512 38262
rect 8528 38262 8580 38298
rect 8528 38246 8541 38262
rect 8541 38246 8575 38262
rect 8575 38246 8580 38262
rect 8392 38228 8397 38234
rect 8397 38228 8431 38234
rect 8431 38228 8444 38234
rect 8392 38187 8444 38228
rect 8392 38182 8397 38187
rect 8397 38182 8431 38187
rect 8431 38182 8444 38187
rect 8460 38228 8469 38234
rect 8469 38228 8503 38234
rect 8503 38228 8512 38234
rect 8460 38187 8512 38228
rect 8460 38182 8469 38187
rect 8469 38182 8503 38187
rect 8503 38182 8512 38187
rect 8528 38228 8541 38234
rect 8541 38228 8575 38234
rect 8575 38228 8580 38234
rect 8528 38187 8580 38228
rect 8528 38182 8541 38187
rect 8541 38182 8575 38187
rect 8575 38182 8580 38187
rect 8392 38153 8397 38170
rect 8397 38153 8431 38170
rect 8431 38153 8444 38170
rect 8392 38118 8444 38153
rect 8460 38153 8469 38170
rect 8469 38153 8503 38170
rect 8503 38153 8512 38170
rect 8460 38118 8512 38153
rect 8528 38153 8541 38170
rect 8541 38153 8575 38170
rect 8575 38153 8580 38170
rect 8528 38118 8580 38153
rect 9312 39006 9364 39009
rect 9312 38972 9317 39006
rect 9317 38972 9351 39006
rect 9351 38972 9364 39006
rect 9312 38957 9364 38972
rect 9380 39006 9432 39009
rect 9380 38972 9389 39006
rect 9389 38972 9423 39006
rect 9423 38972 9432 39006
rect 9380 38957 9432 38972
rect 9448 39006 9500 39009
rect 9448 38972 9461 39006
rect 9461 38972 9495 39006
rect 9495 38972 9500 39006
rect 9448 38957 9500 38972
rect 9312 38932 9364 38944
rect 9312 38898 9317 38932
rect 9317 38898 9351 38932
rect 9351 38898 9364 38932
rect 9312 38892 9364 38898
rect 9380 38932 9432 38944
rect 9380 38898 9389 38932
rect 9389 38898 9423 38932
rect 9423 38898 9432 38932
rect 9380 38892 9432 38898
rect 9448 38932 9500 38944
rect 9448 38898 9461 38932
rect 9461 38898 9495 38932
rect 9495 38898 9500 38932
rect 9448 38892 9500 38898
rect 9312 38858 9364 38879
rect 9312 38827 9317 38858
rect 9317 38827 9351 38858
rect 9351 38827 9364 38858
rect 9380 38858 9432 38879
rect 9380 38827 9389 38858
rect 9389 38827 9423 38858
rect 9423 38827 9432 38858
rect 9448 38858 9500 38879
rect 9448 38827 9461 38858
rect 9461 38827 9495 38858
rect 9495 38827 9500 38858
rect 9312 38784 9364 38814
rect 9312 38762 9317 38784
rect 9317 38762 9351 38784
rect 9351 38762 9364 38784
rect 9380 38784 9432 38814
rect 9380 38762 9389 38784
rect 9389 38762 9423 38784
rect 9423 38762 9432 38784
rect 9448 38784 9500 38814
rect 9448 38762 9461 38784
rect 9461 38762 9495 38784
rect 9495 38762 9500 38784
rect 9312 38710 9364 38749
rect 9312 38697 9317 38710
rect 9317 38697 9351 38710
rect 9351 38697 9364 38710
rect 9380 38710 9432 38749
rect 9380 38697 9389 38710
rect 9389 38697 9423 38710
rect 9423 38697 9432 38710
rect 9448 38710 9500 38749
rect 9448 38697 9461 38710
rect 9461 38697 9495 38710
rect 9495 38697 9500 38710
rect 9312 38676 9317 38684
rect 9317 38676 9351 38684
rect 9351 38676 9364 38684
rect 9312 38636 9364 38676
rect 9312 38632 9317 38636
rect 9317 38632 9351 38636
rect 9351 38632 9364 38636
rect 9380 38676 9389 38684
rect 9389 38676 9423 38684
rect 9423 38676 9432 38684
rect 9380 38636 9432 38676
rect 9380 38632 9389 38636
rect 9389 38632 9423 38636
rect 9423 38632 9432 38636
rect 9448 38676 9461 38684
rect 9461 38676 9495 38684
rect 9495 38676 9500 38684
rect 9448 38636 9500 38676
rect 9448 38632 9461 38636
rect 9461 38632 9495 38636
rect 9495 38632 9500 38636
rect 9312 38602 9317 38619
rect 9317 38602 9351 38619
rect 9351 38602 9364 38619
rect 9312 38567 9364 38602
rect 9380 38602 9389 38619
rect 9389 38602 9423 38619
rect 9423 38602 9432 38619
rect 9380 38567 9432 38602
rect 9448 38602 9461 38619
rect 9461 38602 9495 38619
rect 9495 38602 9500 38619
rect 9448 38567 9500 38602
rect 9312 38528 9317 38554
rect 9317 38528 9351 38554
rect 9351 38528 9364 38554
rect 9312 38502 9364 38528
rect 9380 38528 9389 38554
rect 9389 38528 9423 38554
rect 9423 38528 9432 38554
rect 9380 38502 9432 38528
rect 9448 38528 9461 38554
rect 9461 38528 9495 38554
rect 9495 38528 9500 38554
rect 9448 38502 9500 38528
rect 9312 38487 9364 38490
rect 9312 38453 9317 38487
rect 9317 38453 9351 38487
rect 9351 38453 9364 38487
rect 9312 38438 9364 38453
rect 9380 38487 9432 38490
rect 9380 38453 9389 38487
rect 9389 38453 9423 38487
rect 9423 38453 9432 38487
rect 9380 38438 9432 38453
rect 9448 38487 9500 38490
rect 9448 38453 9461 38487
rect 9461 38453 9495 38487
rect 9495 38453 9500 38487
rect 9448 38438 9500 38453
rect 9312 38412 9364 38426
rect 9312 38378 9317 38412
rect 9317 38378 9351 38412
rect 9351 38378 9364 38412
rect 9312 38374 9364 38378
rect 9380 38412 9432 38426
rect 9380 38378 9389 38412
rect 9389 38378 9423 38412
rect 9423 38378 9432 38412
rect 9380 38374 9432 38378
rect 9448 38412 9500 38426
rect 9448 38378 9461 38412
rect 9461 38378 9495 38412
rect 9495 38378 9500 38412
rect 9448 38374 9500 38378
rect 9312 38337 9364 38362
rect 9312 38310 9317 38337
rect 9317 38310 9351 38337
rect 9351 38310 9364 38337
rect 9380 38337 9432 38362
rect 9380 38310 9389 38337
rect 9389 38310 9423 38337
rect 9423 38310 9432 38337
rect 9448 38337 9500 38362
rect 9448 38310 9461 38337
rect 9461 38310 9495 38337
rect 9495 38310 9500 38337
rect 9312 38262 9364 38298
rect 9312 38246 9317 38262
rect 9317 38246 9351 38262
rect 9351 38246 9364 38262
rect 9380 38262 9432 38298
rect 9380 38246 9389 38262
rect 9389 38246 9423 38262
rect 9423 38246 9432 38262
rect 9448 38262 9500 38298
rect 9448 38246 9461 38262
rect 9461 38246 9495 38262
rect 9495 38246 9500 38262
rect 9312 38228 9317 38234
rect 9317 38228 9351 38234
rect 9351 38228 9364 38234
rect 9312 38187 9364 38228
rect 9312 38182 9317 38187
rect 9317 38182 9351 38187
rect 9351 38182 9364 38187
rect 9380 38228 9389 38234
rect 9389 38228 9423 38234
rect 9423 38228 9432 38234
rect 9380 38187 9432 38228
rect 9380 38182 9389 38187
rect 9389 38182 9423 38187
rect 9423 38182 9432 38187
rect 9448 38228 9461 38234
rect 9461 38228 9495 38234
rect 9495 38228 9500 38234
rect 9448 38187 9500 38228
rect 9448 38182 9461 38187
rect 9461 38182 9495 38187
rect 9495 38182 9500 38187
rect 9312 38153 9317 38170
rect 9317 38153 9351 38170
rect 9351 38153 9364 38170
rect 9312 38118 9364 38153
rect 9380 38153 9389 38170
rect 9389 38153 9423 38170
rect 9423 38153 9432 38170
rect 9380 38118 9432 38153
rect 9448 38153 9461 38170
rect 9461 38153 9495 38170
rect 9495 38153 9500 38170
rect 9448 38118 9500 38153
rect 10232 39006 10284 39009
rect 10232 38972 10237 39006
rect 10237 38972 10271 39006
rect 10271 38972 10284 39006
rect 10232 38957 10284 38972
rect 10300 39006 10352 39009
rect 10300 38972 10309 39006
rect 10309 38972 10343 39006
rect 10343 38972 10352 39006
rect 10300 38957 10352 38972
rect 10368 39006 10420 39009
rect 10368 38972 10381 39006
rect 10381 38972 10415 39006
rect 10415 38972 10420 39006
rect 10368 38957 10420 38972
rect 10232 38932 10284 38944
rect 10232 38898 10237 38932
rect 10237 38898 10271 38932
rect 10271 38898 10284 38932
rect 10232 38892 10284 38898
rect 10300 38932 10352 38944
rect 10300 38898 10309 38932
rect 10309 38898 10343 38932
rect 10343 38898 10352 38932
rect 10300 38892 10352 38898
rect 10368 38932 10420 38944
rect 10368 38898 10381 38932
rect 10381 38898 10415 38932
rect 10415 38898 10420 38932
rect 10368 38892 10420 38898
rect 10232 38858 10284 38879
rect 10232 38827 10237 38858
rect 10237 38827 10271 38858
rect 10271 38827 10284 38858
rect 10300 38858 10352 38879
rect 10300 38827 10309 38858
rect 10309 38827 10343 38858
rect 10343 38827 10352 38858
rect 10368 38858 10420 38879
rect 10368 38827 10381 38858
rect 10381 38827 10415 38858
rect 10415 38827 10420 38858
rect 10232 38784 10284 38814
rect 10232 38762 10237 38784
rect 10237 38762 10271 38784
rect 10271 38762 10284 38784
rect 10300 38784 10352 38814
rect 10300 38762 10309 38784
rect 10309 38762 10343 38784
rect 10343 38762 10352 38784
rect 10368 38784 10420 38814
rect 10368 38762 10381 38784
rect 10381 38762 10415 38784
rect 10415 38762 10420 38784
rect 10232 38710 10284 38749
rect 10232 38697 10237 38710
rect 10237 38697 10271 38710
rect 10271 38697 10284 38710
rect 10300 38710 10352 38749
rect 10300 38697 10309 38710
rect 10309 38697 10343 38710
rect 10343 38697 10352 38710
rect 10368 38710 10420 38749
rect 10368 38697 10381 38710
rect 10381 38697 10415 38710
rect 10415 38697 10420 38710
rect 10232 38676 10237 38684
rect 10237 38676 10271 38684
rect 10271 38676 10284 38684
rect 10232 38636 10284 38676
rect 10232 38632 10237 38636
rect 10237 38632 10271 38636
rect 10271 38632 10284 38636
rect 10300 38676 10309 38684
rect 10309 38676 10343 38684
rect 10343 38676 10352 38684
rect 10300 38636 10352 38676
rect 10300 38632 10309 38636
rect 10309 38632 10343 38636
rect 10343 38632 10352 38636
rect 10368 38676 10381 38684
rect 10381 38676 10415 38684
rect 10415 38676 10420 38684
rect 10368 38636 10420 38676
rect 10368 38632 10381 38636
rect 10381 38632 10415 38636
rect 10415 38632 10420 38636
rect 10232 38602 10237 38619
rect 10237 38602 10271 38619
rect 10271 38602 10284 38619
rect 10232 38567 10284 38602
rect 10300 38602 10309 38619
rect 10309 38602 10343 38619
rect 10343 38602 10352 38619
rect 10300 38567 10352 38602
rect 10368 38602 10381 38619
rect 10381 38602 10415 38619
rect 10415 38602 10420 38619
rect 10368 38567 10420 38602
rect 10232 38528 10237 38554
rect 10237 38528 10271 38554
rect 10271 38528 10284 38554
rect 10232 38502 10284 38528
rect 10300 38528 10309 38554
rect 10309 38528 10343 38554
rect 10343 38528 10352 38554
rect 10300 38502 10352 38528
rect 10368 38528 10381 38554
rect 10381 38528 10415 38554
rect 10415 38528 10420 38554
rect 10368 38502 10420 38528
rect 10232 38487 10284 38490
rect 10232 38453 10237 38487
rect 10237 38453 10271 38487
rect 10271 38453 10284 38487
rect 10232 38438 10284 38453
rect 10300 38487 10352 38490
rect 10300 38453 10309 38487
rect 10309 38453 10343 38487
rect 10343 38453 10352 38487
rect 10300 38438 10352 38453
rect 10368 38487 10420 38490
rect 10368 38453 10381 38487
rect 10381 38453 10415 38487
rect 10415 38453 10420 38487
rect 10368 38438 10420 38453
rect 10232 38412 10284 38426
rect 10232 38378 10237 38412
rect 10237 38378 10271 38412
rect 10271 38378 10284 38412
rect 10232 38374 10284 38378
rect 10300 38412 10352 38426
rect 10300 38378 10309 38412
rect 10309 38378 10343 38412
rect 10343 38378 10352 38412
rect 10300 38374 10352 38378
rect 10368 38412 10420 38426
rect 10368 38378 10381 38412
rect 10381 38378 10415 38412
rect 10415 38378 10420 38412
rect 10368 38374 10420 38378
rect 10232 38337 10284 38362
rect 10232 38310 10237 38337
rect 10237 38310 10271 38337
rect 10271 38310 10284 38337
rect 10300 38337 10352 38362
rect 10300 38310 10309 38337
rect 10309 38310 10343 38337
rect 10343 38310 10352 38337
rect 10368 38337 10420 38362
rect 10368 38310 10381 38337
rect 10381 38310 10415 38337
rect 10415 38310 10420 38337
rect 10232 38262 10284 38298
rect 10232 38246 10237 38262
rect 10237 38246 10271 38262
rect 10271 38246 10284 38262
rect 10300 38262 10352 38298
rect 10300 38246 10309 38262
rect 10309 38246 10343 38262
rect 10343 38246 10352 38262
rect 10368 38262 10420 38298
rect 10368 38246 10381 38262
rect 10381 38246 10415 38262
rect 10415 38246 10420 38262
rect 10232 38228 10237 38234
rect 10237 38228 10271 38234
rect 10271 38228 10284 38234
rect 10232 38187 10284 38228
rect 10232 38182 10237 38187
rect 10237 38182 10271 38187
rect 10271 38182 10284 38187
rect 10300 38228 10309 38234
rect 10309 38228 10343 38234
rect 10343 38228 10352 38234
rect 10300 38187 10352 38228
rect 10300 38182 10309 38187
rect 10309 38182 10343 38187
rect 10343 38182 10352 38187
rect 10368 38228 10381 38234
rect 10381 38228 10415 38234
rect 10415 38228 10420 38234
rect 10368 38187 10420 38228
rect 10368 38182 10381 38187
rect 10381 38182 10415 38187
rect 10415 38182 10420 38187
rect 10232 38153 10237 38170
rect 10237 38153 10271 38170
rect 10271 38153 10284 38170
rect 10232 38118 10284 38153
rect 10300 38153 10309 38170
rect 10309 38153 10343 38170
rect 10343 38153 10352 38170
rect 10300 38118 10352 38153
rect 10368 38153 10381 38170
rect 10381 38153 10415 38170
rect 10415 38153 10420 38170
rect 10368 38118 10420 38153
rect 11152 38957 11157 39009
rect 11157 38957 11204 39009
rect 11220 38957 11272 39009
rect 11288 38957 11335 39009
rect 11335 38957 11340 39009
rect 11152 38892 11157 38944
rect 11157 38892 11204 38944
rect 11220 38892 11272 38944
rect 11288 38892 11335 38944
rect 11335 38892 11340 38944
rect 11152 38827 11157 38879
rect 11157 38827 11204 38879
rect 11220 38827 11272 38879
rect 11288 38827 11335 38879
rect 11335 38827 11340 38879
rect 11152 38762 11157 38814
rect 11157 38762 11204 38814
rect 11220 38762 11272 38814
rect 11288 38762 11335 38814
rect 11335 38762 11340 38814
rect 11152 38697 11157 38749
rect 11157 38697 11204 38749
rect 11220 38697 11272 38749
rect 11288 38697 11335 38749
rect 11335 38697 11340 38749
rect 11152 38632 11157 38684
rect 11157 38632 11204 38684
rect 11220 38632 11272 38684
rect 11288 38632 11335 38684
rect 11335 38632 11340 38684
rect 11152 38567 11157 38619
rect 11157 38567 11204 38619
rect 11220 38567 11272 38619
rect 11288 38567 11335 38619
rect 11335 38567 11340 38619
rect 11152 38502 11157 38554
rect 11157 38502 11204 38554
rect 11220 38502 11272 38554
rect 11288 38502 11335 38554
rect 11335 38502 11340 38554
rect 11152 38451 11204 38490
rect 11152 38438 11157 38451
rect 11157 38438 11191 38451
rect 11191 38438 11204 38451
rect 11220 38451 11272 38490
rect 11220 38438 11229 38451
rect 11229 38438 11263 38451
rect 11263 38438 11272 38451
rect 11288 38451 11340 38490
rect 11288 38438 11301 38451
rect 11301 38438 11335 38451
rect 11335 38438 11340 38451
rect 11152 38417 11157 38426
rect 11157 38417 11191 38426
rect 11191 38417 11204 38426
rect 11152 38378 11204 38417
rect 11152 38374 11157 38378
rect 11157 38374 11191 38378
rect 11191 38374 11204 38378
rect 11220 38417 11229 38426
rect 11229 38417 11263 38426
rect 11263 38417 11272 38426
rect 11220 38378 11272 38417
rect 11220 38374 11229 38378
rect 11229 38374 11263 38378
rect 11263 38374 11272 38378
rect 11288 38417 11301 38426
rect 11301 38417 11335 38426
rect 11335 38417 11340 38426
rect 11288 38378 11340 38417
rect 11288 38374 11301 38378
rect 11301 38374 11335 38378
rect 11335 38374 11340 38378
rect 11152 38344 11157 38362
rect 11157 38344 11191 38362
rect 11191 38344 11204 38362
rect 11152 38310 11204 38344
rect 11220 38344 11229 38362
rect 11229 38344 11263 38362
rect 11263 38344 11272 38362
rect 11220 38310 11272 38344
rect 11288 38344 11301 38362
rect 11301 38344 11335 38362
rect 11335 38344 11340 38362
rect 11288 38310 11340 38344
rect 11152 38271 11157 38298
rect 11157 38271 11191 38298
rect 11191 38271 11204 38298
rect 11152 38246 11204 38271
rect 11220 38271 11229 38298
rect 11229 38271 11263 38298
rect 11263 38271 11272 38298
rect 11220 38246 11272 38271
rect 11288 38271 11301 38298
rect 11301 38271 11335 38298
rect 11335 38271 11340 38298
rect 11288 38246 11340 38271
rect 11152 38232 11204 38234
rect 11152 38198 11157 38232
rect 11157 38198 11191 38232
rect 11191 38198 11204 38232
rect 11152 38182 11204 38198
rect 11220 38232 11272 38234
rect 11220 38198 11229 38232
rect 11229 38198 11263 38232
rect 11263 38198 11272 38232
rect 11220 38182 11272 38198
rect 11288 38232 11340 38234
rect 11288 38198 11301 38232
rect 11301 38198 11335 38232
rect 11335 38198 11340 38232
rect 11288 38182 11340 38198
rect 11152 38159 11204 38170
rect 11152 38125 11157 38159
rect 11157 38125 11191 38159
rect 11191 38125 11204 38159
rect 11152 38118 11204 38125
rect 11220 38159 11272 38170
rect 11220 38125 11229 38159
rect 11229 38125 11263 38159
rect 11263 38125 11272 38159
rect 11220 38118 11272 38125
rect 11288 38159 11340 38170
rect 11288 38125 11301 38159
rect 11301 38125 11335 38159
rect 11335 38125 11340 38159
rect 11288 38118 11340 38125
rect 3792 36238 3797 36290
rect 3797 36238 3844 36290
rect 3860 36238 3912 36290
rect 3928 36238 3975 36290
rect 3975 36238 3980 36290
rect 3792 36174 3797 36226
rect 3797 36174 3844 36226
rect 3860 36174 3912 36226
rect 3928 36174 3975 36226
rect 3975 36174 3980 36226
rect 3792 36110 3797 36162
rect 3797 36110 3844 36162
rect 3860 36110 3912 36162
rect 3928 36110 3975 36162
rect 3975 36110 3980 36162
rect 3792 36046 3797 36098
rect 3797 36046 3844 36098
rect 3860 36046 3912 36098
rect 3928 36046 3975 36098
rect 3975 36046 3980 36098
rect 3792 35982 3797 36034
rect 3797 35982 3844 36034
rect 3860 35982 3912 36034
rect 3928 35982 3975 36034
rect 3975 35982 3980 36034
rect 3792 35918 3797 35970
rect 3797 35918 3844 35970
rect 3860 35918 3912 35970
rect 3928 35918 3975 35970
rect 3975 35918 3980 35970
rect 3792 35854 3797 35906
rect 3797 35854 3844 35906
rect 3860 35854 3912 35906
rect 3928 35854 3975 35906
rect 3975 35854 3980 35906
rect 3792 35790 3797 35842
rect 3797 35790 3844 35842
rect 3860 35790 3912 35842
rect 3928 35790 3975 35842
rect 3975 35790 3980 35842
rect 3792 35726 3797 35778
rect 3797 35726 3844 35778
rect 3860 35726 3912 35778
rect 3928 35726 3975 35778
rect 3975 35726 3980 35778
rect 3792 35662 3797 35714
rect 3797 35662 3844 35714
rect 3860 35662 3912 35714
rect 3928 35662 3975 35714
rect 3975 35662 3980 35714
rect 3792 35598 3797 35650
rect 3797 35598 3844 35650
rect 3860 35598 3912 35650
rect 3928 35598 3975 35650
rect 3975 35598 3980 35650
rect 3792 35534 3797 35586
rect 3797 35534 3844 35586
rect 3860 35534 3912 35586
rect 3928 35534 3975 35586
rect 3975 35534 3980 35586
rect 3792 35470 3797 35522
rect 3797 35470 3844 35522
rect 3860 35470 3912 35522
rect 3928 35470 3975 35522
rect 3975 35470 3980 35522
rect 3792 35406 3797 35458
rect 3797 35406 3844 35458
rect 3860 35406 3912 35458
rect 3928 35406 3975 35458
rect 3975 35406 3980 35458
rect 3792 35342 3797 35394
rect 3797 35342 3844 35394
rect 3860 35342 3912 35394
rect 3928 35342 3975 35394
rect 3975 35342 3980 35394
rect 3792 35277 3797 35329
rect 3797 35277 3844 35329
rect 3860 35277 3912 35329
rect 3928 35277 3975 35329
rect 3975 35277 3980 35329
rect 3792 35212 3797 35264
rect 3797 35212 3844 35264
rect 3860 35212 3912 35264
rect 3928 35212 3975 35264
rect 3975 35212 3980 35264
rect 3792 35147 3797 35199
rect 3797 35147 3844 35199
rect 3860 35147 3912 35199
rect 3928 35147 3975 35199
rect 3975 35147 3980 35199
rect 3792 35082 3797 35134
rect 3797 35082 3844 35134
rect 3860 35082 3912 35134
rect 3928 35082 3975 35134
rect 3975 35082 3980 35134
rect 3792 35017 3797 35069
rect 3797 35017 3844 35069
rect 3860 35017 3912 35069
rect 3928 35017 3975 35069
rect 3975 35017 3980 35069
rect 3792 34952 3797 35004
rect 3797 34952 3844 35004
rect 3860 34952 3912 35004
rect 3928 34952 3975 35004
rect 3975 34952 3980 35004
rect 3792 34887 3797 34939
rect 3797 34887 3844 34939
rect 3860 34887 3912 34939
rect 3928 34887 3975 34939
rect 3975 34887 3980 34939
rect 3792 34822 3797 34874
rect 3797 34822 3844 34874
rect 3860 34822 3912 34874
rect 3928 34822 3975 34874
rect 3975 34822 3980 34874
rect 3792 34757 3797 34809
rect 3797 34757 3844 34809
rect 3860 34757 3912 34809
rect 3928 34757 3975 34809
rect 3975 34757 3980 34809
rect 3792 34692 3797 34744
rect 3797 34692 3844 34744
rect 3860 34692 3912 34744
rect 3928 34692 3975 34744
rect 3975 34692 3980 34744
rect 3792 34627 3797 34679
rect 3797 34627 3844 34679
rect 3860 34627 3912 34679
rect 3928 34627 3975 34679
rect 3975 34627 3980 34679
rect 3792 34562 3797 34614
rect 3797 34562 3844 34614
rect 3860 34562 3912 34614
rect 3928 34562 3975 34614
rect 3975 34562 3980 34614
rect 3792 31638 3797 31690
rect 3797 31638 3844 31690
rect 3860 31638 3912 31690
rect 3928 31638 3975 31690
rect 3975 31638 3980 31690
rect 3792 31574 3797 31626
rect 3797 31574 3844 31626
rect 3860 31574 3912 31626
rect 3928 31574 3975 31626
rect 3975 31574 3980 31626
rect 3792 31510 3797 31562
rect 3797 31510 3844 31562
rect 3860 31510 3912 31562
rect 3928 31510 3975 31562
rect 3975 31510 3980 31562
rect 3792 31446 3797 31498
rect 3797 31446 3844 31498
rect 3860 31446 3912 31498
rect 3928 31446 3975 31498
rect 3975 31446 3980 31498
rect 3792 31382 3797 31434
rect 3797 31382 3844 31434
rect 3860 31382 3912 31434
rect 3928 31382 3975 31434
rect 3975 31382 3980 31434
rect 3792 31318 3797 31370
rect 3797 31318 3844 31370
rect 3860 31318 3912 31370
rect 3928 31318 3975 31370
rect 3975 31318 3980 31370
rect 3792 31254 3797 31306
rect 3797 31254 3844 31306
rect 3860 31254 3912 31306
rect 3928 31254 3975 31306
rect 3975 31254 3980 31306
rect 3792 31190 3797 31242
rect 3797 31190 3844 31242
rect 3860 31190 3912 31242
rect 3928 31190 3975 31242
rect 3975 31190 3980 31242
rect 3792 31126 3797 31178
rect 3797 31126 3844 31178
rect 3860 31126 3912 31178
rect 3928 31126 3975 31178
rect 3975 31126 3980 31178
rect 3792 31062 3797 31114
rect 3797 31062 3844 31114
rect 3860 31062 3912 31114
rect 3928 31062 3975 31114
rect 3975 31062 3980 31114
rect 3792 30998 3797 31050
rect 3797 30998 3844 31050
rect 3860 30998 3912 31050
rect 3928 30998 3975 31050
rect 3975 30998 3980 31050
rect 3792 30934 3797 30986
rect 3797 30934 3844 30986
rect 3860 30934 3912 30986
rect 3928 30934 3975 30986
rect 3975 30934 3980 30986
rect 3792 30870 3797 30922
rect 3797 30870 3844 30922
rect 3860 30870 3912 30922
rect 3928 30870 3975 30922
rect 3975 30870 3980 30922
rect 3792 30806 3797 30858
rect 3797 30806 3844 30858
rect 3860 30806 3912 30858
rect 3928 30806 3975 30858
rect 3975 30806 3980 30858
rect 3792 30742 3797 30794
rect 3797 30742 3844 30794
rect 3860 30742 3912 30794
rect 3928 30742 3975 30794
rect 3975 30742 3980 30794
rect 3792 30677 3797 30729
rect 3797 30677 3844 30729
rect 3860 30677 3912 30729
rect 3928 30677 3975 30729
rect 3975 30677 3980 30729
rect 3792 30612 3797 30664
rect 3797 30612 3844 30664
rect 3860 30612 3912 30664
rect 3928 30612 3975 30664
rect 3975 30612 3980 30664
rect 3792 30547 3797 30599
rect 3797 30547 3844 30599
rect 3860 30547 3912 30599
rect 3928 30547 3975 30599
rect 3975 30547 3980 30599
rect 3792 30482 3797 30534
rect 3797 30482 3844 30534
rect 3860 30482 3912 30534
rect 3928 30482 3975 30534
rect 3975 30482 3980 30534
rect 3792 30417 3797 30469
rect 3797 30417 3844 30469
rect 3860 30417 3912 30469
rect 3928 30417 3975 30469
rect 3975 30417 3980 30469
rect 3792 30352 3797 30404
rect 3797 30352 3844 30404
rect 3860 30352 3912 30404
rect 3928 30352 3975 30404
rect 3975 30352 3980 30404
rect 3792 30287 3797 30339
rect 3797 30287 3844 30339
rect 3860 30287 3912 30339
rect 3928 30287 3975 30339
rect 3975 30287 3980 30339
rect 3792 30222 3797 30274
rect 3797 30222 3844 30274
rect 3860 30222 3912 30274
rect 3928 30222 3975 30274
rect 3975 30222 3980 30274
rect 3792 30157 3797 30209
rect 3797 30157 3844 30209
rect 3860 30157 3912 30209
rect 3928 30157 3975 30209
rect 3975 30157 3980 30209
rect 3792 30092 3797 30144
rect 3797 30092 3844 30144
rect 3860 30092 3912 30144
rect 3928 30092 3975 30144
rect 3975 30092 3980 30144
rect 3792 30027 3797 30079
rect 3797 30027 3844 30079
rect 3860 30027 3912 30079
rect 3928 30027 3975 30079
rect 3975 30027 3980 30079
rect 3792 29962 3797 30014
rect 3797 29962 3844 30014
rect 3860 29962 3912 30014
rect 3928 29962 3975 30014
rect 3975 29962 3980 30014
rect 4281 37945 4333 37997
rect 4359 37945 4411 37997
rect 4281 37877 4333 37929
rect 4359 37877 4411 37929
rect 4281 37809 4333 37861
rect 4359 37809 4411 37861
rect 4281 37741 4333 37793
rect 4359 37741 4411 37793
rect 4281 37673 4333 37725
rect 4359 37673 4411 37725
rect 4281 37605 4333 37657
rect 4359 37605 4411 37657
rect 4281 37537 4333 37589
rect 4359 37537 4411 37589
rect 4281 37469 4333 37521
rect 4359 37469 4411 37521
rect 4281 37401 4333 37453
rect 4359 37401 4411 37453
rect 4281 37333 4333 37385
rect 4359 37333 4411 37385
rect 4281 37266 4333 37318
rect 4359 37266 4411 37318
rect 4281 37199 4333 37251
rect 4359 37199 4411 37251
rect 4281 37132 4333 37184
rect 4359 37132 4411 37184
rect 4281 37065 4333 37117
rect 4359 37065 4411 37117
rect 4281 34173 4333 34225
rect 4359 34173 4411 34225
rect 4281 34109 4333 34161
rect 4359 34109 4411 34161
rect 4281 34045 4333 34097
rect 4359 34045 4411 34097
rect 4281 33981 4333 34033
rect 4359 33981 4411 34033
rect 4281 33917 4333 33969
rect 4359 33917 4411 33969
rect 4281 33853 4333 33905
rect 4359 33853 4411 33905
rect 4281 33789 4333 33841
rect 4359 33789 4411 33841
rect 4281 33725 4333 33777
rect 4359 33725 4411 33777
rect 4281 33661 4333 33713
rect 4359 33661 4411 33713
rect 4281 33597 4333 33649
rect 4359 33597 4411 33649
rect 4281 33533 4333 33585
rect 4359 33533 4411 33585
rect 4281 33469 4333 33521
rect 4359 33469 4411 33521
rect 4281 33405 4333 33457
rect 4359 33405 4411 33457
rect 4281 33341 4333 33393
rect 4359 33341 4411 33393
rect 4281 33277 4333 33329
rect 4359 33277 4411 33329
rect 4281 33212 4333 33264
rect 4359 33212 4411 33264
rect 4281 33147 4333 33199
rect 4359 33147 4411 33199
rect 4281 33082 4333 33134
rect 4359 33082 4411 33134
rect 4281 33017 4333 33069
rect 4359 33017 4411 33069
rect 4281 32952 4333 33004
rect 4359 32952 4411 33004
rect 4281 32887 4333 32939
rect 4359 32887 4411 32939
rect 4281 32822 4333 32874
rect 4359 32822 4411 32874
rect 4281 32757 4333 32809
rect 4359 32757 4411 32809
rect 4281 32692 4333 32744
rect 4359 32692 4411 32744
rect 4281 32627 4333 32679
rect 4359 32627 4411 32679
rect 4281 32562 4333 32614
rect 4359 32562 4411 32614
rect 4281 32497 4333 32549
rect 4359 32497 4411 32549
rect 4281 29573 4333 29625
rect 4359 29573 4411 29625
rect 4281 29509 4333 29561
rect 4359 29509 4411 29561
rect 4281 29445 4333 29497
rect 4359 29445 4411 29497
rect 4281 29381 4333 29433
rect 4359 29381 4411 29433
rect 4281 29317 4333 29369
rect 4359 29317 4411 29369
rect 4281 29253 4333 29305
rect 4359 29253 4411 29305
rect 4281 29189 4333 29241
rect 4359 29189 4411 29241
rect 4281 29125 4333 29177
rect 4359 29125 4411 29177
rect 4281 29061 4333 29113
rect 4359 29061 4411 29113
rect 4281 28997 4333 29049
rect 4359 28997 4411 29049
rect 4281 28933 4333 28985
rect 4359 28933 4411 28985
rect 4281 28869 4333 28921
rect 4359 28869 4411 28921
rect 4281 28805 4333 28857
rect 4359 28805 4411 28857
rect 4281 28741 4333 28793
rect 4359 28741 4411 28793
rect 4281 28677 4333 28729
rect 4359 28677 4411 28729
rect 4281 28612 4333 28664
rect 4359 28612 4411 28664
rect 4281 28547 4333 28599
rect 4359 28547 4411 28599
rect 4281 28482 4333 28534
rect 4359 28482 4411 28534
rect 4281 28417 4333 28469
rect 4359 28417 4411 28469
rect 4281 28352 4333 28404
rect 4359 28352 4411 28404
rect 4281 28287 4333 28339
rect 4359 28287 4411 28339
rect 4281 28222 4333 28274
rect 4359 28222 4411 28274
rect 4281 28157 4333 28209
rect 4359 28157 4411 28209
rect 4281 28092 4333 28144
rect 4359 28092 4411 28144
rect 4281 28027 4333 28079
rect 4359 28027 4411 28079
rect 4281 27962 4333 28014
rect 4359 27962 4411 28014
rect 4281 27897 4333 27949
rect 4359 27897 4411 27949
rect 4712 36238 4717 36290
rect 4717 36238 4764 36290
rect 4780 36238 4832 36290
rect 4848 36238 4895 36290
rect 4895 36238 4900 36290
rect 4712 36174 4717 36226
rect 4717 36174 4764 36226
rect 4780 36174 4832 36226
rect 4848 36174 4895 36226
rect 4895 36174 4900 36226
rect 4712 36110 4717 36162
rect 4717 36110 4764 36162
rect 4780 36110 4832 36162
rect 4848 36110 4895 36162
rect 4895 36110 4900 36162
rect 4712 36046 4717 36098
rect 4717 36046 4764 36098
rect 4780 36046 4832 36098
rect 4848 36046 4895 36098
rect 4895 36046 4900 36098
rect 4712 35982 4717 36034
rect 4717 35982 4764 36034
rect 4780 35982 4832 36034
rect 4848 35982 4895 36034
rect 4895 35982 4900 36034
rect 4712 35918 4717 35970
rect 4717 35918 4764 35970
rect 4780 35918 4832 35970
rect 4848 35918 4895 35970
rect 4895 35918 4900 35970
rect 4712 35854 4717 35906
rect 4717 35854 4764 35906
rect 4780 35854 4832 35906
rect 4848 35854 4895 35906
rect 4895 35854 4900 35906
rect 4712 35790 4717 35842
rect 4717 35790 4764 35842
rect 4780 35790 4832 35842
rect 4848 35790 4895 35842
rect 4895 35790 4900 35842
rect 4712 35726 4717 35778
rect 4717 35726 4764 35778
rect 4780 35726 4832 35778
rect 4848 35726 4895 35778
rect 4895 35726 4900 35778
rect 4712 35662 4717 35714
rect 4717 35662 4764 35714
rect 4780 35662 4832 35714
rect 4848 35662 4895 35714
rect 4895 35662 4900 35714
rect 4712 35598 4717 35650
rect 4717 35598 4764 35650
rect 4780 35598 4832 35650
rect 4848 35598 4895 35650
rect 4895 35598 4900 35650
rect 4712 35534 4717 35586
rect 4717 35534 4764 35586
rect 4780 35534 4832 35586
rect 4848 35534 4895 35586
rect 4895 35534 4900 35586
rect 4712 35470 4717 35522
rect 4717 35470 4764 35522
rect 4780 35470 4832 35522
rect 4848 35470 4895 35522
rect 4895 35470 4900 35522
rect 4712 35406 4717 35458
rect 4717 35406 4764 35458
rect 4780 35406 4832 35458
rect 4848 35406 4895 35458
rect 4895 35406 4900 35458
rect 4712 35342 4717 35394
rect 4717 35342 4764 35394
rect 4780 35342 4832 35394
rect 4848 35342 4895 35394
rect 4895 35342 4900 35394
rect 4712 35277 4717 35329
rect 4717 35277 4764 35329
rect 4780 35277 4832 35329
rect 4848 35277 4895 35329
rect 4895 35277 4900 35329
rect 4712 35212 4717 35264
rect 4717 35212 4764 35264
rect 4780 35212 4832 35264
rect 4848 35212 4895 35264
rect 4895 35212 4900 35264
rect 4712 35147 4717 35199
rect 4717 35147 4764 35199
rect 4780 35147 4832 35199
rect 4848 35147 4895 35199
rect 4895 35147 4900 35199
rect 4712 35082 4717 35134
rect 4717 35082 4764 35134
rect 4780 35082 4832 35134
rect 4848 35082 4895 35134
rect 4895 35082 4900 35134
rect 4712 35017 4717 35069
rect 4717 35017 4764 35069
rect 4780 35017 4832 35069
rect 4848 35017 4895 35069
rect 4895 35017 4900 35069
rect 4712 34952 4717 35004
rect 4717 34952 4764 35004
rect 4780 34952 4832 35004
rect 4848 34952 4895 35004
rect 4895 34952 4900 35004
rect 4712 34887 4717 34939
rect 4717 34887 4764 34939
rect 4780 34887 4832 34939
rect 4848 34887 4895 34939
rect 4895 34887 4900 34939
rect 4712 34822 4717 34874
rect 4717 34822 4764 34874
rect 4780 34822 4832 34874
rect 4848 34822 4895 34874
rect 4895 34822 4900 34874
rect 4712 34757 4717 34809
rect 4717 34757 4764 34809
rect 4780 34757 4832 34809
rect 4848 34757 4895 34809
rect 4895 34757 4900 34809
rect 4712 34692 4717 34744
rect 4717 34692 4764 34744
rect 4780 34692 4832 34744
rect 4848 34692 4895 34744
rect 4895 34692 4900 34744
rect 4712 34627 4717 34679
rect 4717 34627 4764 34679
rect 4780 34627 4832 34679
rect 4848 34627 4895 34679
rect 4895 34627 4900 34679
rect 4712 34562 4717 34614
rect 4717 34562 4764 34614
rect 4780 34562 4832 34614
rect 4848 34562 4895 34614
rect 4895 34562 4900 34614
rect 4712 31638 4717 31690
rect 4717 31638 4764 31690
rect 4780 31638 4832 31690
rect 4848 31638 4895 31690
rect 4895 31638 4900 31690
rect 4712 31574 4717 31626
rect 4717 31574 4764 31626
rect 4780 31574 4832 31626
rect 4848 31574 4895 31626
rect 4895 31574 4900 31626
rect 4712 31510 4717 31562
rect 4717 31510 4764 31562
rect 4780 31510 4832 31562
rect 4848 31510 4895 31562
rect 4895 31510 4900 31562
rect 4712 31446 4717 31498
rect 4717 31446 4764 31498
rect 4780 31446 4832 31498
rect 4848 31446 4895 31498
rect 4895 31446 4900 31498
rect 4712 31382 4717 31434
rect 4717 31382 4764 31434
rect 4780 31382 4832 31434
rect 4848 31382 4895 31434
rect 4895 31382 4900 31434
rect 4712 31318 4717 31370
rect 4717 31318 4764 31370
rect 4780 31318 4832 31370
rect 4848 31318 4895 31370
rect 4895 31318 4900 31370
rect 4712 31254 4717 31306
rect 4717 31254 4764 31306
rect 4780 31254 4832 31306
rect 4848 31254 4895 31306
rect 4895 31254 4900 31306
rect 4712 31190 4717 31242
rect 4717 31190 4764 31242
rect 4780 31190 4832 31242
rect 4848 31190 4895 31242
rect 4895 31190 4900 31242
rect 4712 31126 4717 31178
rect 4717 31126 4764 31178
rect 4780 31126 4832 31178
rect 4848 31126 4895 31178
rect 4895 31126 4900 31178
rect 4712 31062 4717 31114
rect 4717 31062 4764 31114
rect 4780 31062 4832 31114
rect 4848 31062 4895 31114
rect 4895 31062 4900 31114
rect 4712 30998 4717 31050
rect 4717 30998 4764 31050
rect 4780 30998 4832 31050
rect 4848 30998 4895 31050
rect 4895 30998 4900 31050
rect 4712 30934 4717 30986
rect 4717 30934 4764 30986
rect 4780 30934 4832 30986
rect 4848 30934 4895 30986
rect 4895 30934 4900 30986
rect 4712 30870 4717 30922
rect 4717 30870 4764 30922
rect 4780 30870 4832 30922
rect 4848 30870 4895 30922
rect 4895 30870 4900 30922
rect 4712 30806 4717 30858
rect 4717 30806 4764 30858
rect 4780 30806 4832 30858
rect 4848 30806 4895 30858
rect 4895 30806 4900 30858
rect 4712 30742 4717 30794
rect 4717 30742 4764 30794
rect 4780 30742 4832 30794
rect 4848 30742 4895 30794
rect 4895 30742 4900 30794
rect 4712 30677 4717 30729
rect 4717 30677 4764 30729
rect 4780 30677 4832 30729
rect 4848 30677 4895 30729
rect 4895 30677 4900 30729
rect 4712 30612 4717 30664
rect 4717 30612 4764 30664
rect 4780 30612 4832 30664
rect 4848 30612 4895 30664
rect 4895 30612 4900 30664
rect 4712 30547 4717 30599
rect 4717 30547 4764 30599
rect 4780 30547 4832 30599
rect 4848 30547 4895 30599
rect 4895 30547 4900 30599
rect 4712 30482 4717 30534
rect 4717 30482 4764 30534
rect 4780 30482 4832 30534
rect 4848 30482 4895 30534
rect 4895 30482 4900 30534
rect 4712 30417 4717 30469
rect 4717 30417 4764 30469
rect 4780 30417 4832 30469
rect 4848 30417 4895 30469
rect 4895 30417 4900 30469
rect 4712 30352 4717 30404
rect 4717 30352 4764 30404
rect 4780 30352 4832 30404
rect 4848 30352 4895 30404
rect 4895 30352 4900 30404
rect 4712 30287 4717 30339
rect 4717 30287 4764 30339
rect 4780 30287 4832 30339
rect 4848 30287 4895 30339
rect 4895 30287 4900 30339
rect 4712 30222 4717 30274
rect 4717 30222 4764 30274
rect 4780 30222 4832 30274
rect 4848 30222 4895 30274
rect 4895 30222 4900 30274
rect 4712 30157 4717 30209
rect 4717 30157 4764 30209
rect 4780 30157 4832 30209
rect 4848 30157 4895 30209
rect 4895 30157 4900 30209
rect 4712 30092 4717 30144
rect 4717 30092 4764 30144
rect 4780 30092 4832 30144
rect 4848 30092 4895 30144
rect 4895 30092 4900 30144
rect 4712 30027 4717 30079
rect 4717 30027 4764 30079
rect 4780 30027 4832 30079
rect 4848 30027 4895 30079
rect 4895 30027 4900 30079
rect 4712 29962 4717 30014
rect 4717 29962 4764 30014
rect 4780 29962 4832 30014
rect 4848 29962 4895 30014
rect 4895 29962 4900 30014
rect 3456 23380 3508 23432
rect 3456 23305 3508 23357
rect 3456 23230 3508 23282
rect 4780 27089 4832 27090
rect 4780 27055 4783 27089
rect 4783 27055 4817 27089
rect 4817 27055 4832 27089
rect 4780 27038 4832 27055
rect 4848 27089 4900 27090
rect 4848 27055 4861 27089
rect 4861 27055 4895 27089
rect 4895 27055 4900 27089
rect 4848 27038 4900 27055
rect 4780 27016 4832 27026
rect 4780 26982 4783 27016
rect 4783 26982 4817 27016
rect 4817 26982 4832 27016
rect 4780 26974 4832 26982
rect 4848 27016 4900 27026
rect 4848 26982 4861 27016
rect 4861 26982 4895 27016
rect 4895 26982 4900 27016
rect 4848 26974 4900 26982
rect 4780 26943 4832 26962
rect 4780 26910 4783 26943
rect 4783 26910 4817 26943
rect 4817 26910 4832 26943
rect 4848 26943 4900 26962
rect 4848 26910 4861 26943
rect 4861 26910 4895 26943
rect 4895 26910 4900 26943
rect 4780 26870 4832 26898
rect 4780 26846 4783 26870
rect 4783 26846 4817 26870
rect 4817 26846 4832 26870
rect 4848 26870 4900 26898
rect 4848 26846 4861 26870
rect 4861 26846 4895 26870
rect 4895 26846 4900 26870
rect 4780 26797 4832 26834
rect 4780 26782 4783 26797
rect 4783 26782 4817 26797
rect 4817 26782 4832 26797
rect 4848 26797 4900 26834
rect 4848 26782 4861 26797
rect 4861 26782 4895 26797
rect 4895 26782 4900 26797
rect 4780 26763 4783 26770
rect 4783 26763 4817 26770
rect 4817 26763 4832 26770
rect 4780 26724 4832 26763
rect 4780 26718 4783 26724
rect 4783 26718 4817 26724
rect 4817 26718 4832 26724
rect 4848 26763 4861 26770
rect 4861 26763 4895 26770
rect 4895 26763 4900 26770
rect 4848 26724 4900 26763
rect 4848 26718 4861 26724
rect 4861 26718 4895 26724
rect 4895 26718 4900 26724
rect 4780 26690 4783 26706
rect 4783 26690 4817 26706
rect 4817 26690 4832 26706
rect 4780 26654 4832 26690
rect 4848 26690 4861 26706
rect 4861 26690 4895 26706
rect 4895 26690 4900 26706
rect 4848 26654 4900 26690
rect 4780 26617 4783 26642
rect 4783 26617 4817 26642
rect 4817 26617 4832 26642
rect 4780 26590 4832 26617
rect 4848 26617 4861 26642
rect 4861 26617 4895 26642
rect 4895 26617 4900 26642
rect 4848 26590 4900 26617
rect 4780 26544 4783 26578
rect 4783 26544 4817 26578
rect 4817 26544 4832 26578
rect 4780 26526 4832 26544
rect 4848 26544 4861 26578
rect 4861 26544 4895 26578
rect 4895 26544 4900 26578
rect 4848 26526 4900 26544
rect 4780 26505 4832 26514
rect 4780 26471 4783 26505
rect 4783 26471 4817 26505
rect 4817 26471 4832 26505
rect 4780 26462 4832 26471
rect 4848 26505 4900 26514
rect 4848 26471 4861 26505
rect 4861 26471 4895 26505
rect 4895 26471 4900 26505
rect 4848 26462 4900 26471
rect 4780 26432 4832 26450
rect 4780 26398 4783 26432
rect 4783 26398 4817 26432
rect 4817 26398 4832 26432
rect 4848 26432 4900 26450
rect 4848 26398 4861 26432
rect 4861 26398 4895 26432
rect 4895 26398 4900 26432
rect 4780 26359 4832 26386
rect 4780 26334 4783 26359
rect 4783 26334 4817 26359
rect 4817 26334 4832 26359
rect 4848 26359 4900 26386
rect 4848 26334 4861 26359
rect 4861 26334 4895 26359
rect 4895 26334 4900 26359
rect 4780 26286 4832 26322
rect 4780 26270 4783 26286
rect 4783 26270 4817 26286
rect 4817 26270 4832 26286
rect 4848 26286 4900 26322
rect 4848 26270 4861 26286
rect 4861 26270 4895 26286
rect 4895 26270 4900 26286
rect 4780 26252 4783 26258
rect 4783 26252 4817 26258
rect 4817 26252 4832 26258
rect 4780 26213 4832 26252
rect 4780 26206 4783 26213
rect 4783 26206 4817 26213
rect 4817 26206 4832 26213
rect 4848 26252 4861 26258
rect 4861 26252 4895 26258
rect 4895 26252 4900 26258
rect 4848 26213 4900 26252
rect 4848 26206 4861 26213
rect 4861 26206 4895 26213
rect 4895 26206 4900 26213
rect 4780 26179 4783 26194
rect 4783 26179 4817 26194
rect 4817 26179 4832 26194
rect 4780 26142 4832 26179
rect 4848 26179 4861 26194
rect 4861 26179 4895 26194
rect 4895 26179 4900 26194
rect 4848 26142 4900 26179
rect 4780 26106 4783 26129
rect 4783 26106 4817 26129
rect 4817 26106 4832 26129
rect 4780 26077 4832 26106
rect 4848 26106 4861 26129
rect 4861 26106 4895 26129
rect 4895 26106 4900 26129
rect 4848 26077 4900 26106
rect 4780 26033 4783 26064
rect 4783 26033 4817 26064
rect 4817 26033 4832 26064
rect 4780 26012 4832 26033
rect 4848 26033 4861 26064
rect 4861 26033 4895 26064
rect 4895 26033 4900 26064
rect 4848 26012 4900 26033
rect 4780 25994 4832 25999
rect 4780 25960 4783 25994
rect 4783 25960 4817 25994
rect 4817 25960 4832 25994
rect 4780 25947 4832 25960
rect 4848 25994 4900 25999
rect 4848 25960 4861 25994
rect 4861 25960 4895 25994
rect 4895 25960 4900 25994
rect 4848 25947 4900 25960
rect 4780 25921 4832 25934
rect 4780 25887 4783 25921
rect 4783 25887 4817 25921
rect 4817 25887 4832 25921
rect 4780 25882 4832 25887
rect 4848 25921 4900 25934
rect 4848 25887 4861 25921
rect 4861 25887 4895 25921
rect 4895 25887 4900 25921
rect 4848 25882 4900 25887
rect 4780 25848 4832 25869
rect 4780 25817 4783 25848
rect 4783 25817 4817 25848
rect 4817 25817 4832 25848
rect 4848 25848 4900 25869
rect 4848 25817 4861 25848
rect 4861 25817 4895 25848
rect 4895 25817 4900 25848
rect 4780 25775 4832 25804
rect 4780 25752 4783 25775
rect 4783 25752 4817 25775
rect 4817 25752 4832 25775
rect 4848 25775 4900 25804
rect 4848 25752 4861 25775
rect 4861 25752 4895 25775
rect 4895 25752 4900 25775
rect 4780 25702 4832 25739
rect 4780 25687 4783 25702
rect 4783 25687 4817 25702
rect 4817 25687 4832 25702
rect 4848 25702 4900 25739
rect 4848 25687 4861 25702
rect 4861 25687 4895 25702
rect 4895 25687 4900 25702
rect 4780 25668 4783 25674
rect 4783 25668 4817 25674
rect 4817 25668 4832 25674
rect 4780 25629 4832 25668
rect 4780 25622 4783 25629
rect 4783 25622 4817 25629
rect 4817 25622 4832 25629
rect 4848 25668 4861 25674
rect 4861 25668 4895 25674
rect 4895 25668 4900 25674
rect 4848 25629 4900 25668
rect 4848 25622 4861 25629
rect 4861 25622 4895 25629
rect 4895 25622 4900 25629
rect 4780 25595 4783 25609
rect 4783 25595 4817 25609
rect 4817 25595 4832 25609
rect 4780 25557 4832 25595
rect 4848 25595 4861 25609
rect 4861 25595 4895 25609
rect 4895 25595 4900 25609
rect 4848 25557 4900 25595
rect 4780 25522 4783 25544
rect 4783 25522 4817 25544
rect 4817 25522 4832 25544
rect 4780 25492 4832 25522
rect 4848 25522 4861 25544
rect 4861 25522 4895 25544
rect 4895 25522 4900 25544
rect 4848 25492 4900 25522
rect 4780 25449 4783 25479
rect 4783 25449 4817 25479
rect 4817 25449 4832 25479
rect 4780 25427 4832 25449
rect 4848 25449 4861 25479
rect 4861 25449 4895 25479
rect 4895 25449 4900 25479
rect 4848 25427 4900 25449
rect 4780 25410 4832 25414
rect 4780 25376 4783 25410
rect 4783 25376 4817 25410
rect 4817 25376 4832 25410
rect 4780 25362 4832 25376
rect 4848 25410 4900 25414
rect 4848 25376 4861 25410
rect 4861 25376 4895 25410
rect 4895 25376 4900 25410
rect 4848 25362 4900 25376
rect 5201 37945 5253 37997
rect 5279 37945 5331 37997
rect 5201 37877 5253 37929
rect 5279 37877 5331 37929
rect 5201 37809 5253 37861
rect 5279 37809 5331 37861
rect 5201 37741 5253 37793
rect 5279 37741 5331 37793
rect 5201 37673 5253 37725
rect 5279 37673 5331 37725
rect 5201 37605 5253 37657
rect 5279 37605 5331 37657
rect 5201 37537 5253 37589
rect 5279 37537 5331 37589
rect 5201 37469 5253 37521
rect 5279 37469 5331 37521
rect 5201 37401 5253 37453
rect 5279 37401 5331 37453
rect 5201 37333 5253 37385
rect 5279 37333 5331 37385
rect 5201 37266 5253 37318
rect 5279 37266 5331 37318
rect 5201 37199 5253 37251
rect 5279 37199 5331 37251
rect 5201 37132 5253 37184
rect 5279 37132 5331 37184
rect 5201 37065 5253 37117
rect 5279 37065 5331 37117
rect 5201 34173 5253 34225
rect 5279 34173 5331 34225
rect 5201 34109 5253 34161
rect 5279 34109 5331 34161
rect 5201 34045 5253 34097
rect 5279 34045 5331 34097
rect 5201 33981 5253 34033
rect 5279 33981 5331 34033
rect 5201 33917 5253 33969
rect 5279 33917 5331 33969
rect 5201 33853 5253 33905
rect 5279 33853 5331 33905
rect 5201 33789 5253 33841
rect 5279 33789 5331 33841
rect 5201 33725 5253 33777
rect 5279 33725 5331 33777
rect 5201 33661 5253 33713
rect 5279 33661 5331 33713
rect 5201 33597 5253 33649
rect 5279 33597 5331 33649
rect 5201 33533 5253 33585
rect 5279 33533 5331 33585
rect 5201 33469 5253 33521
rect 5279 33469 5331 33521
rect 5201 33405 5253 33457
rect 5279 33405 5331 33457
rect 5201 33341 5253 33393
rect 5279 33341 5331 33393
rect 5201 33277 5253 33329
rect 5279 33277 5331 33329
rect 5201 33212 5253 33264
rect 5279 33212 5331 33264
rect 5201 33147 5253 33199
rect 5279 33147 5331 33199
rect 5201 33082 5253 33134
rect 5279 33082 5331 33134
rect 5201 33017 5253 33069
rect 5279 33017 5331 33069
rect 5201 32952 5253 33004
rect 5279 32952 5331 33004
rect 5201 32887 5253 32939
rect 5279 32887 5331 32939
rect 5201 32822 5253 32874
rect 5279 32822 5331 32874
rect 5201 32757 5253 32809
rect 5279 32757 5331 32809
rect 5201 32692 5253 32744
rect 5279 32692 5331 32744
rect 5201 32627 5253 32679
rect 5279 32627 5331 32679
rect 5201 32562 5253 32614
rect 5279 32562 5331 32614
rect 5201 32497 5253 32549
rect 5279 32497 5331 32549
rect 5201 29573 5253 29625
rect 5279 29573 5331 29625
rect 5201 29509 5253 29561
rect 5279 29509 5331 29561
rect 5201 29445 5253 29497
rect 5279 29445 5331 29497
rect 5201 29381 5253 29433
rect 5279 29381 5331 29433
rect 5201 29317 5253 29369
rect 5279 29317 5331 29369
rect 5201 29253 5253 29305
rect 5279 29253 5331 29305
rect 5201 29189 5253 29241
rect 5279 29189 5331 29241
rect 5201 29125 5253 29177
rect 5279 29125 5331 29177
rect 5201 29061 5253 29113
rect 5279 29061 5331 29113
rect 5201 28997 5253 29049
rect 5279 28997 5331 29049
rect 5201 28933 5253 28985
rect 5279 28933 5331 28985
rect 5201 28869 5253 28921
rect 5279 28869 5331 28921
rect 5201 28805 5253 28857
rect 5279 28805 5331 28857
rect 5201 28741 5253 28793
rect 5279 28741 5331 28793
rect 5201 28677 5253 28729
rect 5279 28677 5331 28729
rect 5201 28612 5253 28664
rect 5279 28612 5331 28664
rect 5201 28547 5253 28599
rect 5279 28547 5331 28599
rect 5201 28482 5253 28534
rect 5279 28482 5331 28534
rect 5201 28417 5253 28469
rect 5279 28417 5331 28469
rect 5201 28352 5253 28404
rect 5279 28352 5331 28404
rect 5201 28287 5253 28339
rect 5279 28287 5331 28339
rect 5201 28222 5253 28274
rect 5279 28222 5331 28274
rect 5201 28157 5253 28209
rect 5279 28157 5331 28209
rect 5201 28092 5253 28144
rect 5279 28092 5331 28144
rect 5201 28027 5253 28079
rect 5279 28027 5331 28079
rect 5201 27962 5253 28014
rect 5279 27962 5331 28014
rect 5201 27897 5253 27949
rect 5279 27897 5331 27949
rect 5201 24973 5253 25025
rect 5279 24973 5331 25025
rect 5201 24909 5253 24961
rect 5279 24909 5331 24961
rect 5201 24845 5253 24897
rect 5279 24845 5331 24897
rect 5201 24781 5253 24833
rect 5279 24781 5331 24833
rect 5201 24717 5253 24769
rect 5279 24717 5331 24769
rect 5201 24653 5253 24705
rect 5279 24653 5331 24705
rect 5201 24589 5253 24641
rect 5279 24589 5331 24641
rect 5201 24525 5253 24577
rect 5279 24525 5331 24577
rect 5201 24461 5253 24513
rect 5279 24461 5331 24513
rect 5201 24397 5253 24449
rect 5279 24397 5331 24449
rect 5201 24333 5253 24385
rect 5279 24333 5331 24385
rect 5201 24269 5253 24321
rect 5279 24269 5331 24321
rect 5201 24205 5253 24257
rect 5279 24205 5331 24257
rect 5201 24141 5253 24193
rect 5279 24141 5331 24193
rect 5201 24077 5253 24129
rect 5279 24077 5331 24129
rect 5201 24012 5253 24064
rect 5279 24012 5331 24064
rect 5201 23947 5253 23999
rect 5279 23947 5331 23999
rect 5201 23882 5253 23934
rect 5279 23882 5331 23934
rect 5201 23817 5253 23869
rect 5279 23817 5331 23869
rect 5201 23752 5253 23804
rect 5279 23752 5331 23804
rect 5201 23687 5253 23739
rect 5279 23687 5331 23739
rect 5201 23622 5253 23674
rect 5279 23622 5331 23674
rect 5201 23557 5253 23609
rect 5279 23557 5331 23609
rect 5201 23492 5253 23544
rect 5279 23492 5331 23544
rect 5201 23427 5253 23479
rect 5279 23427 5331 23479
rect 5201 23362 5253 23414
rect 5279 23362 5331 23414
rect 5201 23297 5253 23349
rect 5279 23297 5331 23349
rect 4783 22993 4835 22995
rect 4783 22959 4789 22993
rect 4789 22959 4823 22993
rect 4823 22959 4835 22993
rect 4783 22943 4835 22959
rect 4783 22921 4835 22931
rect 4783 22887 4789 22921
rect 4789 22887 4823 22921
rect 4823 22887 4835 22921
rect 4783 22879 4835 22887
rect 4777 22484 4829 22490
rect 4849 22484 4901 22490
rect 4777 22438 4784 22484
rect 4784 22438 4829 22484
rect 4849 22438 4890 22484
rect 4890 22438 4901 22484
rect 4777 22374 4784 22426
rect 4784 22374 4829 22426
rect 4849 22374 4890 22426
rect 4890 22374 4901 22426
rect 4777 22310 4784 22362
rect 4784 22310 4829 22362
rect 4849 22310 4890 22362
rect 4890 22310 4901 22362
rect 4777 22246 4784 22298
rect 4784 22246 4829 22298
rect 4849 22246 4890 22298
rect 4890 22246 4901 22298
rect 4777 22182 4784 22234
rect 4784 22182 4829 22234
rect 4849 22182 4890 22234
rect 4890 22182 4901 22234
rect 4777 22118 4784 22170
rect 4784 22118 4829 22170
rect 4849 22118 4890 22170
rect 4890 22118 4901 22170
rect 4777 22054 4784 22106
rect 4784 22054 4829 22106
rect 4849 22054 4890 22106
rect 4890 22054 4901 22106
rect 4777 21990 4784 22042
rect 4784 21990 4829 22042
rect 4849 21990 4890 22042
rect 4890 21990 4901 22042
rect 4777 21926 4784 21978
rect 4784 21926 4829 21978
rect 4849 21926 4890 21978
rect 4890 21926 4901 21978
rect 4777 21862 4784 21914
rect 4784 21862 4829 21914
rect 4849 21862 4890 21914
rect 4890 21862 4901 21914
rect 4777 21798 4784 21850
rect 4784 21798 4829 21850
rect 4849 21798 4890 21850
rect 4890 21798 4901 21850
rect 4777 21734 4784 21786
rect 4784 21734 4829 21786
rect 4849 21734 4890 21786
rect 4890 21734 4901 21786
rect 4777 21670 4784 21722
rect 4784 21670 4829 21722
rect 4849 21670 4890 21722
rect 4890 21670 4901 21722
rect 4777 21606 4784 21658
rect 4784 21606 4829 21658
rect 4849 21606 4890 21658
rect 4890 21606 4901 21658
rect 4777 21542 4784 21594
rect 4784 21542 4829 21594
rect 4849 21542 4890 21594
rect 4890 21542 4901 21594
rect 4777 21477 4784 21529
rect 4784 21477 4829 21529
rect 4849 21477 4890 21529
rect 4890 21477 4901 21529
rect 4777 21412 4784 21464
rect 4784 21412 4829 21464
rect 4849 21412 4890 21464
rect 4890 21412 4901 21464
rect 4777 21347 4784 21399
rect 4784 21347 4829 21399
rect 4849 21347 4890 21399
rect 4890 21347 4901 21399
rect 4777 21282 4784 21334
rect 4784 21282 4829 21334
rect 4849 21282 4890 21334
rect 4890 21282 4901 21334
rect 4777 21217 4784 21269
rect 4784 21217 4829 21269
rect 4849 21217 4890 21269
rect 4890 21217 4901 21269
rect 4777 21152 4784 21204
rect 4784 21152 4829 21204
rect 4849 21152 4890 21204
rect 4890 21152 4901 21204
rect 4777 21087 4784 21139
rect 4784 21087 4829 21139
rect 4849 21087 4890 21139
rect 4890 21087 4901 21139
rect 4777 21022 4784 21074
rect 4784 21022 4829 21074
rect 4849 21022 4890 21074
rect 4890 21022 4901 21074
rect 4777 20957 4784 21009
rect 4784 20957 4829 21009
rect 4849 20957 4890 21009
rect 4890 20957 4901 21009
rect 4777 20892 4784 20944
rect 4784 20892 4829 20944
rect 4849 20892 4890 20944
rect 4890 20892 4901 20944
rect 4777 20827 4784 20879
rect 4784 20827 4829 20879
rect 4849 20827 4890 20879
rect 4890 20827 4901 20879
rect 4777 20762 4784 20814
rect 4784 20762 4829 20814
rect 4849 20762 4890 20814
rect 4890 20762 4901 20814
rect 3688 14874 3740 14883
rect 3688 14840 3694 14874
rect 3694 14840 3728 14874
rect 3728 14840 3740 14874
rect 3688 14831 3740 14840
rect 3754 14874 3806 14883
rect 3754 14840 3766 14874
rect 3766 14840 3800 14874
rect 3800 14840 3806 14874
rect 3754 14831 3806 14840
rect 3359 14650 3411 14702
rect 3448 14650 3500 14702
rect 3367 13642 3419 13651
rect 3456 13642 3508 13651
rect 3367 13608 3376 13642
rect 3376 13608 3410 13642
rect 3410 13608 3419 13642
rect 3456 13608 3483 13642
rect 3483 13608 3508 13642
rect 3367 13599 3419 13608
rect 3456 13599 3508 13608
rect 4712 17838 4717 17890
rect 4717 17838 4764 17890
rect 4780 17838 4832 17890
rect 4848 17838 4895 17890
rect 4895 17838 4900 17890
rect 4712 17774 4717 17826
rect 4717 17774 4764 17826
rect 4780 17774 4832 17826
rect 4848 17774 4895 17826
rect 4895 17774 4900 17826
rect 4712 17710 4717 17762
rect 4717 17710 4764 17762
rect 4780 17710 4832 17762
rect 4848 17710 4895 17762
rect 4895 17710 4900 17762
rect 4712 17646 4717 17698
rect 4717 17646 4764 17698
rect 4780 17646 4832 17698
rect 4848 17646 4895 17698
rect 4895 17646 4900 17698
rect 4712 17582 4717 17634
rect 4717 17582 4764 17634
rect 4780 17582 4832 17634
rect 4848 17582 4895 17634
rect 4895 17582 4900 17634
rect 4712 17518 4717 17570
rect 4717 17518 4764 17570
rect 4780 17518 4832 17570
rect 4848 17518 4895 17570
rect 4895 17518 4900 17570
rect 4712 17454 4717 17506
rect 4717 17454 4764 17506
rect 4780 17454 4832 17506
rect 4848 17454 4895 17506
rect 4895 17454 4900 17506
rect 4712 17390 4717 17442
rect 4717 17390 4764 17442
rect 4780 17390 4832 17442
rect 4848 17390 4895 17442
rect 4895 17390 4900 17442
rect 4712 17326 4717 17378
rect 4717 17326 4764 17378
rect 4780 17326 4832 17378
rect 4848 17326 4895 17378
rect 4895 17326 4900 17378
rect 4712 17262 4717 17314
rect 4717 17262 4764 17314
rect 4780 17262 4832 17314
rect 4848 17262 4895 17314
rect 4895 17262 4900 17314
rect 4712 17198 4717 17250
rect 4717 17198 4764 17250
rect 4780 17198 4832 17250
rect 4848 17198 4895 17250
rect 4895 17198 4900 17250
rect 4712 17134 4717 17186
rect 4717 17134 4764 17186
rect 4780 17134 4832 17186
rect 4848 17134 4895 17186
rect 4895 17134 4900 17186
rect 4712 17070 4717 17122
rect 4717 17070 4764 17122
rect 4780 17070 4832 17122
rect 4848 17070 4895 17122
rect 4895 17070 4900 17122
rect 4712 17006 4717 17058
rect 4717 17006 4764 17058
rect 4780 17006 4832 17058
rect 4848 17006 4895 17058
rect 4895 17006 4900 17058
rect 4712 16942 4717 16994
rect 4717 16942 4764 16994
rect 4780 16942 4832 16994
rect 4848 16942 4895 16994
rect 4895 16942 4900 16994
rect 4712 16877 4717 16929
rect 4717 16877 4764 16929
rect 4780 16877 4832 16929
rect 4848 16877 4895 16929
rect 4895 16877 4900 16929
rect 4712 16812 4717 16864
rect 4717 16812 4764 16864
rect 4780 16812 4832 16864
rect 4848 16812 4895 16864
rect 4895 16812 4900 16864
rect 4712 16747 4717 16799
rect 4717 16747 4764 16799
rect 4780 16747 4832 16799
rect 4848 16747 4895 16799
rect 4895 16747 4900 16799
rect 4712 16682 4717 16734
rect 4717 16682 4764 16734
rect 4780 16682 4832 16734
rect 4848 16682 4895 16734
rect 4895 16682 4900 16734
rect 4712 16617 4717 16669
rect 4717 16617 4764 16669
rect 4780 16617 4832 16669
rect 4848 16617 4895 16669
rect 4895 16617 4900 16669
rect 4712 16552 4717 16604
rect 4717 16552 4764 16604
rect 4780 16552 4832 16604
rect 4848 16552 4895 16604
rect 4895 16552 4900 16604
rect 4712 16487 4717 16539
rect 4717 16487 4764 16539
rect 4780 16487 4832 16539
rect 4848 16487 4895 16539
rect 4895 16487 4900 16539
rect 4712 16422 4717 16474
rect 4717 16422 4764 16474
rect 4780 16422 4832 16474
rect 4848 16422 4895 16474
rect 4895 16422 4900 16474
rect 4712 16357 4717 16409
rect 4717 16357 4764 16409
rect 4780 16357 4832 16409
rect 4848 16357 4895 16409
rect 4895 16357 4900 16409
rect 4712 16292 4717 16344
rect 4717 16292 4764 16344
rect 4780 16292 4832 16344
rect 4848 16292 4895 16344
rect 4895 16292 4900 16344
rect 4712 16227 4717 16279
rect 4717 16227 4764 16279
rect 4780 16227 4832 16279
rect 4848 16227 4895 16279
rect 4895 16227 4900 16279
rect 4712 16162 4717 16214
rect 4717 16162 4764 16214
rect 4780 16162 4832 16214
rect 4848 16162 4895 16214
rect 4895 16162 4900 16214
rect 2233 13544 2285 13550
rect 2335 13544 2387 13550
rect 2233 13498 2285 13544
rect 2335 13498 2387 13544
rect 2233 13434 2285 13486
rect 2335 13434 2387 13486
rect 2233 13370 2285 13422
rect 2335 13370 2387 13422
rect 2233 13306 2285 13358
rect 2335 13306 2387 13358
rect 2233 13242 2285 13294
rect 2335 13242 2387 13294
rect 2233 13178 2285 13230
rect 2335 13178 2387 13230
rect 2233 13114 2285 13166
rect 2335 13114 2387 13166
rect 2233 13050 2285 13102
rect 2335 13050 2387 13102
rect 2233 12986 2285 13038
rect 2335 12986 2387 13038
rect 2233 12922 2285 12974
rect 2335 12922 2387 12974
rect 2233 12858 2285 12910
rect 2335 12858 2387 12910
rect 2233 12794 2285 12846
rect 2335 12794 2387 12846
rect 2233 12730 2285 12782
rect 2335 12730 2387 12782
rect 2233 12666 2285 12718
rect 2335 12666 2387 12718
rect 2233 12602 2285 12654
rect 2335 12602 2387 12654
rect 2233 12538 2285 12590
rect 2335 12538 2387 12590
rect 2233 12474 2285 12526
rect 2335 12474 2387 12526
rect 2233 12410 2285 12462
rect 2335 12410 2387 12462
rect 2233 12346 2285 12398
rect 2335 12346 2387 12398
rect 2233 12282 2285 12334
rect 2335 12282 2387 12334
rect 2233 12218 2285 12270
rect 2335 12218 2387 12270
rect 2233 12154 2285 12206
rect 2335 12154 2387 12206
rect 2233 12090 2285 12142
rect 2335 12090 2387 12142
rect 2233 12026 2285 12078
rect 2335 12026 2387 12078
rect 2233 11962 2285 12014
rect 2335 11962 2387 12014
rect 2233 11898 2285 11950
rect 2335 11898 2387 11950
rect 2233 11834 2285 11886
rect 2335 11834 2387 11886
rect 2233 11770 2285 11822
rect 2335 11770 2387 11822
rect 2233 11705 2285 11757
rect 2335 11705 2387 11757
rect 2233 11640 2285 11692
rect 2335 11640 2387 11692
rect 2233 11575 2285 11627
rect 2335 11575 2387 11627
rect 2233 11510 2285 11562
rect 2335 11510 2387 11562
rect 2233 11445 2285 11497
rect 2335 11445 2387 11497
rect 2233 11380 2285 11432
rect 2335 11380 2387 11432
rect 2233 11315 2285 11367
rect 2335 11315 2387 11367
rect 2233 11250 2285 11302
rect 2335 11250 2387 11302
rect 2233 11185 2285 11237
rect 2335 11185 2387 11237
rect 2233 11120 2285 11172
rect 2335 11134 2387 11172
rect 2335 11120 2387 11134
rect 2233 11062 2285 11107
rect 2335 11095 2387 11107
rect 2233 11055 2285 11062
rect 2335 11061 2365 11095
rect 2365 11061 2387 11095
rect 2335 11055 2387 11061
rect 2233 11023 2285 11042
rect 2233 10990 2255 11023
rect 2255 10990 2285 11023
rect 2335 11022 2387 11042
rect 2335 10990 2365 11022
rect 2365 10990 2387 11022
rect 2233 10950 2285 10977
rect 2233 10925 2255 10950
rect 2255 10925 2285 10950
rect 2335 10949 2387 10977
rect 2335 10925 2365 10949
rect 2365 10925 2387 10949
rect 2233 10877 2285 10912
rect 2233 10860 2255 10877
rect 2255 10860 2285 10877
rect 2233 10843 2255 10847
rect 2255 10843 2285 10847
rect 2335 10876 2387 10912
rect 2335 10860 2365 10876
rect 2365 10860 2387 10876
rect 2233 10804 2285 10843
rect 2335 10842 2365 10847
rect 2365 10842 2387 10847
rect 2233 10795 2255 10804
rect 2255 10795 2285 10804
rect 2233 10770 2255 10782
rect 2255 10770 2285 10782
rect 2335 10803 2387 10842
rect 2335 10795 2365 10803
rect 2365 10795 2387 10803
rect 2233 10731 2285 10770
rect 2335 10769 2365 10782
rect 2365 10769 2387 10782
rect 2233 10730 2255 10731
rect 2255 10730 2285 10731
rect 2233 10697 2255 10717
rect 2255 10697 2285 10717
rect 2335 10730 2387 10769
rect 2233 10665 2285 10697
rect 2335 10696 2365 10717
rect 2365 10696 2387 10717
rect 2335 10665 2387 10696
rect 2233 10624 2255 10652
rect 2255 10624 2285 10652
rect 2233 10600 2285 10624
rect 2335 10623 2365 10652
rect 2365 10623 2387 10652
rect 2335 10600 2387 10623
rect 2233 10585 2285 10587
rect 2233 10551 2255 10585
rect 2255 10551 2285 10585
rect 2335 10584 2387 10587
rect 2233 10535 2285 10551
rect 2335 10550 2365 10584
rect 2365 10550 2387 10584
rect 2335 10535 2387 10550
rect 2233 10512 2285 10522
rect 2233 10478 2255 10512
rect 2255 10478 2285 10512
rect 2335 10511 2387 10522
rect 2233 10470 2285 10478
rect 2335 10477 2365 10511
rect 2365 10477 2387 10511
rect 2335 10470 2387 10477
rect 2233 10439 2285 10457
rect 2233 10405 2255 10439
rect 2255 10405 2285 10439
rect 2335 10438 2387 10457
rect 2335 10405 2365 10438
rect 2365 10405 2387 10438
rect 2233 10366 2285 10392
rect 2233 10340 2255 10366
rect 2255 10340 2285 10366
rect 2335 10365 2387 10392
rect 2335 10340 2365 10365
rect 2365 10340 2387 10365
rect 2233 10293 2285 10327
rect 2233 10275 2255 10293
rect 2255 10275 2285 10293
rect 2233 10259 2255 10262
rect 2255 10259 2285 10262
rect 2335 10292 2387 10327
rect 2335 10275 2365 10292
rect 2365 10275 2387 10292
rect 2233 10220 2285 10259
rect 2335 10258 2365 10262
rect 2365 10258 2387 10262
rect 2233 10210 2255 10220
rect 2255 10210 2285 10220
rect 2233 10186 2255 10197
rect 2255 10186 2285 10197
rect 2335 10219 2387 10258
rect 2335 10210 2365 10219
rect 2365 10210 2387 10219
rect 2233 10147 2285 10186
rect 2335 10185 2365 10197
rect 2365 10185 2387 10197
rect 2233 10145 2255 10147
rect 2255 10145 2285 10147
rect 2233 10113 2255 10132
rect 2255 10113 2285 10132
rect 2335 10146 2387 10185
rect 2335 10145 2365 10146
rect 2365 10145 2387 10146
rect 2233 10080 2285 10113
rect 2335 10112 2365 10132
rect 2365 10112 2387 10132
rect 2335 10080 2387 10112
rect 2233 10040 2255 10067
rect 2255 10040 2285 10067
rect 2233 10015 2285 10040
rect 2335 10039 2365 10067
rect 2365 10039 2387 10067
rect 2335 10015 2387 10039
rect 2233 10001 2285 10002
rect 2233 9967 2255 10001
rect 2255 9967 2285 10001
rect 2335 10000 2387 10002
rect 2233 9950 2285 9967
rect 2335 9966 2365 10000
rect 2365 9966 2387 10000
rect 2335 9950 2387 9966
rect 2233 9928 2285 9937
rect 2233 9894 2255 9928
rect 2255 9894 2285 9928
rect 2335 9927 2387 9937
rect 2233 9885 2285 9894
rect 2335 9893 2365 9927
rect 2365 9893 2387 9927
rect 2335 9885 2387 9893
rect 2233 9855 2285 9872
rect 2233 9821 2255 9855
rect 2255 9821 2285 9855
rect 2335 9854 2387 9872
rect 2233 9820 2285 9821
rect 2335 9820 2365 9854
rect 2365 9820 2387 9854
rect 2233 9782 2285 9807
rect 2233 9755 2255 9782
rect 2255 9755 2285 9782
rect 2335 9781 2387 9807
rect 2335 9755 2365 9781
rect 2365 9755 2387 9781
rect 2233 9709 2285 9742
rect 2233 9690 2255 9709
rect 2255 9690 2285 9709
rect 2233 9675 2255 9677
rect 2255 9675 2285 9677
rect 2335 9708 2387 9742
rect 2335 9690 2365 9708
rect 2365 9690 2387 9708
rect 2233 9636 2285 9675
rect 2335 9674 2365 9677
rect 2365 9674 2387 9677
rect 2233 9625 2255 9636
rect 2255 9625 2285 9636
rect 2233 9602 2255 9612
rect 2255 9602 2285 9612
rect 2335 9635 2387 9674
rect 2335 9625 2365 9635
rect 2365 9625 2387 9635
rect 2233 9563 2285 9602
rect 2335 9601 2365 9612
rect 2365 9601 2387 9612
rect 2233 9560 2255 9563
rect 2255 9560 2285 9563
rect 2233 9529 2255 9547
rect 2255 9529 2285 9547
rect 2335 9562 2387 9601
rect 2335 9560 2365 9562
rect 2365 9560 2387 9562
rect 2233 9495 2285 9529
rect 2335 9528 2365 9547
rect 2365 9528 2387 9547
rect 2335 9495 2387 9528
rect 2233 9456 2255 9482
rect 2255 9456 2285 9482
rect 2233 9430 2285 9456
rect 2335 9455 2365 9482
rect 2365 9455 2387 9482
rect 2335 9430 2387 9455
rect 2233 9383 2255 9417
rect 2255 9383 2285 9417
rect 2335 9416 2387 9417
rect 2233 9365 2285 9383
rect 2335 9382 2365 9416
rect 2365 9382 2387 9416
rect 2335 9365 2387 9382
rect 2872 13371 2924 13377
rect 2940 13371 2992 13377
rect 3008 13371 3060 13377
rect 2872 13325 2877 13371
rect 2877 13325 2924 13371
rect 2940 13325 2992 13371
rect 3008 13325 3055 13371
rect 3055 13325 3060 13371
rect 2872 13260 2877 13312
rect 2877 13260 2924 13312
rect 2940 13260 2992 13312
rect 3008 13260 3055 13312
rect 3055 13260 3060 13312
rect 2872 13195 2877 13247
rect 2877 13195 2924 13247
rect 2940 13195 2992 13247
rect 3008 13195 3055 13247
rect 3055 13195 3060 13247
rect 2872 13130 2877 13182
rect 2877 13130 2924 13182
rect 2940 13130 2992 13182
rect 3008 13130 3055 13182
rect 3055 13130 3060 13182
rect 2872 13065 2877 13117
rect 2877 13065 2924 13117
rect 2940 13065 2992 13117
rect 3008 13065 3055 13117
rect 3055 13065 3060 13117
rect 2872 13000 2877 13052
rect 2877 13000 2924 13052
rect 2940 13000 2992 13052
rect 3008 13000 3055 13052
rect 3055 13000 3060 13052
rect 2872 12935 2877 12987
rect 2877 12935 2924 12987
rect 2940 12935 2992 12987
rect 3008 12935 3055 12987
rect 3055 12935 3060 12987
rect 2872 12870 2877 12922
rect 2877 12870 2924 12922
rect 2940 12870 2992 12922
rect 3008 12870 3055 12922
rect 3055 12870 3060 12922
rect 2872 12805 2877 12857
rect 2877 12805 2924 12857
rect 2940 12805 2992 12857
rect 3008 12805 3055 12857
rect 3055 12805 3060 12857
rect 2872 12740 2877 12792
rect 2877 12740 2924 12792
rect 2940 12740 2992 12792
rect 3008 12740 3055 12792
rect 3055 12740 3060 12792
rect 2872 12675 2877 12727
rect 2877 12675 2924 12727
rect 2940 12675 2992 12727
rect 3008 12675 3055 12727
rect 3055 12675 3060 12727
rect 2872 12610 2877 12662
rect 2877 12610 2924 12662
rect 2940 12610 2992 12662
rect 3008 12610 3055 12662
rect 3055 12610 3060 12662
rect 2872 12545 2877 12597
rect 2877 12545 2924 12597
rect 2940 12545 2992 12597
rect 3008 12545 3055 12597
rect 3055 12545 3060 12597
rect 2872 12480 2877 12532
rect 2877 12480 2924 12532
rect 2940 12480 2992 12532
rect 3008 12480 3055 12532
rect 3055 12480 3060 12532
rect 2872 12415 2877 12467
rect 2877 12415 2924 12467
rect 2940 12415 2992 12467
rect 3008 12415 3055 12467
rect 3055 12415 3060 12467
rect 2872 12350 2877 12402
rect 2877 12350 2924 12402
rect 2940 12350 2992 12402
rect 3008 12350 3055 12402
rect 3055 12350 3060 12402
rect 2872 12285 2877 12337
rect 2877 12285 2924 12337
rect 2940 12285 2992 12337
rect 3008 12285 3055 12337
rect 3055 12285 3060 12337
rect 2872 12220 2877 12272
rect 2877 12220 2924 12272
rect 2940 12220 2992 12272
rect 3008 12220 3055 12272
rect 3055 12220 3060 12272
rect 2872 12155 2877 12207
rect 2877 12155 2924 12207
rect 2940 12155 2992 12207
rect 3008 12155 3055 12207
rect 3055 12155 3060 12207
rect 2872 12090 2877 12142
rect 2877 12090 2924 12142
rect 2940 12090 2992 12142
rect 3008 12090 3055 12142
rect 3055 12090 3060 12142
rect 2872 12024 2877 12076
rect 2877 12024 2924 12076
rect 2940 12024 2992 12076
rect 3008 12024 3055 12076
rect 3055 12024 3060 12076
rect 2872 11958 2877 12010
rect 2877 11958 2924 12010
rect 2940 11958 2992 12010
rect 3008 11958 3055 12010
rect 3055 11958 3060 12010
rect 2872 11892 2877 11944
rect 2877 11892 2924 11944
rect 2940 11892 2992 11944
rect 3008 11892 3055 11944
rect 3055 11892 3060 11944
rect 2872 11826 2877 11878
rect 2877 11826 2924 11878
rect 2940 11826 2992 11878
rect 3008 11826 3055 11878
rect 3055 11826 3060 11878
rect 2872 11760 2877 11812
rect 2877 11760 2924 11812
rect 2940 11760 2992 11812
rect 3008 11760 3055 11812
rect 3055 11760 3060 11812
rect 2872 11694 2877 11746
rect 2877 11694 2924 11746
rect 2940 11694 2992 11746
rect 3008 11694 3055 11746
rect 3055 11694 3060 11746
rect 2872 11628 2877 11680
rect 2877 11628 2924 11680
rect 2940 11628 2992 11680
rect 3008 11628 3055 11680
rect 3055 11628 3060 11680
rect 2872 11562 2877 11614
rect 2877 11562 2924 11614
rect 2940 11562 2992 11614
rect 3008 11562 3055 11614
rect 3055 11562 3060 11614
rect 3792 13238 3797 13290
rect 3797 13238 3844 13290
rect 3860 13238 3912 13290
rect 3928 13238 3975 13290
rect 3975 13238 3980 13290
rect 3792 13174 3797 13226
rect 3797 13174 3844 13226
rect 3860 13174 3912 13226
rect 3928 13174 3975 13226
rect 3975 13174 3980 13226
rect 3792 13110 3797 13162
rect 3797 13110 3844 13162
rect 3860 13110 3912 13162
rect 3928 13110 3975 13162
rect 3975 13110 3980 13162
rect 3792 13046 3797 13098
rect 3797 13046 3844 13098
rect 3860 13046 3912 13098
rect 3928 13046 3975 13098
rect 3975 13046 3980 13098
rect 3792 12982 3797 13034
rect 3797 12982 3844 13034
rect 3860 12982 3912 13034
rect 3928 12982 3975 13034
rect 3975 12982 3980 13034
rect 3792 12918 3797 12970
rect 3797 12918 3844 12970
rect 3860 12918 3912 12970
rect 3928 12918 3975 12970
rect 3975 12918 3980 12970
rect 3792 12854 3797 12906
rect 3797 12854 3844 12906
rect 3860 12854 3912 12906
rect 3928 12854 3975 12906
rect 3975 12854 3980 12906
rect 3792 12790 3797 12842
rect 3797 12790 3844 12842
rect 3860 12790 3912 12842
rect 3928 12790 3975 12842
rect 3975 12790 3980 12842
rect 3792 12726 3797 12778
rect 3797 12726 3844 12778
rect 3860 12726 3912 12778
rect 3928 12726 3975 12778
rect 3975 12726 3980 12778
rect 3792 12662 3797 12714
rect 3797 12662 3844 12714
rect 3860 12662 3912 12714
rect 3928 12662 3975 12714
rect 3975 12662 3980 12714
rect 3792 12598 3797 12650
rect 3797 12598 3844 12650
rect 3860 12598 3912 12650
rect 3928 12598 3975 12650
rect 3975 12598 3980 12650
rect 3792 12534 3797 12586
rect 3797 12534 3844 12586
rect 3860 12534 3912 12586
rect 3928 12534 3975 12586
rect 3975 12534 3980 12586
rect 3792 12470 3797 12522
rect 3797 12470 3844 12522
rect 3860 12470 3912 12522
rect 3928 12470 3975 12522
rect 3975 12470 3980 12522
rect 3792 12406 3797 12458
rect 3797 12406 3844 12458
rect 3860 12406 3912 12458
rect 3928 12406 3975 12458
rect 3975 12406 3980 12458
rect 3792 12342 3797 12394
rect 3797 12342 3844 12394
rect 3860 12342 3912 12394
rect 3928 12342 3975 12394
rect 3975 12342 3980 12394
rect 3792 12277 3797 12329
rect 3797 12277 3844 12329
rect 3860 12277 3912 12329
rect 3928 12277 3975 12329
rect 3975 12277 3980 12329
rect 3792 12212 3797 12264
rect 3797 12212 3844 12264
rect 3860 12212 3912 12264
rect 3928 12212 3975 12264
rect 3975 12212 3980 12264
rect 3792 12147 3797 12199
rect 3797 12147 3844 12199
rect 3860 12147 3912 12199
rect 3928 12147 3975 12199
rect 3975 12147 3980 12199
rect 3792 12082 3797 12134
rect 3797 12082 3844 12134
rect 3860 12082 3912 12134
rect 3928 12082 3975 12134
rect 3975 12082 3980 12134
rect 3792 12017 3797 12069
rect 3797 12017 3844 12069
rect 3860 12017 3912 12069
rect 3928 12017 3975 12069
rect 3975 12017 3980 12069
rect 3792 11952 3797 12004
rect 3797 11952 3844 12004
rect 3860 11952 3912 12004
rect 3928 11952 3975 12004
rect 3975 11952 3980 12004
rect 3792 11887 3797 11939
rect 3797 11887 3844 11939
rect 3860 11887 3912 11939
rect 3928 11887 3975 11939
rect 3975 11887 3980 11939
rect 3792 11822 3797 11874
rect 3797 11822 3844 11874
rect 3860 11822 3912 11874
rect 3928 11822 3975 11874
rect 3975 11822 3980 11874
rect 3792 11757 3797 11809
rect 3797 11757 3844 11809
rect 3860 11757 3912 11809
rect 3928 11757 3975 11809
rect 3975 11757 3980 11809
rect 3792 11692 3797 11744
rect 3797 11692 3844 11744
rect 3860 11692 3912 11744
rect 3928 11692 3975 11744
rect 3975 11692 3980 11744
rect 3792 11627 3797 11679
rect 3797 11627 3844 11679
rect 3860 11627 3912 11679
rect 3928 11627 3975 11679
rect 3975 11627 3980 11679
rect 3792 11562 3797 11614
rect 3797 11562 3844 11614
rect 3860 11562 3912 11614
rect 3928 11562 3975 11614
rect 3975 11562 3980 11614
rect 3361 10895 3413 10947
rect 3439 10895 3491 10947
rect 3361 10829 3413 10881
rect 3439 10829 3491 10881
rect 3361 10763 3413 10815
rect 3439 10763 3491 10815
rect 3361 10697 3413 10749
rect 3439 10697 3491 10749
rect 3361 10631 3413 10683
rect 3439 10631 3491 10683
rect 3361 10565 3413 10617
rect 3439 10565 3491 10617
rect 3361 10499 3413 10551
rect 3439 10499 3491 10551
rect 3361 10433 3413 10485
rect 3439 10433 3491 10485
rect 3361 10367 3413 10419
rect 3439 10367 3491 10419
rect 3361 10301 3413 10353
rect 3439 10301 3491 10353
rect 3361 10234 3413 10286
rect 3439 10234 3491 10286
rect 3361 10167 3413 10219
rect 3439 10167 3491 10219
rect 3361 10100 3413 10152
rect 3439 10100 3491 10152
rect 3361 10033 3413 10085
rect 3439 10033 3491 10085
rect 3361 9966 3413 10018
rect 3439 9966 3491 10018
rect 3361 9899 3413 9951
rect 3439 9899 3491 9951
rect 3361 9832 3413 9884
rect 3439 9832 3491 9884
rect 3361 9765 3413 9817
rect 3439 9765 3491 9817
rect 3361 9698 3413 9750
rect 3439 9698 3491 9750
rect 3361 9631 3413 9683
rect 3439 9631 3491 9683
rect 3361 9564 3413 9616
rect 3439 9564 3491 9616
rect 3361 9497 3413 9549
rect 3439 9497 3491 9549
rect 4712 13238 4717 13290
rect 4717 13238 4764 13290
rect 4780 13238 4832 13290
rect 4848 13238 4895 13290
rect 4895 13238 4900 13290
rect 4712 13174 4717 13226
rect 4717 13174 4764 13226
rect 4780 13174 4832 13226
rect 4848 13174 4895 13226
rect 4895 13174 4900 13226
rect 4712 13110 4717 13162
rect 4717 13110 4764 13162
rect 4780 13110 4832 13162
rect 4848 13110 4895 13162
rect 4895 13110 4900 13162
rect 4712 13046 4717 13098
rect 4717 13046 4764 13098
rect 4780 13046 4832 13098
rect 4848 13046 4895 13098
rect 4895 13046 4900 13098
rect 4712 12982 4717 13034
rect 4717 12982 4764 13034
rect 4780 12982 4832 13034
rect 4848 12982 4895 13034
rect 4895 12982 4900 13034
rect 4712 12918 4717 12970
rect 4717 12918 4764 12970
rect 4780 12918 4832 12970
rect 4848 12918 4895 12970
rect 4895 12918 4900 12970
rect 4712 12854 4717 12906
rect 4717 12854 4764 12906
rect 4780 12854 4832 12906
rect 4848 12854 4895 12906
rect 4895 12854 4900 12906
rect 4712 12790 4717 12842
rect 4717 12790 4764 12842
rect 4780 12790 4832 12842
rect 4848 12790 4895 12842
rect 4895 12790 4900 12842
rect 4712 12726 4717 12778
rect 4717 12726 4764 12778
rect 4780 12726 4832 12778
rect 4848 12726 4895 12778
rect 4895 12726 4900 12778
rect 4712 12662 4717 12714
rect 4717 12662 4764 12714
rect 4780 12662 4832 12714
rect 4848 12662 4895 12714
rect 4895 12662 4900 12714
rect 4712 12598 4717 12650
rect 4717 12598 4764 12650
rect 4780 12598 4832 12650
rect 4848 12598 4895 12650
rect 4895 12598 4900 12650
rect 4712 12534 4717 12586
rect 4717 12534 4764 12586
rect 4780 12534 4832 12586
rect 4848 12534 4895 12586
rect 4895 12534 4900 12586
rect 4712 12470 4717 12522
rect 4717 12470 4764 12522
rect 4780 12470 4832 12522
rect 4848 12470 4895 12522
rect 4895 12470 4900 12522
rect 4712 12406 4717 12458
rect 4717 12406 4764 12458
rect 4780 12406 4832 12458
rect 4848 12406 4895 12458
rect 4895 12406 4900 12458
rect 4712 12342 4717 12394
rect 4717 12342 4764 12394
rect 4780 12342 4832 12394
rect 4848 12342 4895 12394
rect 4895 12342 4900 12394
rect 4712 12277 4717 12329
rect 4717 12277 4764 12329
rect 4780 12277 4832 12329
rect 4848 12277 4895 12329
rect 4895 12277 4900 12329
rect 4712 12212 4717 12264
rect 4717 12212 4764 12264
rect 4780 12212 4832 12264
rect 4848 12212 4895 12264
rect 4895 12212 4900 12264
rect 4712 12147 4717 12199
rect 4717 12147 4764 12199
rect 4780 12147 4832 12199
rect 4848 12147 4895 12199
rect 4895 12147 4900 12199
rect 4712 12082 4717 12134
rect 4717 12082 4764 12134
rect 4780 12082 4832 12134
rect 4848 12082 4895 12134
rect 4895 12082 4900 12134
rect 4712 12017 4717 12069
rect 4717 12017 4764 12069
rect 4780 12017 4832 12069
rect 4848 12017 4895 12069
rect 4895 12017 4900 12069
rect 4712 11952 4717 12004
rect 4717 11952 4764 12004
rect 4780 11952 4832 12004
rect 4848 11952 4895 12004
rect 4895 11952 4900 12004
rect 4712 11887 4717 11939
rect 4717 11887 4764 11939
rect 4780 11887 4832 11939
rect 4848 11887 4895 11939
rect 4895 11887 4900 11939
rect 4712 11822 4717 11874
rect 4717 11822 4764 11874
rect 4780 11822 4832 11874
rect 4848 11822 4895 11874
rect 4895 11822 4900 11874
rect 4712 11757 4717 11809
rect 4717 11757 4764 11809
rect 4780 11757 4832 11809
rect 4848 11757 4895 11809
rect 4895 11757 4900 11809
rect 4712 11692 4717 11744
rect 4717 11692 4764 11744
rect 4780 11692 4832 11744
rect 4848 11692 4895 11744
rect 4895 11692 4900 11744
rect 4712 11627 4717 11679
rect 4717 11627 4764 11679
rect 4780 11627 4832 11679
rect 4848 11627 4895 11679
rect 4895 11627 4900 11679
rect 4712 11562 4717 11614
rect 4717 11562 4764 11614
rect 4780 11562 4832 11614
rect 4848 11562 4895 11614
rect 4895 11562 4900 11614
rect 4281 11173 4333 11225
rect 4359 11173 4411 11225
rect 4281 11109 4333 11161
rect 4359 11109 4411 11161
rect 4281 11045 4333 11097
rect 4359 11045 4411 11097
rect 4281 10981 4333 11033
rect 4359 10981 4411 11033
rect 4281 10917 4333 10969
rect 4359 10917 4411 10969
rect 4281 10853 4333 10905
rect 4359 10853 4411 10905
rect 4281 10789 4333 10841
rect 4359 10789 4411 10841
rect 4281 10725 4333 10777
rect 4359 10725 4411 10777
rect 4281 10661 4333 10713
rect 4359 10661 4411 10713
rect 4281 10597 4333 10649
rect 4359 10597 4411 10649
rect 4281 10533 4333 10585
rect 4359 10533 4411 10585
rect 4281 10469 4333 10521
rect 4359 10469 4411 10521
rect 4281 10405 4333 10457
rect 4359 10405 4411 10457
rect 4281 10341 4333 10393
rect 4359 10341 4411 10393
rect 4281 10277 4333 10329
rect 4359 10277 4411 10329
rect 4281 10212 4333 10264
rect 4359 10212 4411 10264
rect 4281 10147 4333 10199
rect 4359 10147 4411 10199
rect 4281 10082 4333 10134
rect 4359 10082 4411 10134
rect 4281 10017 4333 10069
rect 4359 10017 4411 10069
rect 4281 9952 4333 10004
rect 4359 9952 4411 10004
rect 4281 9887 4333 9939
rect 4359 9887 4411 9939
rect 4281 9822 4333 9874
rect 4359 9822 4411 9874
rect 4281 9757 4333 9809
rect 4359 9757 4411 9809
rect 4281 9692 4333 9744
rect 4359 9692 4411 9744
rect 4281 9627 4333 9679
rect 4359 9627 4411 9679
rect 4281 9562 4333 9614
rect 4359 9562 4411 9614
rect 4281 9497 4333 9549
rect 4359 9497 4411 9549
rect 5201 20373 5253 20425
rect 5279 20373 5331 20425
rect 5201 20309 5253 20361
rect 5279 20309 5331 20361
rect 5201 20245 5253 20297
rect 5279 20245 5331 20297
rect 5201 20181 5253 20233
rect 5279 20181 5331 20233
rect 5201 20117 5253 20169
rect 5279 20117 5331 20169
rect 5201 20053 5253 20105
rect 5279 20053 5331 20105
rect 5201 19989 5253 20041
rect 5279 19989 5331 20041
rect 5201 19925 5253 19977
rect 5279 19925 5331 19977
rect 5201 19861 5253 19913
rect 5279 19861 5331 19913
rect 5201 19797 5253 19849
rect 5279 19797 5331 19849
rect 5201 19733 5253 19785
rect 5279 19733 5331 19785
rect 5201 19669 5253 19721
rect 5279 19669 5331 19721
rect 5201 19605 5253 19657
rect 5279 19605 5331 19657
rect 5201 19541 5253 19593
rect 5279 19541 5331 19593
rect 5201 19477 5253 19529
rect 5279 19477 5331 19529
rect 5201 19412 5253 19464
rect 5279 19412 5331 19464
rect 5201 19347 5253 19399
rect 5279 19347 5331 19399
rect 5201 19282 5253 19334
rect 5279 19282 5331 19334
rect 5201 19217 5253 19269
rect 5279 19217 5331 19269
rect 5201 19152 5253 19204
rect 5279 19152 5331 19204
rect 5201 19087 5253 19139
rect 5279 19087 5331 19139
rect 5201 19022 5253 19074
rect 5279 19022 5331 19074
rect 5201 18957 5253 19009
rect 5279 18957 5331 19009
rect 5201 18892 5253 18944
rect 5279 18892 5331 18944
rect 5201 18827 5253 18879
rect 5279 18827 5331 18879
rect 5201 18762 5253 18814
rect 5279 18762 5331 18814
rect 5201 18697 5253 18749
rect 5279 18697 5331 18749
rect 5201 15773 5253 15825
rect 5279 15773 5331 15825
rect 5201 15709 5253 15761
rect 5279 15709 5331 15761
rect 5201 15645 5253 15697
rect 5279 15645 5331 15697
rect 5201 15581 5253 15633
rect 5279 15581 5331 15633
rect 5201 15517 5253 15569
rect 5279 15517 5331 15569
rect 5201 15453 5253 15505
rect 5279 15453 5331 15505
rect 5201 15389 5253 15441
rect 5279 15389 5331 15441
rect 5201 15325 5253 15377
rect 5279 15325 5331 15377
rect 5201 15261 5253 15313
rect 5279 15261 5331 15313
rect 5201 15197 5253 15249
rect 5279 15197 5331 15249
rect 5201 15133 5253 15185
rect 5279 15133 5331 15185
rect 5201 15069 5253 15121
rect 5279 15069 5331 15121
rect 5201 15005 5253 15057
rect 5279 15005 5331 15057
rect 5201 14941 5253 14993
rect 5279 14941 5331 14993
rect 5201 14877 5253 14929
rect 5279 14877 5331 14929
rect 5201 14812 5253 14864
rect 5279 14812 5331 14864
rect 5201 14747 5253 14799
rect 5279 14747 5331 14799
rect 5201 14682 5253 14734
rect 5279 14682 5331 14734
rect 5201 14617 5253 14669
rect 5279 14617 5331 14669
rect 5201 14552 5253 14604
rect 5279 14552 5331 14604
rect 5201 14487 5253 14539
rect 5279 14487 5331 14539
rect 5201 14422 5253 14474
rect 5279 14422 5331 14474
rect 5201 14357 5253 14409
rect 5279 14357 5331 14409
rect 5201 14292 5253 14344
rect 5279 14292 5331 14344
rect 5201 14227 5253 14279
rect 5279 14227 5331 14279
rect 5201 14162 5253 14214
rect 5279 14162 5331 14214
rect 5201 14097 5253 14149
rect 5279 14097 5331 14149
rect 5201 11173 5253 11225
rect 5279 11173 5331 11225
rect 5201 11109 5253 11161
rect 5279 11109 5331 11161
rect 5201 11045 5253 11097
rect 5279 11045 5331 11097
rect 5201 10981 5253 11033
rect 5279 10981 5331 11033
rect 5201 10917 5253 10969
rect 5279 10917 5331 10969
rect 5201 10853 5253 10905
rect 5279 10853 5331 10905
rect 5201 10789 5253 10841
rect 5279 10789 5331 10841
rect 5201 10725 5253 10777
rect 5279 10725 5331 10777
rect 5201 10661 5253 10713
rect 5279 10661 5331 10713
rect 5201 10597 5253 10649
rect 5279 10597 5331 10649
rect 5201 10533 5253 10585
rect 5279 10533 5331 10585
rect 5201 10469 5253 10521
rect 5279 10469 5331 10521
rect 5201 10405 5253 10457
rect 5279 10405 5331 10457
rect 5201 10341 5253 10393
rect 5279 10341 5331 10393
rect 5201 10277 5253 10329
rect 5279 10277 5331 10329
rect 5201 10212 5253 10264
rect 5279 10212 5331 10264
rect 5201 10147 5253 10199
rect 5279 10147 5331 10199
rect 5201 10082 5253 10134
rect 5279 10082 5331 10134
rect 5201 10017 5253 10069
rect 5279 10017 5331 10069
rect 5201 9952 5253 10004
rect 5279 9952 5331 10004
rect 5201 9887 5253 9939
rect 5279 9887 5331 9939
rect 5201 9822 5253 9874
rect 5279 9822 5331 9874
rect 5201 9757 5253 9809
rect 5279 9757 5331 9809
rect 5201 9692 5253 9744
rect 5279 9692 5331 9744
rect 5201 9627 5253 9679
rect 5279 9627 5331 9679
rect 5201 9562 5253 9614
rect 5279 9562 5331 9614
rect 5201 9497 5253 9549
rect 5279 9497 5331 9549
rect 5632 36238 5637 36290
rect 5637 36238 5684 36290
rect 5700 36238 5752 36290
rect 5768 36238 5815 36290
rect 5815 36238 5820 36290
rect 5632 36174 5637 36226
rect 5637 36174 5684 36226
rect 5700 36174 5752 36226
rect 5768 36174 5815 36226
rect 5815 36174 5820 36226
rect 5632 36110 5637 36162
rect 5637 36110 5684 36162
rect 5700 36110 5752 36162
rect 5768 36110 5815 36162
rect 5815 36110 5820 36162
rect 5632 36046 5637 36098
rect 5637 36046 5684 36098
rect 5700 36046 5752 36098
rect 5768 36046 5815 36098
rect 5815 36046 5820 36098
rect 5632 35982 5637 36034
rect 5637 35982 5684 36034
rect 5700 35982 5752 36034
rect 5768 35982 5815 36034
rect 5815 35982 5820 36034
rect 5632 35918 5637 35970
rect 5637 35918 5684 35970
rect 5700 35918 5752 35970
rect 5768 35918 5815 35970
rect 5815 35918 5820 35970
rect 5632 35854 5637 35906
rect 5637 35854 5684 35906
rect 5700 35854 5752 35906
rect 5768 35854 5815 35906
rect 5815 35854 5820 35906
rect 5632 35790 5637 35842
rect 5637 35790 5684 35842
rect 5700 35790 5752 35842
rect 5768 35790 5815 35842
rect 5815 35790 5820 35842
rect 5632 35726 5637 35778
rect 5637 35726 5684 35778
rect 5700 35726 5752 35778
rect 5768 35726 5815 35778
rect 5815 35726 5820 35778
rect 5632 35662 5637 35714
rect 5637 35662 5684 35714
rect 5700 35662 5752 35714
rect 5768 35662 5815 35714
rect 5815 35662 5820 35714
rect 5632 35598 5637 35650
rect 5637 35598 5684 35650
rect 5700 35598 5752 35650
rect 5768 35598 5815 35650
rect 5815 35598 5820 35650
rect 5632 35534 5637 35586
rect 5637 35534 5684 35586
rect 5700 35534 5752 35586
rect 5768 35534 5815 35586
rect 5815 35534 5820 35586
rect 5632 35470 5637 35522
rect 5637 35470 5684 35522
rect 5700 35470 5752 35522
rect 5768 35470 5815 35522
rect 5815 35470 5820 35522
rect 5632 35406 5637 35458
rect 5637 35406 5684 35458
rect 5700 35406 5752 35458
rect 5768 35406 5815 35458
rect 5815 35406 5820 35458
rect 5632 35342 5637 35394
rect 5637 35342 5684 35394
rect 5700 35342 5752 35394
rect 5768 35342 5815 35394
rect 5815 35342 5820 35394
rect 5632 35277 5637 35329
rect 5637 35277 5684 35329
rect 5700 35277 5752 35329
rect 5768 35277 5815 35329
rect 5815 35277 5820 35329
rect 5632 35212 5637 35264
rect 5637 35212 5684 35264
rect 5700 35212 5752 35264
rect 5768 35212 5815 35264
rect 5815 35212 5820 35264
rect 5632 35147 5637 35199
rect 5637 35147 5684 35199
rect 5700 35147 5752 35199
rect 5768 35147 5815 35199
rect 5815 35147 5820 35199
rect 5632 35082 5637 35134
rect 5637 35082 5684 35134
rect 5700 35082 5752 35134
rect 5768 35082 5815 35134
rect 5815 35082 5820 35134
rect 5632 35017 5637 35069
rect 5637 35017 5684 35069
rect 5700 35017 5752 35069
rect 5768 35017 5815 35069
rect 5815 35017 5820 35069
rect 5632 34952 5637 35004
rect 5637 34952 5684 35004
rect 5700 34952 5752 35004
rect 5768 34952 5815 35004
rect 5815 34952 5820 35004
rect 5632 34887 5637 34939
rect 5637 34887 5684 34939
rect 5700 34887 5752 34939
rect 5768 34887 5815 34939
rect 5815 34887 5820 34939
rect 5632 34822 5637 34874
rect 5637 34822 5684 34874
rect 5700 34822 5752 34874
rect 5768 34822 5815 34874
rect 5815 34822 5820 34874
rect 5632 34757 5637 34809
rect 5637 34757 5684 34809
rect 5700 34757 5752 34809
rect 5768 34757 5815 34809
rect 5815 34757 5820 34809
rect 5632 34692 5637 34744
rect 5637 34692 5684 34744
rect 5700 34692 5752 34744
rect 5768 34692 5815 34744
rect 5815 34692 5820 34744
rect 5632 34627 5637 34679
rect 5637 34627 5684 34679
rect 5700 34627 5752 34679
rect 5768 34627 5815 34679
rect 5815 34627 5820 34679
rect 5632 34562 5637 34614
rect 5637 34562 5684 34614
rect 5700 34562 5752 34614
rect 5768 34562 5815 34614
rect 5815 34562 5820 34614
rect 5632 31638 5637 31690
rect 5637 31638 5684 31690
rect 5700 31638 5752 31690
rect 5768 31638 5815 31690
rect 5815 31638 5820 31690
rect 5632 31574 5637 31626
rect 5637 31574 5684 31626
rect 5700 31574 5752 31626
rect 5768 31574 5815 31626
rect 5815 31574 5820 31626
rect 5632 31510 5637 31562
rect 5637 31510 5684 31562
rect 5700 31510 5752 31562
rect 5768 31510 5815 31562
rect 5815 31510 5820 31562
rect 5632 31446 5637 31498
rect 5637 31446 5684 31498
rect 5700 31446 5752 31498
rect 5768 31446 5815 31498
rect 5815 31446 5820 31498
rect 5632 31382 5637 31434
rect 5637 31382 5684 31434
rect 5700 31382 5752 31434
rect 5768 31382 5815 31434
rect 5815 31382 5820 31434
rect 5632 31318 5637 31370
rect 5637 31318 5684 31370
rect 5700 31318 5752 31370
rect 5768 31318 5815 31370
rect 5815 31318 5820 31370
rect 5632 31254 5637 31306
rect 5637 31254 5684 31306
rect 5700 31254 5752 31306
rect 5768 31254 5815 31306
rect 5815 31254 5820 31306
rect 5632 31190 5637 31242
rect 5637 31190 5684 31242
rect 5700 31190 5752 31242
rect 5768 31190 5815 31242
rect 5815 31190 5820 31242
rect 5632 31126 5637 31178
rect 5637 31126 5684 31178
rect 5700 31126 5752 31178
rect 5768 31126 5815 31178
rect 5815 31126 5820 31178
rect 5632 31062 5637 31114
rect 5637 31062 5684 31114
rect 5700 31062 5752 31114
rect 5768 31062 5815 31114
rect 5815 31062 5820 31114
rect 5632 30998 5637 31050
rect 5637 30998 5684 31050
rect 5700 30998 5752 31050
rect 5768 30998 5815 31050
rect 5815 30998 5820 31050
rect 5632 30934 5637 30986
rect 5637 30934 5684 30986
rect 5700 30934 5752 30986
rect 5768 30934 5815 30986
rect 5815 30934 5820 30986
rect 5632 30870 5637 30922
rect 5637 30870 5684 30922
rect 5700 30870 5752 30922
rect 5768 30870 5815 30922
rect 5815 30870 5820 30922
rect 5632 30806 5637 30858
rect 5637 30806 5684 30858
rect 5700 30806 5752 30858
rect 5768 30806 5815 30858
rect 5815 30806 5820 30858
rect 5632 30742 5637 30794
rect 5637 30742 5684 30794
rect 5700 30742 5752 30794
rect 5768 30742 5815 30794
rect 5815 30742 5820 30794
rect 5632 30677 5637 30729
rect 5637 30677 5684 30729
rect 5700 30677 5752 30729
rect 5768 30677 5815 30729
rect 5815 30677 5820 30729
rect 5632 30612 5637 30664
rect 5637 30612 5684 30664
rect 5700 30612 5752 30664
rect 5768 30612 5815 30664
rect 5815 30612 5820 30664
rect 5632 30547 5637 30599
rect 5637 30547 5684 30599
rect 5700 30547 5752 30599
rect 5768 30547 5815 30599
rect 5815 30547 5820 30599
rect 5632 30482 5637 30534
rect 5637 30482 5684 30534
rect 5700 30482 5752 30534
rect 5768 30482 5815 30534
rect 5815 30482 5820 30534
rect 5632 30417 5637 30469
rect 5637 30417 5684 30469
rect 5700 30417 5752 30469
rect 5768 30417 5815 30469
rect 5815 30417 5820 30469
rect 5632 30352 5637 30404
rect 5637 30352 5684 30404
rect 5700 30352 5752 30404
rect 5768 30352 5815 30404
rect 5815 30352 5820 30404
rect 5632 30287 5637 30339
rect 5637 30287 5684 30339
rect 5700 30287 5752 30339
rect 5768 30287 5815 30339
rect 5815 30287 5820 30339
rect 5632 30222 5637 30274
rect 5637 30222 5684 30274
rect 5700 30222 5752 30274
rect 5768 30222 5815 30274
rect 5815 30222 5820 30274
rect 5632 30157 5637 30209
rect 5637 30157 5684 30209
rect 5700 30157 5752 30209
rect 5768 30157 5815 30209
rect 5815 30157 5820 30209
rect 5632 30092 5637 30144
rect 5637 30092 5684 30144
rect 5700 30092 5752 30144
rect 5768 30092 5815 30144
rect 5815 30092 5820 30144
rect 5632 30027 5637 30079
rect 5637 30027 5684 30079
rect 5700 30027 5752 30079
rect 5768 30027 5815 30079
rect 5815 30027 5820 30079
rect 5632 29962 5637 30014
rect 5637 29962 5684 30014
rect 5700 29962 5752 30014
rect 5768 29962 5815 30014
rect 5815 29962 5820 30014
rect 5632 27038 5637 27090
rect 5637 27038 5684 27090
rect 5700 27038 5752 27090
rect 5768 27038 5815 27090
rect 5815 27038 5820 27090
rect 5632 26974 5637 27026
rect 5637 26974 5684 27026
rect 5700 26974 5752 27026
rect 5768 26974 5815 27026
rect 5815 26974 5820 27026
rect 5632 26910 5637 26962
rect 5637 26910 5684 26962
rect 5700 26910 5752 26962
rect 5768 26910 5815 26962
rect 5815 26910 5820 26962
rect 5632 26846 5637 26898
rect 5637 26846 5684 26898
rect 5700 26846 5752 26898
rect 5768 26846 5815 26898
rect 5815 26846 5820 26898
rect 5632 26782 5637 26834
rect 5637 26782 5684 26834
rect 5700 26782 5752 26834
rect 5768 26782 5815 26834
rect 5815 26782 5820 26834
rect 5632 26718 5637 26770
rect 5637 26718 5684 26770
rect 5700 26718 5752 26770
rect 5768 26718 5815 26770
rect 5815 26718 5820 26770
rect 5632 26654 5637 26706
rect 5637 26654 5684 26706
rect 5700 26654 5752 26706
rect 5768 26654 5815 26706
rect 5815 26654 5820 26706
rect 5632 26590 5637 26642
rect 5637 26590 5684 26642
rect 5700 26590 5752 26642
rect 5768 26590 5815 26642
rect 5815 26590 5820 26642
rect 5632 26526 5637 26578
rect 5637 26526 5684 26578
rect 5700 26526 5752 26578
rect 5768 26526 5815 26578
rect 5815 26526 5820 26578
rect 5632 26462 5637 26514
rect 5637 26462 5684 26514
rect 5700 26462 5752 26514
rect 5768 26462 5815 26514
rect 5815 26462 5820 26514
rect 5632 26398 5637 26450
rect 5637 26398 5684 26450
rect 5700 26398 5752 26450
rect 5768 26398 5815 26450
rect 5815 26398 5820 26450
rect 5632 26334 5637 26386
rect 5637 26334 5684 26386
rect 5700 26334 5752 26386
rect 5768 26334 5815 26386
rect 5815 26334 5820 26386
rect 5632 26270 5637 26322
rect 5637 26270 5684 26322
rect 5700 26270 5752 26322
rect 5768 26270 5815 26322
rect 5815 26270 5820 26322
rect 5632 26206 5637 26258
rect 5637 26206 5684 26258
rect 5700 26206 5752 26258
rect 5768 26206 5815 26258
rect 5815 26206 5820 26258
rect 5632 26142 5637 26194
rect 5637 26142 5684 26194
rect 5700 26142 5752 26194
rect 5768 26142 5815 26194
rect 5815 26142 5820 26194
rect 5632 26077 5637 26129
rect 5637 26077 5684 26129
rect 5700 26077 5752 26129
rect 5768 26077 5815 26129
rect 5815 26077 5820 26129
rect 5632 26012 5637 26064
rect 5637 26012 5684 26064
rect 5700 26012 5752 26064
rect 5768 26012 5815 26064
rect 5815 26012 5820 26064
rect 5632 25947 5637 25999
rect 5637 25947 5684 25999
rect 5700 25947 5752 25999
rect 5768 25947 5815 25999
rect 5815 25947 5820 25999
rect 5632 25882 5637 25934
rect 5637 25882 5684 25934
rect 5700 25882 5752 25934
rect 5768 25882 5815 25934
rect 5815 25882 5820 25934
rect 5632 25817 5637 25869
rect 5637 25817 5684 25869
rect 5700 25817 5752 25869
rect 5768 25817 5815 25869
rect 5815 25817 5820 25869
rect 5632 25752 5637 25804
rect 5637 25752 5684 25804
rect 5700 25752 5752 25804
rect 5768 25752 5815 25804
rect 5815 25752 5820 25804
rect 5632 25687 5637 25739
rect 5637 25687 5684 25739
rect 5700 25687 5752 25739
rect 5768 25687 5815 25739
rect 5815 25687 5820 25739
rect 5632 25622 5637 25674
rect 5637 25622 5684 25674
rect 5700 25622 5752 25674
rect 5768 25622 5815 25674
rect 5815 25622 5820 25674
rect 5632 25557 5637 25609
rect 5637 25557 5684 25609
rect 5700 25557 5752 25609
rect 5768 25557 5815 25609
rect 5815 25557 5820 25609
rect 5632 25492 5637 25544
rect 5637 25492 5684 25544
rect 5700 25492 5752 25544
rect 5768 25492 5815 25544
rect 5815 25492 5820 25544
rect 5632 25427 5637 25479
rect 5637 25427 5684 25479
rect 5700 25427 5752 25479
rect 5768 25427 5815 25479
rect 5815 25427 5820 25479
rect 5632 25362 5637 25414
rect 5637 25362 5684 25414
rect 5700 25362 5752 25414
rect 5768 25362 5815 25414
rect 5815 25362 5820 25414
rect 5632 22438 5637 22490
rect 5637 22438 5684 22490
rect 5700 22438 5752 22490
rect 5768 22438 5815 22490
rect 5815 22438 5820 22490
rect 5632 22374 5637 22426
rect 5637 22374 5684 22426
rect 5700 22374 5752 22426
rect 5768 22374 5815 22426
rect 5815 22374 5820 22426
rect 5632 22310 5637 22362
rect 5637 22310 5684 22362
rect 5700 22310 5752 22362
rect 5768 22310 5815 22362
rect 5815 22310 5820 22362
rect 5632 22246 5637 22298
rect 5637 22246 5684 22298
rect 5700 22246 5752 22298
rect 5768 22246 5815 22298
rect 5815 22246 5820 22298
rect 5632 22182 5637 22234
rect 5637 22182 5684 22234
rect 5700 22182 5752 22234
rect 5768 22182 5815 22234
rect 5815 22182 5820 22234
rect 5632 22118 5637 22170
rect 5637 22118 5684 22170
rect 5700 22118 5752 22170
rect 5768 22118 5815 22170
rect 5815 22118 5820 22170
rect 5632 22054 5637 22106
rect 5637 22054 5684 22106
rect 5700 22054 5752 22106
rect 5768 22054 5815 22106
rect 5815 22054 5820 22106
rect 5632 21990 5637 22042
rect 5637 21990 5684 22042
rect 5700 21990 5752 22042
rect 5768 21990 5815 22042
rect 5815 21990 5820 22042
rect 5632 21926 5637 21978
rect 5637 21926 5684 21978
rect 5700 21926 5752 21978
rect 5768 21926 5815 21978
rect 5815 21926 5820 21978
rect 5632 21862 5637 21914
rect 5637 21862 5684 21914
rect 5700 21862 5752 21914
rect 5768 21862 5815 21914
rect 5815 21862 5820 21914
rect 5632 21798 5637 21850
rect 5637 21798 5684 21850
rect 5700 21798 5752 21850
rect 5768 21798 5815 21850
rect 5815 21798 5820 21850
rect 5632 21734 5637 21786
rect 5637 21734 5684 21786
rect 5700 21734 5752 21786
rect 5768 21734 5815 21786
rect 5815 21734 5820 21786
rect 5632 21670 5637 21722
rect 5637 21670 5684 21722
rect 5700 21670 5752 21722
rect 5768 21670 5815 21722
rect 5815 21670 5820 21722
rect 5632 21606 5637 21658
rect 5637 21606 5684 21658
rect 5700 21606 5752 21658
rect 5768 21606 5815 21658
rect 5815 21606 5820 21658
rect 5632 21542 5637 21594
rect 5637 21542 5684 21594
rect 5700 21542 5752 21594
rect 5768 21542 5815 21594
rect 5815 21542 5820 21594
rect 5632 21477 5637 21529
rect 5637 21477 5684 21529
rect 5700 21477 5752 21529
rect 5768 21477 5815 21529
rect 5815 21477 5820 21529
rect 5632 21412 5637 21464
rect 5637 21412 5684 21464
rect 5700 21412 5752 21464
rect 5768 21412 5815 21464
rect 5815 21412 5820 21464
rect 5632 21347 5637 21399
rect 5637 21347 5684 21399
rect 5700 21347 5752 21399
rect 5768 21347 5815 21399
rect 5815 21347 5820 21399
rect 5632 21282 5637 21334
rect 5637 21282 5684 21334
rect 5700 21282 5752 21334
rect 5768 21282 5815 21334
rect 5815 21282 5820 21334
rect 5632 21217 5637 21269
rect 5637 21217 5684 21269
rect 5700 21217 5752 21269
rect 5768 21217 5815 21269
rect 5815 21217 5820 21269
rect 5632 21152 5637 21204
rect 5637 21152 5684 21204
rect 5700 21152 5752 21204
rect 5768 21152 5815 21204
rect 5815 21152 5820 21204
rect 5632 21087 5637 21139
rect 5637 21087 5684 21139
rect 5700 21087 5752 21139
rect 5768 21087 5815 21139
rect 5815 21087 5820 21139
rect 5632 21022 5637 21074
rect 5637 21022 5684 21074
rect 5700 21022 5752 21074
rect 5768 21022 5815 21074
rect 5815 21022 5820 21074
rect 5632 20957 5637 21009
rect 5637 20957 5684 21009
rect 5700 20957 5752 21009
rect 5768 20957 5815 21009
rect 5815 20957 5820 21009
rect 5632 20892 5637 20944
rect 5637 20892 5684 20944
rect 5700 20892 5752 20944
rect 5768 20892 5815 20944
rect 5815 20892 5820 20944
rect 5632 20827 5637 20879
rect 5637 20827 5684 20879
rect 5700 20827 5752 20879
rect 5768 20827 5815 20879
rect 5815 20827 5820 20879
rect 5632 20762 5637 20814
rect 5637 20762 5684 20814
rect 5700 20762 5752 20814
rect 5768 20762 5815 20814
rect 5815 20762 5820 20814
rect 5632 17838 5637 17890
rect 5637 17838 5684 17890
rect 5700 17838 5752 17890
rect 5768 17838 5815 17890
rect 5815 17838 5820 17890
rect 5632 17774 5637 17826
rect 5637 17774 5684 17826
rect 5700 17774 5752 17826
rect 5768 17774 5815 17826
rect 5815 17774 5820 17826
rect 5632 17710 5637 17762
rect 5637 17710 5684 17762
rect 5700 17710 5752 17762
rect 5768 17710 5815 17762
rect 5815 17710 5820 17762
rect 5632 17646 5637 17698
rect 5637 17646 5684 17698
rect 5700 17646 5752 17698
rect 5768 17646 5815 17698
rect 5815 17646 5820 17698
rect 5632 17582 5637 17634
rect 5637 17582 5684 17634
rect 5700 17582 5752 17634
rect 5768 17582 5815 17634
rect 5815 17582 5820 17634
rect 5632 17518 5637 17570
rect 5637 17518 5684 17570
rect 5700 17518 5752 17570
rect 5768 17518 5815 17570
rect 5815 17518 5820 17570
rect 5632 17454 5637 17506
rect 5637 17454 5684 17506
rect 5700 17454 5752 17506
rect 5768 17454 5815 17506
rect 5815 17454 5820 17506
rect 5632 17390 5637 17442
rect 5637 17390 5684 17442
rect 5700 17390 5752 17442
rect 5768 17390 5815 17442
rect 5815 17390 5820 17442
rect 5632 17326 5637 17378
rect 5637 17326 5684 17378
rect 5700 17326 5752 17378
rect 5768 17326 5815 17378
rect 5815 17326 5820 17378
rect 5632 17262 5637 17314
rect 5637 17262 5684 17314
rect 5700 17262 5752 17314
rect 5768 17262 5815 17314
rect 5815 17262 5820 17314
rect 5632 17198 5637 17250
rect 5637 17198 5684 17250
rect 5700 17198 5752 17250
rect 5768 17198 5815 17250
rect 5815 17198 5820 17250
rect 5632 17134 5637 17186
rect 5637 17134 5684 17186
rect 5700 17134 5752 17186
rect 5768 17134 5815 17186
rect 5815 17134 5820 17186
rect 5632 17070 5637 17122
rect 5637 17070 5684 17122
rect 5700 17070 5752 17122
rect 5768 17070 5815 17122
rect 5815 17070 5820 17122
rect 5632 17006 5637 17058
rect 5637 17006 5684 17058
rect 5700 17006 5752 17058
rect 5768 17006 5815 17058
rect 5815 17006 5820 17058
rect 5632 16942 5637 16994
rect 5637 16942 5684 16994
rect 5700 16942 5752 16994
rect 5768 16942 5815 16994
rect 5815 16942 5820 16994
rect 5632 16877 5637 16929
rect 5637 16877 5684 16929
rect 5700 16877 5752 16929
rect 5768 16877 5815 16929
rect 5815 16877 5820 16929
rect 5632 16812 5637 16864
rect 5637 16812 5684 16864
rect 5700 16812 5752 16864
rect 5768 16812 5815 16864
rect 5815 16812 5820 16864
rect 5632 16747 5637 16799
rect 5637 16747 5684 16799
rect 5700 16747 5752 16799
rect 5768 16747 5815 16799
rect 5815 16747 5820 16799
rect 5632 16682 5637 16734
rect 5637 16682 5684 16734
rect 5700 16682 5752 16734
rect 5768 16682 5815 16734
rect 5815 16682 5820 16734
rect 5632 16617 5637 16669
rect 5637 16617 5684 16669
rect 5700 16617 5752 16669
rect 5768 16617 5815 16669
rect 5815 16617 5820 16669
rect 5632 16552 5637 16604
rect 5637 16552 5684 16604
rect 5700 16552 5752 16604
rect 5768 16552 5815 16604
rect 5815 16552 5820 16604
rect 5632 16487 5637 16539
rect 5637 16487 5684 16539
rect 5700 16487 5752 16539
rect 5768 16487 5815 16539
rect 5815 16487 5820 16539
rect 5632 16422 5637 16474
rect 5637 16422 5684 16474
rect 5700 16422 5752 16474
rect 5768 16422 5815 16474
rect 5815 16422 5820 16474
rect 5632 16357 5637 16409
rect 5637 16357 5684 16409
rect 5700 16357 5752 16409
rect 5768 16357 5815 16409
rect 5815 16357 5820 16409
rect 5632 16292 5637 16344
rect 5637 16292 5684 16344
rect 5700 16292 5752 16344
rect 5768 16292 5815 16344
rect 5815 16292 5820 16344
rect 5632 16227 5637 16279
rect 5637 16227 5684 16279
rect 5700 16227 5752 16279
rect 5768 16227 5815 16279
rect 5815 16227 5820 16279
rect 5632 16162 5637 16214
rect 5637 16162 5684 16214
rect 5700 16162 5752 16214
rect 5768 16162 5815 16214
rect 5815 16162 5820 16214
rect 5632 13238 5637 13290
rect 5637 13238 5684 13290
rect 5700 13238 5752 13290
rect 5768 13238 5815 13290
rect 5815 13238 5820 13290
rect 5632 13174 5637 13226
rect 5637 13174 5684 13226
rect 5700 13174 5752 13226
rect 5768 13174 5815 13226
rect 5815 13174 5820 13226
rect 5632 13110 5637 13162
rect 5637 13110 5684 13162
rect 5700 13110 5752 13162
rect 5768 13110 5815 13162
rect 5815 13110 5820 13162
rect 5632 13046 5637 13098
rect 5637 13046 5684 13098
rect 5700 13046 5752 13098
rect 5768 13046 5815 13098
rect 5815 13046 5820 13098
rect 5632 12982 5637 13034
rect 5637 12982 5684 13034
rect 5700 12982 5752 13034
rect 5768 12982 5815 13034
rect 5815 12982 5820 13034
rect 5632 12918 5637 12970
rect 5637 12918 5684 12970
rect 5700 12918 5752 12970
rect 5768 12918 5815 12970
rect 5815 12918 5820 12970
rect 5632 12854 5637 12906
rect 5637 12854 5684 12906
rect 5700 12854 5752 12906
rect 5768 12854 5815 12906
rect 5815 12854 5820 12906
rect 5632 12790 5637 12842
rect 5637 12790 5684 12842
rect 5700 12790 5752 12842
rect 5768 12790 5815 12842
rect 5815 12790 5820 12842
rect 5632 12726 5637 12778
rect 5637 12726 5684 12778
rect 5700 12726 5752 12778
rect 5768 12726 5815 12778
rect 5815 12726 5820 12778
rect 5632 12662 5637 12714
rect 5637 12662 5684 12714
rect 5700 12662 5752 12714
rect 5768 12662 5815 12714
rect 5815 12662 5820 12714
rect 5632 12598 5637 12650
rect 5637 12598 5684 12650
rect 5700 12598 5752 12650
rect 5768 12598 5815 12650
rect 5815 12598 5820 12650
rect 5632 12534 5637 12586
rect 5637 12534 5684 12586
rect 5700 12534 5752 12586
rect 5768 12534 5815 12586
rect 5815 12534 5820 12586
rect 5632 12470 5637 12522
rect 5637 12470 5684 12522
rect 5700 12470 5752 12522
rect 5768 12470 5815 12522
rect 5815 12470 5820 12522
rect 5632 12406 5637 12458
rect 5637 12406 5684 12458
rect 5700 12406 5752 12458
rect 5768 12406 5815 12458
rect 5815 12406 5820 12458
rect 5632 12342 5637 12394
rect 5637 12342 5684 12394
rect 5700 12342 5752 12394
rect 5768 12342 5815 12394
rect 5815 12342 5820 12394
rect 5632 12277 5637 12329
rect 5637 12277 5684 12329
rect 5700 12277 5752 12329
rect 5768 12277 5815 12329
rect 5815 12277 5820 12329
rect 5632 12212 5637 12264
rect 5637 12212 5684 12264
rect 5700 12212 5752 12264
rect 5768 12212 5815 12264
rect 5815 12212 5820 12264
rect 5632 12147 5637 12199
rect 5637 12147 5684 12199
rect 5700 12147 5752 12199
rect 5768 12147 5815 12199
rect 5815 12147 5820 12199
rect 5632 12082 5637 12134
rect 5637 12082 5684 12134
rect 5700 12082 5752 12134
rect 5768 12082 5815 12134
rect 5815 12082 5820 12134
rect 5632 12017 5637 12069
rect 5637 12017 5684 12069
rect 5700 12017 5752 12069
rect 5768 12017 5815 12069
rect 5815 12017 5820 12069
rect 5632 11952 5637 12004
rect 5637 11952 5684 12004
rect 5700 11952 5752 12004
rect 5768 11952 5815 12004
rect 5815 11952 5820 12004
rect 5632 11887 5637 11939
rect 5637 11887 5684 11939
rect 5700 11887 5752 11939
rect 5768 11887 5815 11939
rect 5815 11887 5820 11939
rect 5632 11822 5637 11874
rect 5637 11822 5684 11874
rect 5700 11822 5752 11874
rect 5768 11822 5815 11874
rect 5815 11822 5820 11874
rect 5632 11757 5637 11809
rect 5637 11757 5684 11809
rect 5700 11757 5752 11809
rect 5768 11757 5815 11809
rect 5815 11757 5820 11809
rect 5632 11692 5637 11744
rect 5637 11692 5684 11744
rect 5700 11692 5752 11744
rect 5768 11692 5815 11744
rect 5815 11692 5820 11744
rect 5632 11627 5637 11679
rect 5637 11627 5684 11679
rect 5700 11627 5752 11679
rect 5768 11627 5815 11679
rect 5815 11627 5820 11679
rect 5632 11562 5637 11614
rect 5637 11562 5684 11614
rect 5700 11562 5752 11614
rect 5768 11562 5815 11614
rect 5815 11562 5820 11614
rect 6121 37945 6173 37997
rect 6199 37945 6251 37997
rect 6121 37877 6173 37929
rect 6199 37877 6251 37929
rect 6121 37809 6173 37861
rect 6199 37809 6251 37861
rect 6121 37741 6173 37793
rect 6199 37741 6251 37793
rect 6121 37673 6173 37725
rect 6199 37673 6251 37725
rect 6121 37605 6173 37657
rect 6199 37605 6251 37657
rect 6121 37537 6173 37589
rect 6199 37537 6251 37589
rect 6121 37469 6173 37521
rect 6199 37469 6251 37521
rect 6121 37401 6173 37453
rect 6199 37401 6251 37453
rect 6121 37333 6173 37385
rect 6199 37333 6251 37385
rect 6121 37266 6173 37318
rect 6199 37266 6251 37318
rect 6121 37199 6173 37251
rect 6199 37199 6251 37251
rect 6121 37132 6173 37184
rect 6199 37132 6251 37184
rect 6121 37065 6173 37117
rect 6199 37065 6251 37117
rect 6121 34173 6173 34225
rect 6199 34173 6251 34225
rect 6121 34109 6173 34161
rect 6199 34109 6251 34161
rect 6121 34045 6173 34097
rect 6199 34045 6251 34097
rect 6121 33981 6173 34033
rect 6199 33981 6251 34033
rect 6121 33917 6173 33969
rect 6199 33917 6251 33969
rect 6121 33853 6173 33905
rect 6199 33853 6251 33905
rect 6121 33789 6173 33841
rect 6199 33789 6251 33841
rect 6121 33725 6173 33777
rect 6199 33725 6251 33777
rect 6121 33661 6173 33713
rect 6199 33661 6251 33713
rect 6121 33597 6173 33649
rect 6199 33597 6251 33649
rect 6121 33533 6173 33585
rect 6199 33533 6251 33585
rect 6121 33469 6173 33521
rect 6199 33469 6251 33521
rect 6121 33405 6173 33457
rect 6199 33405 6251 33457
rect 6121 33341 6173 33393
rect 6199 33341 6251 33393
rect 6121 33277 6173 33329
rect 6199 33277 6251 33329
rect 6121 33212 6173 33264
rect 6199 33212 6251 33264
rect 6121 33147 6173 33199
rect 6199 33147 6251 33199
rect 6121 33082 6173 33134
rect 6199 33082 6251 33134
rect 6121 33017 6173 33069
rect 6199 33017 6251 33069
rect 6121 32952 6173 33004
rect 6199 32952 6251 33004
rect 6121 32887 6173 32939
rect 6199 32887 6251 32939
rect 6121 32822 6173 32874
rect 6199 32822 6251 32874
rect 6121 32757 6173 32809
rect 6199 32757 6251 32809
rect 6121 32692 6173 32744
rect 6199 32692 6251 32744
rect 6121 32627 6173 32679
rect 6199 32627 6251 32679
rect 6121 32562 6173 32614
rect 6199 32562 6251 32614
rect 6121 32497 6173 32549
rect 6199 32497 6251 32549
rect 6121 29573 6173 29625
rect 6199 29573 6251 29625
rect 6121 29509 6173 29561
rect 6199 29509 6251 29561
rect 6121 29445 6173 29497
rect 6199 29445 6251 29497
rect 6121 29381 6173 29433
rect 6199 29381 6251 29433
rect 6121 29317 6173 29369
rect 6199 29317 6251 29369
rect 6121 29253 6173 29305
rect 6199 29253 6251 29305
rect 6121 29189 6173 29241
rect 6199 29189 6251 29241
rect 6121 29125 6173 29177
rect 6199 29125 6251 29177
rect 6121 29061 6173 29113
rect 6199 29061 6251 29113
rect 6121 28997 6173 29049
rect 6199 28997 6251 29049
rect 6121 28933 6173 28985
rect 6199 28933 6251 28985
rect 6121 28869 6173 28921
rect 6199 28869 6251 28921
rect 6121 28805 6173 28857
rect 6199 28805 6251 28857
rect 6121 28741 6173 28793
rect 6199 28741 6251 28793
rect 6121 28677 6173 28729
rect 6199 28677 6251 28729
rect 6121 28612 6173 28664
rect 6199 28612 6251 28664
rect 6121 28547 6173 28599
rect 6199 28547 6251 28599
rect 6121 28482 6173 28534
rect 6199 28482 6251 28534
rect 6121 28417 6173 28469
rect 6199 28417 6251 28469
rect 6121 28352 6173 28404
rect 6199 28352 6251 28404
rect 6121 28287 6173 28339
rect 6199 28287 6251 28339
rect 6121 28222 6173 28274
rect 6199 28222 6251 28274
rect 6121 28157 6173 28209
rect 6199 28157 6251 28209
rect 6121 28092 6173 28144
rect 6199 28092 6251 28144
rect 6121 28027 6173 28079
rect 6199 28027 6251 28079
rect 6121 27962 6173 28014
rect 6199 27962 6251 28014
rect 6121 27897 6173 27949
rect 6199 27897 6251 27949
rect 6121 24973 6173 25025
rect 6199 24973 6251 25025
rect 6121 24909 6173 24961
rect 6199 24909 6251 24961
rect 6121 24845 6173 24897
rect 6199 24845 6251 24897
rect 6121 24781 6173 24833
rect 6199 24781 6251 24833
rect 6121 24717 6173 24769
rect 6199 24717 6251 24769
rect 6121 24653 6173 24705
rect 6199 24653 6251 24705
rect 6121 24589 6173 24641
rect 6199 24589 6251 24641
rect 6121 24525 6173 24577
rect 6199 24525 6251 24577
rect 6121 24461 6173 24513
rect 6199 24461 6251 24513
rect 6121 24397 6173 24449
rect 6199 24397 6251 24449
rect 6121 24333 6173 24385
rect 6199 24333 6251 24385
rect 6121 24269 6173 24321
rect 6199 24269 6251 24321
rect 6121 24205 6173 24257
rect 6199 24205 6251 24257
rect 6121 24141 6173 24193
rect 6199 24141 6251 24193
rect 6121 24077 6173 24129
rect 6199 24077 6251 24129
rect 6121 24012 6173 24064
rect 6199 24012 6251 24064
rect 6121 23947 6173 23999
rect 6199 23947 6251 23999
rect 6121 23882 6173 23934
rect 6199 23882 6251 23934
rect 6121 23817 6173 23869
rect 6199 23817 6251 23869
rect 6121 23752 6173 23804
rect 6199 23752 6251 23804
rect 6121 23687 6173 23739
rect 6199 23687 6251 23739
rect 6121 23622 6173 23674
rect 6199 23622 6251 23674
rect 6121 23557 6173 23609
rect 6199 23557 6251 23609
rect 6121 23492 6173 23544
rect 6199 23492 6251 23544
rect 6121 23427 6173 23479
rect 6199 23427 6251 23479
rect 6121 23362 6173 23414
rect 6199 23362 6251 23414
rect 6121 23297 6173 23349
rect 6199 23297 6251 23349
rect 6121 20373 6173 20425
rect 6199 20373 6251 20425
rect 6121 20309 6173 20361
rect 6199 20309 6251 20361
rect 6121 20245 6173 20297
rect 6199 20245 6251 20297
rect 6121 20181 6173 20233
rect 6199 20181 6251 20233
rect 6121 20117 6173 20169
rect 6199 20117 6251 20169
rect 6121 20053 6173 20105
rect 6199 20053 6251 20105
rect 6121 19989 6173 20041
rect 6199 19989 6251 20041
rect 6121 19925 6173 19977
rect 6199 19925 6251 19977
rect 6121 19861 6173 19913
rect 6199 19861 6251 19913
rect 6121 19797 6173 19849
rect 6199 19797 6251 19849
rect 6121 19733 6173 19785
rect 6199 19733 6251 19785
rect 6121 19669 6173 19721
rect 6199 19669 6251 19721
rect 6121 19605 6173 19657
rect 6199 19605 6251 19657
rect 6121 19541 6173 19593
rect 6199 19541 6251 19593
rect 6121 19477 6173 19529
rect 6199 19477 6251 19529
rect 6121 19412 6173 19464
rect 6199 19412 6251 19464
rect 6121 19347 6173 19399
rect 6199 19347 6251 19399
rect 6121 19282 6173 19334
rect 6199 19282 6251 19334
rect 6121 19217 6173 19269
rect 6199 19217 6251 19269
rect 6121 19152 6173 19204
rect 6199 19152 6251 19204
rect 6121 19087 6173 19139
rect 6199 19087 6251 19139
rect 6121 19022 6173 19074
rect 6199 19022 6251 19074
rect 6121 18957 6173 19009
rect 6199 18957 6251 19009
rect 6121 18892 6173 18944
rect 6199 18892 6251 18944
rect 6121 18827 6173 18879
rect 6199 18827 6251 18879
rect 6121 18762 6173 18814
rect 6199 18762 6251 18814
rect 6121 18697 6173 18749
rect 6199 18697 6251 18749
rect 6121 15773 6173 15825
rect 6199 15773 6251 15825
rect 6121 15709 6173 15761
rect 6199 15709 6251 15761
rect 6121 15645 6173 15697
rect 6199 15645 6251 15697
rect 6121 15581 6173 15633
rect 6199 15581 6251 15633
rect 6121 15517 6173 15569
rect 6199 15517 6251 15569
rect 6121 15453 6173 15505
rect 6199 15453 6251 15505
rect 6121 15389 6173 15441
rect 6199 15389 6251 15441
rect 6121 15325 6173 15377
rect 6199 15325 6251 15377
rect 6121 15261 6173 15313
rect 6199 15261 6251 15313
rect 6121 15197 6173 15249
rect 6199 15197 6251 15249
rect 6121 15133 6173 15185
rect 6199 15133 6251 15185
rect 6121 15069 6173 15121
rect 6199 15069 6251 15121
rect 6121 15005 6173 15057
rect 6199 15005 6251 15057
rect 6121 14941 6173 14993
rect 6199 14941 6251 14993
rect 6121 14877 6173 14929
rect 6199 14877 6251 14929
rect 6121 14812 6173 14864
rect 6199 14812 6251 14864
rect 6121 14747 6173 14799
rect 6199 14747 6251 14799
rect 6121 14682 6173 14734
rect 6199 14682 6251 14734
rect 6121 14617 6173 14669
rect 6199 14617 6251 14669
rect 6121 14552 6173 14604
rect 6199 14552 6251 14604
rect 6121 14487 6173 14539
rect 6199 14487 6251 14539
rect 6121 14422 6173 14474
rect 6199 14422 6251 14474
rect 6121 14357 6173 14409
rect 6199 14357 6251 14409
rect 6121 14292 6173 14344
rect 6199 14292 6251 14344
rect 6121 14227 6173 14279
rect 6199 14227 6251 14279
rect 6121 14162 6173 14214
rect 6199 14162 6251 14214
rect 6121 14097 6173 14149
rect 6199 14097 6251 14149
rect 6121 11173 6173 11225
rect 6199 11173 6251 11225
rect 6121 11109 6173 11161
rect 6199 11109 6251 11161
rect 6121 11045 6173 11097
rect 6199 11045 6251 11097
rect 6121 10981 6173 11033
rect 6199 10981 6251 11033
rect 6121 10917 6173 10969
rect 6199 10917 6251 10969
rect 6121 10853 6173 10905
rect 6199 10853 6251 10905
rect 6121 10789 6173 10841
rect 6199 10789 6251 10841
rect 6121 10725 6173 10777
rect 6199 10725 6251 10777
rect 6121 10661 6173 10713
rect 6199 10661 6251 10713
rect 6121 10597 6173 10649
rect 6199 10597 6251 10649
rect 6121 10533 6173 10585
rect 6199 10533 6251 10585
rect 6121 10469 6173 10521
rect 6199 10469 6251 10521
rect 6121 10405 6173 10457
rect 6199 10405 6251 10457
rect 6121 10341 6173 10393
rect 6199 10341 6251 10393
rect 6121 10277 6173 10329
rect 6199 10277 6251 10329
rect 6121 10212 6173 10264
rect 6199 10212 6251 10264
rect 6121 10147 6173 10199
rect 6199 10147 6251 10199
rect 6121 10082 6173 10134
rect 6199 10082 6251 10134
rect 6121 10017 6173 10069
rect 6199 10017 6251 10069
rect 6121 9952 6173 10004
rect 6199 9952 6251 10004
rect 6121 9887 6173 9939
rect 6199 9887 6251 9939
rect 6121 9822 6173 9874
rect 6199 9822 6251 9874
rect 6121 9757 6173 9809
rect 6199 9757 6251 9809
rect 6121 9692 6173 9744
rect 6199 9692 6251 9744
rect 6121 9627 6173 9679
rect 6199 9627 6251 9679
rect 6121 9562 6173 9614
rect 6199 9562 6251 9614
rect 6121 9497 6173 9549
rect 6199 9497 6251 9549
rect 6552 36238 6557 36290
rect 6557 36238 6604 36290
rect 6620 36238 6672 36290
rect 6688 36238 6735 36290
rect 6735 36238 6740 36290
rect 6552 36174 6557 36226
rect 6557 36174 6604 36226
rect 6620 36174 6672 36226
rect 6688 36174 6735 36226
rect 6735 36174 6740 36226
rect 6552 36110 6557 36162
rect 6557 36110 6604 36162
rect 6620 36110 6672 36162
rect 6688 36110 6735 36162
rect 6735 36110 6740 36162
rect 6552 36046 6557 36098
rect 6557 36046 6604 36098
rect 6620 36046 6672 36098
rect 6688 36046 6735 36098
rect 6735 36046 6740 36098
rect 6552 35982 6557 36034
rect 6557 35982 6604 36034
rect 6620 35982 6672 36034
rect 6688 35982 6735 36034
rect 6735 35982 6740 36034
rect 6552 35918 6557 35970
rect 6557 35918 6604 35970
rect 6620 35918 6672 35970
rect 6688 35918 6735 35970
rect 6735 35918 6740 35970
rect 6552 35854 6557 35906
rect 6557 35854 6604 35906
rect 6620 35854 6672 35906
rect 6688 35854 6735 35906
rect 6735 35854 6740 35906
rect 6552 35790 6557 35842
rect 6557 35790 6604 35842
rect 6620 35790 6672 35842
rect 6688 35790 6735 35842
rect 6735 35790 6740 35842
rect 6552 35726 6557 35778
rect 6557 35726 6604 35778
rect 6620 35726 6672 35778
rect 6688 35726 6735 35778
rect 6735 35726 6740 35778
rect 6552 35662 6557 35714
rect 6557 35662 6604 35714
rect 6620 35662 6672 35714
rect 6688 35662 6735 35714
rect 6735 35662 6740 35714
rect 6552 35598 6557 35650
rect 6557 35598 6604 35650
rect 6620 35598 6672 35650
rect 6688 35598 6735 35650
rect 6735 35598 6740 35650
rect 6552 35534 6557 35586
rect 6557 35534 6604 35586
rect 6620 35534 6672 35586
rect 6688 35534 6735 35586
rect 6735 35534 6740 35586
rect 6552 35470 6557 35522
rect 6557 35470 6604 35522
rect 6620 35470 6672 35522
rect 6688 35470 6735 35522
rect 6735 35470 6740 35522
rect 6552 35406 6557 35458
rect 6557 35406 6604 35458
rect 6620 35406 6672 35458
rect 6688 35406 6735 35458
rect 6735 35406 6740 35458
rect 6552 35342 6557 35394
rect 6557 35342 6604 35394
rect 6620 35342 6672 35394
rect 6688 35342 6735 35394
rect 6735 35342 6740 35394
rect 6552 35277 6557 35329
rect 6557 35277 6604 35329
rect 6620 35277 6672 35329
rect 6688 35277 6735 35329
rect 6735 35277 6740 35329
rect 6552 35212 6557 35264
rect 6557 35212 6604 35264
rect 6620 35212 6672 35264
rect 6688 35212 6735 35264
rect 6735 35212 6740 35264
rect 6552 35147 6557 35199
rect 6557 35147 6604 35199
rect 6620 35147 6672 35199
rect 6688 35147 6735 35199
rect 6735 35147 6740 35199
rect 6552 35082 6557 35134
rect 6557 35082 6604 35134
rect 6620 35082 6672 35134
rect 6688 35082 6735 35134
rect 6735 35082 6740 35134
rect 6552 35017 6557 35069
rect 6557 35017 6604 35069
rect 6620 35017 6672 35069
rect 6688 35017 6735 35069
rect 6735 35017 6740 35069
rect 6552 34952 6557 35004
rect 6557 34952 6604 35004
rect 6620 34952 6672 35004
rect 6688 34952 6735 35004
rect 6735 34952 6740 35004
rect 6552 34887 6557 34939
rect 6557 34887 6604 34939
rect 6620 34887 6672 34939
rect 6688 34887 6735 34939
rect 6735 34887 6740 34939
rect 6552 34822 6557 34874
rect 6557 34822 6604 34874
rect 6620 34822 6672 34874
rect 6688 34822 6735 34874
rect 6735 34822 6740 34874
rect 6552 34757 6557 34809
rect 6557 34757 6604 34809
rect 6620 34757 6672 34809
rect 6688 34757 6735 34809
rect 6735 34757 6740 34809
rect 6552 34692 6557 34744
rect 6557 34692 6604 34744
rect 6620 34692 6672 34744
rect 6688 34692 6735 34744
rect 6735 34692 6740 34744
rect 6552 34627 6557 34679
rect 6557 34627 6604 34679
rect 6620 34627 6672 34679
rect 6688 34627 6735 34679
rect 6735 34627 6740 34679
rect 6552 34562 6557 34614
rect 6557 34562 6604 34614
rect 6620 34562 6672 34614
rect 6688 34562 6735 34614
rect 6735 34562 6740 34614
rect 6552 31638 6557 31690
rect 6557 31638 6604 31690
rect 6620 31638 6672 31690
rect 6688 31638 6735 31690
rect 6735 31638 6740 31690
rect 6552 31574 6557 31626
rect 6557 31574 6604 31626
rect 6620 31574 6672 31626
rect 6688 31574 6735 31626
rect 6735 31574 6740 31626
rect 6552 31510 6557 31562
rect 6557 31510 6604 31562
rect 6620 31510 6672 31562
rect 6688 31510 6735 31562
rect 6735 31510 6740 31562
rect 6552 31446 6557 31498
rect 6557 31446 6604 31498
rect 6620 31446 6672 31498
rect 6688 31446 6735 31498
rect 6735 31446 6740 31498
rect 6552 31382 6557 31434
rect 6557 31382 6604 31434
rect 6620 31382 6672 31434
rect 6688 31382 6735 31434
rect 6735 31382 6740 31434
rect 6552 31318 6557 31370
rect 6557 31318 6604 31370
rect 6620 31318 6672 31370
rect 6688 31318 6735 31370
rect 6735 31318 6740 31370
rect 6552 31254 6557 31306
rect 6557 31254 6604 31306
rect 6620 31254 6672 31306
rect 6688 31254 6735 31306
rect 6735 31254 6740 31306
rect 6552 31190 6557 31242
rect 6557 31190 6604 31242
rect 6620 31190 6672 31242
rect 6688 31190 6735 31242
rect 6735 31190 6740 31242
rect 6552 31126 6557 31178
rect 6557 31126 6604 31178
rect 6620 31126 6672 31178
rect 6688 31126 6735 31178
rect 6735 31126 6740 31178
rect 6552 31062 6557 31114
rect 6557 31062 6604 31114
rect 6620 31062 6672 31114
rect 6688 31062 6735 31114
rect 6735 31062 6740 31114
rect 6552 30998 6557 31050
rect 6557 30998 6604 31050
rect 6620 30998 6672 31050
rect 6688 30998 6735 31050
rect 6735 30998 6740 31050
rect 6552 30934 6557 30986
rect 6557 30934 6604 30986
rect 6620 30934 6672 30986
rect 6688 30934 6735 30986
rect 6735 30934 6740 30986
rect 6552 30870 6557 30922
rect 6557 30870 6604 30922
rect 6620 30870 6672 30922
rect 6688 30870 6735 30922
rect 6735 30870 6740 30922
rect 6552 30806 6557 30858
rect 6557 30806 6604 30858
rect 6620 30806 6672 30858
rect 6688 30806 6735 30858
rect 6735 30806 6740 30858
rect 6552 30742 6557 30794
rect 6557 30742 6604 30794
rect 6620 30742 6672 30794
rect 6688 30742 6735 30794
rect 6735 30742 6740 30794
rect 6552 30677 6557 30729
rect 6557 30677 6604 30729
rect 6620 30677 6672 30729
rect 6688 30677 6735 30729
rect 6735 30677 6740 30729
rect 6552 30612 6557 30664
rect 6557 30612 6604 30664
rect 6620 30612 6672 30664
rect 6688 30612 6735 30664
rect 6735 30612 6740 30664
rect 6552 30547 6557 30599
rect 6557 30547 6604 30599
rect 6620 30547 6672 30599
rect 6688 30547 6735 30599
rect 6735 30547 6740 30599
rect 6552 30482 6557 30534
rect 6557 30482 6604 30534
rect 6620 30482 6672 30534
rect 6688 30482 6735 30534
rect 6735 30482 6740 30534
rect 6552 30417 6557 30469
rect 6557 30417 6604 30469
rect 6620 30417 6672 30469
rect 6688 30417 6735 30469
rect 6735 30417 6740 30469
rect 6552 30352 6557 30404
rect 6557 30352 6604 30404
rect 6620 30352 6672 30404
rect 6688 30352 6735 30404
rect 6735 30352 6740 30404
rect 6552 30287 6557 30339
rect 6557 30287 6604 30339
rect 6620 30287 6672 30339
rect 6688 30287 6735 30339
rect 6735 30287 6740 30339
rect 6552 30222 6557 30274
rect 6557 30222 6604 30274
rect 6620 30222 6672 30274
rect 6688 30222 6735 30274
rect 6735 30222 6740 30274
rect 6552 30157 6557 30209
rect 6557 30157 6604 30209
rect 6620 30157 6672 30209
rect 6688 30157 6735 30209
rect 6735 30157 6740 30209
rect 6552 30092 6557 30144
rect 6557 30092 6604 30144
rect 6620 30092 6672 30144
rect 6688 30092 6735 30144
rect 6735 30092 6740 30144
rect 6552 30027 6557 30079
rect 6557 30027 6604 30079
rect 6620 30027 6672 30079
rect 6688 30027 6735 30079
rect 6735 30027 6740 30079
rect 6552 29962 6557 30014
rect 6557 29962 6604 30014
rect 6620 29962 6672 30014
rect 6688 29962 6735 30014
rect 6735 29962 6740 30014
rect 6552 27038 6557 27090
rect 6557 27038 6604 27090
rect 6620 27038 6672 27090
rect 6688 27038 6735 27090
rect 6735 27038 6740 27090
rect 6552 26974 6557 27026
rect 6557 26974 6604 27026
rect 6620 26974 6672 27026
rect 6688 26974 6735 27026
rect 6735 26974 6740 27026
rect 6552 26910 6557 26962
rect 6557 26910 6604 26962
rect 6620 26910 6672 26962
rect 6688 26910 6735 26962
rect 6735 26910 6740 26962
rect 6552 26846 6557 26898
rect 6557 26846 6604 26898
rect 6620 26846 6672 26898
rect 6688 26846 6735 26898
rect 6735 26846 6740 26898
rect 6552 26782 6557 26834
rect 6557 26782 6604 26834
rect 6620 26782 6672 26834
rect 6688 26782 6735 26834
rect 6735 26782 6740 26834
rect 6552 26718 6557 26770
rect 6557 26718 6604 26770
rect 6620 26718 6672 26770
rect 6688 26718 6735 26770
rect 6735 26718 6740 26770
rect 6552 26654 6557 26706
rect 6557 26654 6604 26706
rect 6620 26654 6672 26706
rect 6688 26654 6735 26706
rect 6735 26654 6740 26706
rect 6552 26590 6557 26642
rect 6557 26590 6604 26642
rect 6620 26590 6672 26642
rect 6688 26590 6735 26642
rect 6735 26590 6740 26642
rect 6552 26526 6557 26578
rect 6557 26526 6604 26578
rect 6620 26526 6672 26578
rect 6688 26526 6735 26578
rect 6735 26526 6740 26578
rect 6552 26462 6557 26514
rect 6557 26462 6604 26514
rect 6620 26462 6672 26514
rect 6688 26462 6735 26514
rect 6735 26462 6740 26514
rect 6552 26398 6557 26450
rect 6557 26398 6604 26450
rect 6620 26398 6672 26450
rect 6688 26398 6735 26450
rect 6735 26398 6740 26450
rect 6552 26334 6557 26386
rect 6557 26334 6604 26386
rect 6620 26334 6672 26386
rect 6688 26334 6735 26386
rect 6735 26334 6740 26386
rect 6552 26270 6557 26322
rect 6557 26270 6604 26322
rect 6620 26270 6672 26322
rect 6688 26270 6735 26322
rect 6735 26270 6740 26322
rect 6552 26206 6557 26258
rect 6557 26206 6604 26258
rect 6620 26206 6672 26258
rect 6688 26206 6735 26258
rect 6735 26206 6740 26258
rect 6552 26142 6557 26194
rect 6557 26142 6604 26194
rect 6620 26142 6672 26194
rect 6688 26142 6735 26194
rect 6735 26142 6740 26194
rect 6552 26077 6557 26129
rect 6557 26077 6604 26129
rect 6620 26077 6672 26129
rect 6688 26077 6735 26129
rect 6735 26077 6740 26129
rect 6552 26012 6557 26064
rect 6557 26012 6604 26064
rect 6620 26012 6672 26064
rect 6688 26012 6735 26064
rect 6735 26012 6740 26064
rect 6552 25947 6557 25999
rect 6557 25947 6604 25999
rect 6620 25947 6672 25999
rect 6688 25947 6735 25999
rect 6735 25947 6740 25999
rect 6552 25882 6557 25934
rect 6557 25882 6604 25934
rect 6620 25882 6672 25934
rect 6688 25882 6735 25934
rect 6735 25882 6740 25934
rect 6552 25817 6557 25869
rect 6557 25817 6604 25869
rect 6620 25817 6672 25869
rect 6688 25817 6735 25869
rect 6735 25817 6740 25869
rect 6552 25752 6557 25804
rect 6557 25752 6604 25804
rect 6620 25752 6672 25804
rect 6688 25752 6735 25804
rect 6735 25752 6740 25804
rect 6552 25687 6557 25739
rect 6557 25687 6604 25739
rect 6620 25687 6672 25739
rect 6688 25687 6735 25739
rect 6735 25687 6740 25739
rect 6552 25622 6557 25674
rect 6557 25622 6604 25674
rect 6620 25622 6672 25674
rect 6688 25622 6735 25674
rect 6735 25622 6740 25674
rect 6552 25557 6557 25609
rect 6557 25557 6604 25609
rect 6620 25557 6672 25609
rect 6688 25557 6735 25609
rect 6735 25557 6740 25609
rect 6552 25492 6557 25544
rect 6557 25492 6604 25544
rect 6620 25492 6672 25544
rect 6688 25492 6735 25544
rect 6735 25492 6740 25544
rect 6552 25427 6557 25479
rect 6557 25427 6604 25479
rect 6620 25427 6672 25479
rect 6688 25427 6735 25479
rect 6735 25427 6740 25479
rect 6552 25362 6557 25414
rect 6557 25362 6604 25414
rect 6620 25362 6672 25414
rect 6688 25362 6735 25414
rect 6735 25362 6740 25414
rect 6552 22438 6557 22490
rect 6557 22438 6604 22490
rect 6620 22438 6672 22490
rect 6688 22438 6735 22490
rect 6735 22438 6740 22490
rect 6552 22374 6557 22426
rect 6557 22374 6604 22426
rect 6620 22374 6672 22426
rect 6688 22374 6735 22426
rect 6735 22374 6740 22426
rect 6552 22310 6557 22362
rect 6557 22310 6604 22362
rect 6620 22310 6672 22362
rect 6688 22310 6735 22362
rect 6735 22310 6740 22362
rect 6552 22246 6557 22298
rect 6557 22246 6604 22298
rect 6620 22246 6672 22298
rect 6688 22246 6735 22298
rect 6735 22246 6740 22298
rect 6552 22182 6557 22234
rect 6557 22182 6604 22234
rect 6620 22182 6672 22234
rect 6688 22182 6735 22234
rect 6735 22182 6740 22234
rect 6552 22118 6557 22170
rect 6557 22118 6604 22170
rect 6620 22118 6672 22170
rect 6688 22118 6735 22170
rect 6735 22118 6740 22170
rect 6552 22054 6557 22106
rect 6557 22054 6604 22106
rect 6620 22054 6672 22106
rect 6688 22054 6735 22106
rect 6735 22054 6740 22106
rect 6552 21990 6557 22042
rect 6557 21990 6604 22042
rect 6620 21990 6672 22042
rect 6688 21990 6735 22042
rect 6735 21990 6740 22042
rect 6552 21926 6557 21978
rect 6557 21926 6604 21978
rect 6620 21926 6672 21978
rect 6688 21926 6735 21978
rect 6735 21926 6740 21978
rect 6552 21862 6557 21914
rect 6557 21862 6604 21914
rect 6620 21862 6672 21914
rect 6688 21862 6735 21914
rect 6735 21862 6740 21914
rect 6552 21798 6557 21850
rect 6557 21798 6604 21850
rect 6620 21798 6672 21850
rect 6688 21798 6735 21850
rect 6735 21798 6740 21850
rect 6552 21734 6557 21786
rect 6557 21734 6604 21786
rect 6620 21734 6672 21786
rect 6688 21734 6735 21786
rect 6735 21734 6740 21786
rect 6552 21670 6557 21722
rect 6557 21670 6604 21722
rect 6620 21670 6672 21722
rect 6688 21670 6735 21722
rect 6735 21670 6740 21722
rect 6552 21606 6557 21658
rect 6557 21606 6604 21658
rect 6620 21606 6672 21658
rect 6688 21606 6735 21658
rect 6735 21606 6740 21658
rect 6552 21542 6557 21594
rect 6557 21542 6604 21594
rect 6620 21542 6672 21594
rect 6688 21542 6735 21594
rect 6735 21542 6740 21594
rect 6552 21477 6557 21529
rect 6557 21477 6604 21529
rect 6620 21477 6672 21529
rect 6688 21477 6735 21529
rect 6735 21477 6740 21529
rect 6552 21412 6557 21464
rect 6557 21412 6604 21464
rect 6620 21412 6672 21464
rect 6688 21412 6735 21464
rect 6735 21412 6740 21464
rect 6552 21347 6557 21399
rect 6557 21347 6604 21399
rect 6620 21347 6672 21399
rect 6688 21347 6735 21399
rect 6735 21347 6740 21399
rect 6552 21282 6557 21334
rect 6557 21282 6604 21334
rect 6620 21282 6672 21334
rect 6688 21282 6735 21334
rect 6735 21282 6740 21334
rect 6552 21217 6557 21269
rect 6557 21217 6604 21269
rect 6620 21217 6672 21269
rect 6688 21217 6735 21269
rect 6735 21217 6740 21269
rect 6552 21152 6557 21204
rect 6557 21152 6604 21204
rect 6620 21152 6672 21204
rect 6688 21152 6735 21204
rect 6735 21152 6740 21204
rect 6552 21087 6557 21139
rect 6557 21087 6604 21139
rect 6620 21087 6672 21139
rect 6688 21087 6735 21139
rect 6735 21087 6740 21139
rect 6552 21022 6557 21074
rect 6557 21022 6604 21074
rect 6620 21022 6672 21074
rect 6688 21022 6735 21074
rect 6735 21022 6740 21074
rect 6552 20957 6557 21009
rect 6557 20957 6604 21009
rect 6620 20957 6672 21009
rect 6688 20957 6735 21009
rect 6735 20957 6740 21009
rect 6552 20892 6557 20944
rect 6557 20892 6604 20944
rect 6620 20892 6672 20944
rect 6688 20892 6735 20944
rect 6735 20892 6740 20944
rect 6552 20827 6557 20879
rect 6557 20827 6604 20879
rect 6620 20827 6672 20879
rect 6688 20827 6735 20879
rect 6735 20827 6740 20879
rect 6552 20762 6557 20814
rect 6557 20762 6604 20814
rect 6620 20762 6672 20814
rect 6688 20762 6735 20814
rect 6735 20762 6740 20814
rect 6552 17838 6557 17890
rect 6557 17838 6604 17890
rect 6620 17838 6672 17890
rect 6688 17838 6735 17890
rect 6735 17838 6740 17890
rect 6552 17774 6557 17826
rect 6557 17774 6604 17826
rect 6620 17774 6672 17826
rect 6688 17774 6735 17826
rect 6735 17774 6740 17826
rect 6552 17710 6557 17762
rect 6557 17710 6604 17762
rect 6620 17710 6672 17762
rect 6688 17710 6735 17762
rect 6735 17710 6740 17762
rect 6552 17646 6557 17698
rect 6557 17646 6604 17698
rect 6620 17646 6672 17698
rect 6688 17646 6735 17698
rect 6735 17646 6740 17698
rect 6552 17582 6557 17634
rect 6557 17582 6604 17634
rect 6620 17582 6672 17634
rect 6688 17582 6735 17634
rect 6735 17582 6740 17634
rect 6552 17518 6557 17570
rect 6557 17518 6604 17570
rect 6620 17518 6672 17570
rect 6688 17518 6735 17570
rect 6735 17518 6740 17570
rect 6552 17454 6557 17506
rect 6557 17454 6604 17506
rect 6620 17454 6672 17506
rect 6688 17454 6735 17506
rect 6735 17454 6740 17506
rect 6552 17390 6557 17442
rect 6557 17390 6604 17442
rect 6620 17390 6672 17442
rect 6688 17390 6735 17442
rect 6735 17390 6740 17442
rect 6552 17326 6557 17378
rect 6557 17326 6604 17378
rect 6620 17326 6672 17378
rect 6688 17326 6735 17378
rect 6735 17326 6740 17378
rect 6552 17262 6557 17314
rect 6557 17262 6604 17314
rect 6620 17262 6672 17314
rect 6688 17262 6735 17314
rect 6735 17262 6740 17314
rect 6552 17198 6557 17250
rect 6557 17198 6604 17250
rect 6620 17198 6672 17250
rect 6688 17198 6735 17250
rect 6735 17198 6740 17250
rect 6552 17134 6557 17186
rect 6557 17134 6604 17186
rect 6620 17134 6672 17186
rect 6688 17134 6735 17186
rect 6735 17134 6740 17186
rect 6552 17070 6557 17122
rect 6557 17070 6604 17122
rect 6620 17070 6672 17122
rect 6688 17070 6735 17122
rect 6735 17070 6740 17122
rect 6552 17006 6557 17058
rect 6557 17006 6604 17058
rect 6620 17006 6672 17058
rect 6688 17006 6735 17058
rect 6735 17006 6740 17058
rect 6552 16942 6557 16994
rect 6557 16942 6604 16994
rect 6620 16942 6672 16994
rect 6688 16942 6735 16994
rect 6735 16942 6740 16994
rect 6552 16877 6557 16929
rect 6557 16877 6604 16929
rect 6620 16877 6672 16929
rect 6688 16877 6735 16929
rect 6735 16877 6740 16929
rect 6552 16812 6557 16864
rect 6557 16812 6604 16864
rect 6620 16812 6672 16864
rect 6688 16812 6735 16864
rect 6735 16812 6740 16864
rect 6552 16747 6557 16799
rect 6557 16747 6604 16799
rect 6620 16747 6672 16799
rect 6688 16747 6735 16799
rect 6735 16747 6740 16799
rect 6552 16682 6557 16734
rect 6557 16682 6604 16734
rect 6620 16682 6672 16734
rect 6688 16682 6735 16734
rect 6735 16682 6740 16734
rect 6552 16617 6557 16669
rect 6557 16617 6604 16669
rect 6620 16617 6672 16669
rect 6688 16617 6735 16669
rect 6735 16617 6740 16669
rect 6552 16552 6557 16604
rect 6557 16552 6604 16604
rect 6620 16552 6672 16604
rect 6688 16552 6735 16604
rect 6735 16552 6740 16604
rect 6552 16487 6557 16539
rect 6557 16487 6604 16539
rect 6620 16487 6672 16539
rect 6688 16487 6735 16539
rect 6735 16487 6740 16539
rect 6552 16422 6557 16474
rect 6557 16422 6604 16474
rect 6620 16422 6672 16474
rect 6688 16422 6735 16474
rect 6735 16422 6740 16474
rect 6552 16357 6557 16409
rect 6557 16357 6604 16409
rect 6620 16357 6672 16409
rect 6688 16357 6735 16409
rect 6735 16357 6740 16409
rect 6552 16292 6557 16344
rect 6557 16292 6604 16344
rect 6620 16292 6672 16344
rect 6688 16292 6735 16344
rect 6735 16292 6740 16344
rect 6552 16227 6557 16279
rect 6557 16227 6604 16279
rect 6620 16227 6672 16279
rect 6688 16227 6735 16279
rect 6735 16227 6740 16279
rect 6552 16162 6557 16214
rect 6557 16162 6604 16214
rect 6620 16162 6672 16214
rect 6688 16162 6735 16214
rect 6735 16162 6740 16214
rect 6552 13238 6557 13290
rect 6557 13238 6604 13290
rect 6620 13238 6672 13290
rect 6688 13238 6735 13290
rect 6735 13238 6740 13290
rect 6552 13174 6557 13226
rect 6557 13174 6604 13226
rect 6620 13174 6672 13226
rect 6688 13174 6735 13226
rect 6735 13174 6740 13226
rect 6552 13110 6557 13162
rect 6557 13110 6604 13162
rect 6620 13110 6672 13162
rect 6688 13110 6735 13162
rect 6735 13110 6740 13162
rect 6552 13046 6557 13098
rect 6557 13046 6604 13098
rect 6620 13046 6672 13098
rect 6688 13046 6735 13098
rect 6735 13046 6740 13098
rect 6552 12982 6557 13034
rect 6557 12982 6604 13034
rect 6620 12982 6672 13034
rect 6688 12982 6735 13034
rect 6735 12982 6740 13034
rect 6552 12918 6557 12970
rect 6557 12918 6604 12970
rect 6620 12918 6672 12970
rect 6688 12918 6735 12970
rect 6735 12918 6740 12970
rect 6552 12854 6557 12906
rect 6557 12854 6604 12906
rect 6620 12854 6672 12906
rect 6688 12854 6735 12906
rect 6735 12854 6740 12906
rect 6552 12790 6557 12842
rect 6557 12790 6604 12842
rect 6620 12790 6672 12842
rect 6688 12790 6735 12842
rect 6735 12790 6740 12842
rect 6552 12726 6557 12778
rect 6557 12726 6604 12778
rect 6620 12726 6672 12778
rect 6688 12726 6735 12778
rect 6735 12726 6740 12778
rect 6552 12662 6557 12714
rect 6557 12662 6604 12714
rect 6620 12662 6672 12714
rect 6688 12662 6735 12714
rect 6735 12662 6740 12714
rect 6552 12598 6557 12650
rect 6557 12598 6604 12650
rect 6620 12598 6672 12650
rect 6688 12598 6735 12650
rect 6735 12598 6740 12650
rect 6552 12534 6557 12586
rect 6557 12534 6604 12586
rect 6620 12534 6672 12586
rect 6688 12534 6735 12586
rect 6735 12534 6740 12586
rect 6552 12470 6557 12522
rect 6557 12470 6604 12522
rect 6620 12470 6672 12522
rect 6688 12470 6735 12522
rect 6735 12470 6740 12522
rect 6552 12406 6557 12458
rect 6557 12406 6604 12458
rect 6620 12406 6672 12458
rect 6688 12406 6735 12458
rect 6735 12406 6740 12458
rect 6552 12342 6557 12394
rect 6557 12342 6604 12394
rect 6620 12342 6672 12394
rect 6688 12342 6735 12394
rect 6735 12342 6740 12394
rect 6552 12277 6557 12329
rect 6557 12277 6604 12329
rect 6620 12277 6672 12329
rect 6688 12277 6735 12329
rect 6735 12277 6740 12329
rect 6552 12212 6557 12264
rect 6557 12212 6604 12264
rect 6620 12212 6672 12264
rect 6688 12212 6735 12264
rect 6735 12212 6740 12264
rect 6552 12147 6557 12199
rect 6557 12147 6604 12199
rect 6620 12147 6672 12199
rect 6688 12147 6735 12199
rect 6735 12147 6740 12199
rect 6552 12082 6557 12134
rect 6557 12082 6604 12134
rect 6620 12082 6672 12134
rect 6688 12082 6735 12134
rect 6735 12082 6740 12134
rect 6552 12017 6557 12069
rect 6557 12017 6604 12069
rect 6620 12017 6672 12069
rect 6688 12017 6735 12069
rect 6735 12017 6740 12069
rect 6552 11952 6557 12004
rect 6557 11952 6604 12004
rect 6620 11952 6672 12004
rect 6688 11952 6735 12004
rect 6735 11952 6740 12004
rect 6552 11887 6557 11939
rect 6557 11887 6604 11939
rect 6620 11887 6672 11939
rect 6688 11887 6735 11939
rect 6735 11887 6740 11939
rect 6552 11822 6557 11874
rect 6557 11822 6604 11874
rect 6620 11822 6672 11874
rect 6688 11822 6735 11874
rect 6735 11822 6740 11874
rect 6552 11757 6557 11809
rect 6557 11757 6604 11809
rect 6620 11757 6672 11809
rect 6688 11757 6735 11809
rect 6735 11757 6740 11809
rect 6552 11692 6557 11744
rect 6557 11692 6604 11744
rect 6620 11692 6672 11744
rect 6688 11692 6735 11744
rect 6735 11692 6740 11744
rect 6552 11627 6557 11679
rect 6557 11627 6604 11679
rect 6620 11627 6672 11679
rect 6688 11627 6735 11679
rect 6735 11627 6740 11679
rect 6552 11562 6557 11614
rect 6557 11562 6604 11614
rect 6620 11562 6672 11614
rect 6688 11562 6735 11614
rect 6735 11562 6740 11614
rect 7041 37945 7093 37997
rect 7119 37945 7171 37997
rect 7041 37877 7093 37929
rect 7119 37877 7171 37929
rect 7041 37809 7093 37861
rect 7119 37809 7171 37861
rect 7041 37741 7093 37793
rect 7119 37741 7171 37793
rect 7041 37673 7093 37725
rect 7119 37673 7171 37725
rect 7041 37605 7093 37657
rect 7119 37605 7171 37657
rect 7041 37537 7093 37589
rect 7119 37537 7171 37589
rect 7041 37469 7093 37521
rect 7119 37469 7171 37521
rect 7041 37401 7093 37453
rect 7119 37401 7171 37453
rect 7041 37333 7093 37385
rect 7119 37333 7171 37385
rect 7041 37266 7093 37318
rect 7119 37266 7171 37318
rect 7041 37199 7093 37251
rect 7119 37199 7171 37251
rect 7041 37132 7093 37184
rect 7119 37132 7171 37184
rect 7041 37065 7093 37117
rect 7119 37065 7171 37117
rect 7041 34173 7093 34225
rect 7119 34173 7171 34225
rect 7041 34109 7093 34161
rect 7119 34109 7171 34161
rect 7041 34045 7093 34097
rect 7119 34045 7171 34097
rect 7041 33981 7093 34033
rect 7119 33981 7171 34033
rect 7041 33917 7093 33969
rect 7119 33917 7171 33969
rect 7041 33853 7093 33905
rect 7119 33853 7171 33905
rect 7041 33789 7093 33841
rect 7119 33789 7171 33841
rect 7041 33725 7093 33777
rect 7119 33725 7171 33777
rect 7041 33661 7093 33713
rect 7119 33661 7171 33713
rect 7041 33597 7093 33649
rect 7119 33597 7171 33649
rect 7041 33533 7093 33585
rect 7119 33533 7171 33585
rect 7041 33469 7093 33521
rect 7119 33469 7171 33521
rect 7041 33405 7093 33457
rect 7119 33405 7171 33457
rect 7041 33341 7093 33393
rect 7119 33341 7171 33393
rect 7041 33277 7093 33329
rect 7119 33277 7171 33329
rect 7041 33212 7093 33264
rect 7119 33212 7171 33264
rect 7041 33147 7093 33199
rect 7119 33147 7171 33199
rect 7041 33082 7093 33134
rect 7119 33082 7171 33134
rect 7041 33017 7093 33069
rect 7119 33017 7171 33069
rect 7041 32952 7093 33004
rect 7119 32952 7171 33004
rect 7041 32887 7093 32939
rect 7119 32887 7171 32939
rect 7041 32822 7093 32874
rect 7119 32822 7171 32874
rect 7041 32757 7093 32809
rect 7119 32757 7171 32809
rect 7041 32692 7093 32744
rect 7119 32692 7171 32744
rect 7041 32627 7093 32679
rect 7119 32627 7171 32679
rect 7041 32562 7093 32614
rect 7119 32562 7171 32614
rect 7041 32497 7093 32549
rect 7119 32497 7171 32549
rect 7041 29573 7093 29625
rect 7119 29573 7171 29625
rect 7041 29509 7093 29561
rect 7119 29509 7171 29561
rect 7041 29445 7093 29497
rect 7119 29445 7171 29497
rect 7041 29381 7093 29433
rect 7119 29381 7171 29433
rect 7041 29317 7093 29369
rect 7119 29317 7171 29369
rect 7041 29253 7093 29305
rect 7119 29253 7171 29305
rect 7041 29189 7093 29241
rect 7119 29189 7171 29241
rect 7041 29125 7093 29177
rect 7119 29125 7171 29177
rect 7041 29061 7093 29113
rect 7119 29061 7171 29113
rect 7041 28997 7093 29049
rect 7119 28997 7171 29049
rect 7041 28933 7093 28985
rect 7119 28933 7171 28985
rect 7041 28869 7093 28921
rect 7119 28869 7171 28921
rect 7041 28805 7093 28857
rect 7119 28805 7171 28857
rect 7041 28741 7093 28793
rect 7119 28741 7171 28793
rect 7041 28677 7093 28729
rect 7119 28677 7171 28729
rect 7041 28612 7093 28664
rect 7119 28612 7171 28664
rect 7041 28547 7093 28599
rect 7119 28547 7171 28599
rect 7041 28482 7093 28534
rect 7119 28482 7171 28534
rect 7041 28417 7093 28469
rect 7119 28417 7171 28469
rect 7041 28352 7093 28404
rect 7119 28352 7171 28404
rect 7041 28287 7093 28339
rect 7119 28287 7171 28339
rect 7041 28222 7093 28274
rect 7119 28222 7171 28274
rect 7041 28157 7093 28209
rect 7119 28157 7171 28209
rect 7041 28092 7093 28144
rect 7119 28092 7171 28144
rect 7041 28027 7093 28079
rect 7119 28027 7171 28079
rect 7041 27962 7093 28014
rect 7119 27962 7171 28014
rect 7041 27897 7093 27949
rect 7119 27897 7171 27949
rect 7041 24973 7093 25025
rect 7119 24973 7171 25025
rect 7041 24909 7093 24961
rect 7119 24909 7171 24961
rect 7041 24845 7093 24897
rect 7119 24845 7171 24897
rect 7041 24781 7093 24833
rect 7119 24781 7171 24833
rect 7041 24717 7093 24769
rect 7119 24717 7171 24769
rect 7041 24653 7093 24705
rect 7119 24653 7171 24705
rect 7041 24589 7093 24641
rect 7119 24589 7171 24641
rect 7041 24525 7093 24577
rect 7119 24525 7171 24577
rect 7041 24461 7093 24513
rect 7119 24461 7171 24513
rect 7041 24397 7093 24449
rect 7119 24397 7171 24449
rect 7041 24333 7093 24385
rect 7119 24333 7171 24385
rect 7041 24269 7093 24321
rect 7119 24269 7171 24321
rect 7041 24205 7093 24257
rect 7119 24205 7171 24257
rect 7041 24141 7093 24193
rect 7119 24141 7171 24193
rect 7041 24077 7093 24129
rect 7119 24077 7171 24129
rect 7041 24012 7093 24064
rect 7119 24012 7171 24064
rect 7041 23947 7093 23999
rect 7119 23947 7171 23999
rect 7041 23882 7093 23934
rect 7119 23882 7171 23934
rect 7041 23817 7093 23869
rect 7119 23817 7171 23869
rect 7041 23752 7093 23804
rect 7119 23752 7171 23804
rect 7041 23687 7093 23739
rect 7119 23687 7171 23739
rect 7041 23622 7093 23674
rect 7119 23622 7171 23674
rect 7041 23557 7093 23609
rect 7119 23557 7171 23609
rect 7041 23492 7093 23544
rect 7119 23492 7171 23544
rect 7041 23427 7093 23479
rect 7119 23427 7171 23479
rect 7041 23362 7093 23414
rect 7119 23362 7171 23414
rect 7041 23297 7093 23349
rect 7119 23297 7171 23349
rect 7041 20373 7093 20425
rect 7119 20373 7171 20425
rect 7041 20309 7093 20361
rect 7119 20309 7171 20361
rect 7041 20245 7093 20297
rect 7119 20245 7171 20297
rect 7041 20181 7093 20233
rect 7119 20181 7171 20233
rect 7041 20117 7093 20169
rect 7119 20117 7171 20169
rect 7041 20053 7093 20105
rect 7119 20053 7171 20105
rect 7041 19989 7093 20041
rect 7119 19989 7171 20041
rect 7041 19925 7093 19977
rect 7119 19925 7171 19977
rect 7041 19861 7093 19913
rect 7119 19861 7171 19913
rect 7041 19797 7093 19849
rect 7119 19797 7171 19849
rect 7041 19733 7093 19785
rect 7119 19733 7171 19785
rect 7041 19669 7093 19721
rect 7119 19669 7171 19721
rect 7041 19605 7093 19657
rect 7119 19605 7171 19657
rect 7041 19541 7093 19593
rect 7119 19541 7171 19593
rect 7041 19477 7093 19529
rect 7119 19477 7171 19529
rect 7041 19412 7093 19464
rect 7119 19412 7171 19464
rect 7041 19347 7093 19399
rect 7119 19347 7171 19399
rect 7041 19282 7093 19334
rect 7119 19282 7171 19334
rect 7041 19217 7093 19269
rect 7119 19217 7171 19269
rect 7041 19152 7093 19204
rect 7119 19152 7171 19204
rect 7041 19087 7093 19139
rect 7119 19087 7171 19139
rect 7041 19022 7093 19074
rect 7119 19022 7171 19074
rect 7041 18957 7093 19009
rect 7119 18957 7171 19009
rect 7041 18892 7093 18944
rect 7119 18892 7171 18944
rect 7041 18827 7093 18879
rect 7119 18827 7171 18879
rect 7041 18762 7093 18814
rect 7119 18762 7171 18814
rect 7041 18697 7093 18749
rect 7119 18697 7171 18749
rect 7041 15773 7093 15825
rect 7119 15773 7171 15825
rect 7041 15709 7093 15761
rect 7119 15709 7171 15761
rect 7041 15645 7093 15697
rect 7119 15645 7171 15697
rect 7041 15581 7093 15633
rect 7119 15581 7171 15633
rect 7041 15517 7093 15569
rect 7119 15517 7171 15569
rect 7041 15453 7093 15505
rect 7119 15453 7171 15505
rect 7041 15389 7093 15441
rect 7119 15389 7171 15441
rect 7041 15325 7093 15377
rect 7119 15325 7171 15377
rect 7041 15261 7093 15313
rect 7119 15261 7171 15313
rect 7041 15197 7093 15249
rect 7119 15197 7171 15249
rect 7041 15133 7093 15185
rect 7119 15133 7171 15185
rect 7041 15069 7093 15121
rect 7119 15069 7171 15121
rect 7041 15005 7093 15057
rect 7119 15005 7171 15057
rect 7041 14941 7093 14993
rect 7119 14941 7171 14993
rect 7041 14877 7093 14929
rect 7119 14877 7171 14929
rect 7041 14812 7093 14864
rect 7119 14812 7171 14864
rect 7041 14747 7093 14799
rect 7119 14747 7171 14799
rect 7041 14682 7093 14734
rect 7119 14682 7171 14734
rect 7041 14617 7093 14669
rect 7119 14617 7171 14669
rect 7041 14552 7093 14604
rect 7119 14552 7171 14604
rect 7041 14487 7093 14539
rect 7119 14487 7171 14539
rect 7041 14422 7093 14474
rect 7119 14422 7171 14474
rect 7041 14357 7093 14409
rect 7119 14357 7171 14409
rect 7041 14292 7093 14344
rect 7119 14292 7171 14344
rect 7041 14227 7093 14279
rect 7119 14227 7171 14279
rect 7041 14162 7093 14214
rect 7119 14162 7171 14214
rect 7041 14097 7093 14149
rect 7119 14097 7171 14149
rect 7041 11173 7093 11225
rect 7119 11173 7171 11225
rect 7041 11109 7093 11161
rect 7119 11109 7171 11161
rect 7041 11045 7093 11097
rect 7119 11045 7171 11097
rect 7041 10981 7093 11033
rect 7119 10981 7171 11033
rect 7041 10917 7093 10969
rect 7119 10917 7171 10969
rect 7041 10853 7093 10905
rect 7119 10853 7171 10905
rect 7041 10789 7093 10841
rect 7119 10789 7171 10841
rect 7041 10725 7093 10777
rect 7119 10725 7171 10777
rect 7041 10661 7093 10713
rect 7119 10661 7171 10713
rect 7041 10597 7093 10649
rect 7119 10597 7171 10649
rect 7041 10533 7093 10585
rect 7119 10533 7171 10585
rect 7041 10469 7093 10521
rect 7119 10469 7171 10521
rect 7041 10405 7093 10457
rect 7119 10405 7171 10457
rect 7041 10341 7093 10393
rect 7119 10341 7171 10393
rect 7041 10277 7093 10329
rect 7119 10277 7171 10329
rect 7041 10212 7093 10264
rect 7119 10212 7171 10264
rect 7041 10147 7093 10199
rect 7119 10147 7171 10199
rect 7041 10082 7093 10134
rect 7119 10082 7171 10134
rect 7041 10017 7093 10069
rect 7119 10017 7171 10069
rect 7041 9952 7093 10004
rect 7119 9952 7171 10004
rect 7041 9887 7093 9939
rect 7119 9887 7171 9939
rect 7041 9822 7093 9874
rect 7119 9822 7171 9874
rect 7041 9757 7093 9809
rect 7119 9757 7171 9809
rect 7041 9692 7093 9744
rect 7119 9692 7171 9744
rect 7041 9627 7093 9679
rect 7119 9627 7171 9679
rect 7041 9562 7093 9614
rect 7119 9562 7171 9614
rect 7041 9497 7093 9549
rect 7119 9497 7171 9549
rect 7472 36238 7477 36290
rect 7477 36238 7524 36290
rect 7540 36238 7592 36290
rect 7608 36238 7655 36290
rect 7655 36238 7660 36290
rect 7472 36174 7477 36226
rect 7477 36174 7524 36226
rect 7540 36174 7592 36226
rect 7608 36174 7655 36226
rect 7655 36174 7660 36226
rect 7472 36110 7477 36162
rect 7477 36110 7524 36162
rect 7540 36110 7592 36162
rect 7608 36110 7655 36162
rect 7655 36110 7660 36162
rect 7472 36046 7477 36098
rect 7477 36046 7524 36098
rect 7540 36046 7592 36098
rect 7608 36046 7655 36098
rect 7655 36046 7660 36098
rect 7472 35982 7477 36034
rect 7477 35982 7524 36034
rect 7540 35982 7592 36034
rect 7608 35982 7655 36034
rect 7655 35982 7660 36034
rect 7472 35918 7477 35970
rect 7477 35918 7524 35970
rect 7540 35918 7592 35970
rect 7608 35918 7655 35970
rect 7655 35918 7660 35970
rect 7472 35854 7477 35906
rect 7477 35854 7524 35906
rect 7540 35854 7592 35906
rect 7608 35854 7655 35906
rect 7655 35854 7660 35906
rect 7472 35790 7477 35842
rect 7477 35790 7524 35842
rect 7540 35790 7592 35842
rect 7608 35790 7655 35842
rect 7655 35790 7660 35842
rect 7472 35726 7477 35778
rect 7477 35726 7524 35778
rect 7540 35726 7592 35778
rect 7608 35726 7655 35778
rect 7655 35726 7660 35778
rect 7472 35662 7477 35714
rect 7477 35662 7524 35714
rect 7540 35662 7592 35714
rect 7608 35662 7655 35714
rect 7655 35662 7660 35714
rect 7472 35598 7477 35650
rect 7477 35598 7524 35650
rect 7540 35598 7592 35650
rect 7608 35598 7655 35650
rect 7655 35598 7660 35650
rect 7472 35534 7477 35586
rect 7477 35534 7524 35586
rect 7540 35534 7592 35586
rect 7608 35534 7655 35586
rect 7655 35534 7660 35586
rect 7472 35470 7477 35522
rect 7477 35470 7524 35522
rect 7540 35470 7592 35522
rect 7608 35470 7655 35522
rect 7655 35470 7660 35522
rect 7472 35406 7477 35458
rect 7477 35406 7524 35458
rect 7540 35406 7592 35458
rect 7608 35406 7655 35458
rect 7655 35406 7660 35458
rect 7472 35342 7477 35394
rect 7477 35342 7524 35394
rect 7540 35342 7592 35394
rect 7608 35342 7655 35394
rect 7655 35342 7660 35394
rect 7472 35277 7477 35329
rect 7477 35277 7524 35329
rect 7540 35277 7592 35329
rect 7608 35277 7655 35329
rect 7655 35277 7660 35329
rect 7472 35212 7477 35264
rect 7477 35212 7524 35264
rect 7540 35212 7592 35264
rect 7608 35212 7655 35264
rect 7655 35212 7660 35264
rect 7472 35147 7477 35199
rect 7477 35147 7524 35199
rect 7540 35147 7592 35199
rect 7608 35147 7655 35199
rect 7655 35147 7660 35199
rect 7472 35082 7477 35134
rect 7477 35082 7524 35134
rect 7540 35082 7592 35134
rect 7608 35082 7655 35134
rect 7655 35082 7660 35134
rect 7472 35017 7477 35069
rect 7477 35017 7524 35069
rect 7540 35017 7592 35069
rect 7608 35017 7655 35069
rect 7655 35017 7660 35069
rect 7472 34952 7477 35004
rect 7477 34952 7524 35004
rect 7540 34952 7592 35004
rect 7608 34952 7655 35004
rect 7655 34952 7660 35004
rect 7472 34887 7477 34939
rect 7477 34887 7524 34939
rect 7540 34887 7592 34939
rect 7608 34887 7655 34939
rect 7655 34887 7660 34939
rect 7472 34822 7477 34874
rect 7477 34822 7524 34874
rect 7540 34822 7592 34874
rect 7608 34822 7655 34874
rect 7655 34822 7660 34874
rect 7472 34757 7477 34809
rect 7477 34757 7524 34809
rect 7540 34757 7592 34809
rect 7608 34757 7655 34809
rect 7655 34757 7660 34809
rect 7472 34692 7477 34744
rect 7477 34692 7524 34744
rect 7540 34692 7592 34744
rect 7608 34692 7655 34744
rect 7655 34692 7660 34744
rect 7472 34627 7477 34679
rect 7477 34627 7524 34679
rect 7540 34627 7592 34679
rect 7608 34627 7655 34679
rect 7655 34627 7660 34679
rect 7472 34562 7477 34614
rect 7477 34562 7524 34614
rect 7540 34562 7592 34614
rect 7608 34562 7655 34614
rect 7655 34562 7660 34614
rect 7472 31638 7477 31690
rect 7477 31638 7524 31690
rect 7540 31638 7592 31690
rect 7608 31638 7655 31690
rect 7655 31638 7660 31690
rect 7472 31574 7477 31626
rect 7477 31574 7524 31626
rect 7540 31574 7592 31626
rect 7608 31574 7655 31626
rect 7655 31574 7660 31626
rect 7472 31510 7477 31562
rect 7477 31510 7524 31562
rect 7540 31510 7592 31562
rect 7608 31510 7655 31562
rect 7655 31510 7660 31562
rect 7472 31446 7477 31498
rect 7477 31446 7524 31498
rect 7540 31446 7592 31498
rect 7608 31446 7655 31498
rect 7655 31446 7660 31498
rect 7472 31382 7477 31434
rect 7477 31382 7524 31434
rect 7540 31382 7592 31434
rect 7608 31382 7655 31434
rect 7655 31382 7660 31434
rect 7472 31318 7477 31370
rect 7477 31318 7524 31370
rect 7540 31318 7592 31370
rect 7608 31318 7655 31370
rect 7655 31318 7660 31370
rect 7472 31254 7477 31306
rect 7477 31254 7524 31306
rect 7540 31254 7592 31306
rect 7608 31254 7655 31306
rect 7655 31254 7660 31306
rect 7472 31190 7477 31242
rect 7477 31190 7524 31242
rect 7540 31190 7592 31242
rect 7608 31190 7655 31242
rect 7655 31190 7660 31242
rect 7472 31126 7477 31178
rect 7477 31126 7524 31178
rect 7540 31126 7592 31178
rect 7608 31126 7655 31178
rect 7655 31126 7660 31178
rect 7472 31062 7477 31114
rect 7477 31062 7524 31114
rect 7540 31062 7592 31114
rect 7608 31062 7655 31114
rect 7655 31062 7660 31114
rect 7472 30998 7477 31050
rect 7477 30998 7524 31050
rect 7540 30998 7592 31050
rect 7608 30998 7655 31050
rect 7655 30998 7660 31050
rect 7472 30934 7477 30986
rect 7477 30934 7524 30986
rect 7540 30934 7592 30986
rect 7608 30934 7655 30986
rect 7655 30934 7660 30986
rect 7472 30870 7477 30922
rect 7477 30870 7524 30922
rect 7540 30870 7592 30922
rect 7608 30870 7655 30922
rect 7655 30870 7660 30922
rect 7472 30806 7477 30858
rect 7477 30806 7524 30858
rect 7540 30806 7592 30858
rect 7608 30806 7655 30858
rect 7655 30806 7660 30858
rect 7472 30742 7477 30794
rect 7477 30742 7524 30794
rect 7540 30742 7592 30794
rect 7608 30742 7655 30794
rect 7655 30742 7660 30794
rect 7472 30677 7477 30729
rect 7477 30677 7524 30729
rect 7540 30677 7592 30729
rect 7608 30677 7655 30729
rect 7655 30677 7660 30729
rect 7472 30612 7477 30664
rect 7477 30612 7524 30664
rect 7540 30612 7592 30664
rect 7608 30612 7655 30664
rect 7655 30612 7660 30664
rect 7472 30547 7477 30599
rect 7477 30547 7524 30599
rect 7540 30547 7592 30599
rect 7608 30547 7655 30599
rect 7655 30547 7660 30599
rect 7472 30482 7477 30534
rect 7477 30482 7524 30534
rect 7540 30482 7592 30534
rect 7608 30482 7655 30534
rect 7655 30482 7660 30534
rect 7472 30417 7477 30469
rect 7477 30417 7524 30469
rect 7540 30417 7592 30469
rect 7608 30417 7655 30469
rect 7655 30417 7660 30469
rect 7472 30352 7477 30404
rect 7477 30352 7524 30404
rect 7540 30352 7592 30404
rect 7608 30352 7655 30404
rect 7655 30352 7660 30404
rect 7472 30287 7477 30339
rect 7477 30287 7524 30339
rect 7540 30287 7592 30339
rect 7608 30287 7655 30339
rect 7655 30287 7660 30339
rect 7472 30222 7477 30274
rect 7477 30222 7524 30274
rect 7540 30222 7592 30274
rect 7608 30222 7655 30274
rect 7655 30222 7660 30274
rect 7472 30157 7477 30209
rect 7477 30157 7524 30209
rect 7540 30157 7592 30209
rect 7608 30157 7655 30209
rect 7655 30157 7660 30209
rect 7472 30092 7477 30144
rect 7477 30092 7524 30144
rect 7540 30092 7592 30144
rect 7608 30092 7655 30144
rect 7655 30092 7660 30144
rect 7472 30027 7477 30079
rect 7477 30027 7524 30079
rect 7540 30027 7592 30079
rect 7608 30027 7655 30079
rect 7655 30027 7660 30079
rect 7472 29962 7477 30014
rect 7477 29962 7524 30014
rect 7540 29962 7592 30014
rect 7608 29962 7655 30014
rect 7655 29962 7660 30014
rect 7472 27038 7477 27090
rect 7477 27038 7524 27090
rect 7540 27038 7592 27090
rect 7608 27038 7655 27090
rect 7655 27038 7660 27090
rect 7472 26974 7477 27026
rect 7477 26974 7524 27026
rect 7540 26974 7592 27026
rect 7608 26974 7655 27026
rect 7655 26974 7660 27026
rect 7472 26910 7477 26962
rect 7477 26910 7524 26962
rect 7540 26910 7592 26962
rect 7608 26910 7655 26962
rect 7655 26910 7660 26962
rect 7472 26846 7477 26898
rect 7477 26846 7524 26898
rect 7540 26846 7592 26898
rect 7608 26846 7655 26898
rect 7655 26846 7660 26898
rect 7472 26782 7477 26834
rect 7477 26782 7524 26834
rect 7540 26782 7592 26834
rect 7608 26782 7655 26834
rect 7655 26782 7660 26834
rect 7472 26718 7477 26770
rect 7477 26718 7524 26770
rect 7540 26718 7592 26770
rect 7608 26718 7655 26770
rect 7655 26718 7660 26770
rect 7472 26654 7477 26706
rect 7477 26654 7524 26706
rect 7540 26654 7592 26706
rect 7608 26654 7655 26706
rect 7655 26654 7660 26706
rect 7472 26590 7477 26642
rect 7477 26590 7524 26642
rect 7540 26590 7592 26642
rect 7608 26590 7655 26642
rect 7655 26590 7660 26642
rect 7472 26526 7477 26578
rect 7477 26526 7524 26578
rect 7540 26526 7592 26578
rect 7608 26526 7655 26578
rect 7655 26526 7660 26578
rect 7472 26462 7477 26514
rect 7477 26462 7524 26514
rect 7540 26462 7592 26514
rect 7608 26462 7655 26514
rect 7655 26462 7660 26514
rect 7472 26398 7477 26450
rect 7477 26398 7524 26450
rect 7540 26398 7592 26450
rect 7608 26398 7655 26450
rect 7655 26398 7660 26450
rect 7472 26334 7477 26386
rect 7477 26334 7524 26386
rect 7540 26334 7592 26386
rect 7608 26334 7655 26386
rect 7655 26334 7660 26386
rect 7472 26270 7477 26322
rect 7477 26270 7524 26322
rect 7540 26270 7592 26322
rect 7608 26270 7655 26322
rect 7655 26270 7660 26322
rect 7472 26206 7477 26258
rect 7477 26206 7524 26258
rect 7540 26206 7592 26258
rect 7608 26206 7655 26258
rect 7655 26206 7660 26258
rect 7472 26142 7477 26194
rect 7477 26142 7524 26194
rect 7540 26142 7592 26194
rect 7608 26142 7655 26194
rect 7655 26142 7660 26194
rect 7472 26077 7477 26129
rect 7477 26077 7524 26129
rect 7540 26077 7592 26129
rect 7608 26077 7655 26129
rect 7655 26077 7660 26129
rect 7472 26012 7477 26064
rect 7477 26012 7524 26064
rect 7540 26012 7592 26064
rect 7608 26012 7655 26064
rect 7655 26012 7660 26064
rect 7472 25947 7477 25999
rect 7477 25947 7524 25999
rect 7540 25947 7592 25999
rect 7608 25947 7655 25999
rect 7655 25947 7660 25999
rect 7472 25882 7477 25934
rect 7477 25882 7524 25934
rect 7540 25882 7592 25934
rect 7608 25882 7655 25934
rect 7655 25882 7660 25934
rect 7472 25817 7477 25869
rect 7477 25817 7524 25869
rect 7540 25817 7592 25869
rect 7608 25817 7655 25869
rect 7655 25817 7660 25869
rect 7472 25752 7477 25804
rect 7477 25752 7524 25804
rect 7540 25752 7592 25804
rect 7608 25752 7655 25804
rect 7655 25752 7660 25804
rect 7472 25687 7477 25739
rect 7477 25687 7524 25739
rect 7540 25687 7592 25739
rect 7608 25687 7655 25739
rect 7655 25687 7660 25739
rect 7472 25622 7477 25674
rect 7477 25622 7524 25674
rect 7540 25622 7592 25674
rect 7608 25622 7655 25674
rect 7655 25622 7660 25674
rect 7472 25557 7477 25609
rect 7477 25557 7524 25609
rect 7540 25557 7592 25609
rect 7608 25557 7655 25609
rect 7655 25557 7660 25609
rect 7472 25492 7477 25544
rect 7477 25492 7524 25544
rect 7540 25492 7592 25544
rect 7608 25492 7655 25544
rect 7655 25492 7660 25544
rect 7472 25427 7477 25479
rect 7477 25427 7524 25479
rect 7540 25427 7592 25479
rect 7608 25427 7655 25479
rect 7655 25427 7660 25479
rect 7472 25362 7477 25414
rect 7477 25362 7524 25414
rect 7540 25362 7592 25414
rect 7608 25362 7655 25414
rect 7655 25362 7660 25414
rect 7472 22438 7477 22490
rect 7477 22438 7524 22490
rect 7540 22438 7592 22490
rect 7608 22438 7655 22490
rect 7655 22438 7660 22490
rect 7472 22374 7477 22426
rect 7477 22374 7524 22426
rect 7540 22374 7592 22426
rect 7608 22374 7655 22426
rect 7655 22374 7660 22426
rect 7472 22310 7477 22362
rect 7477 22310 7524 22362
rect 7540 22310 7592 22362
rect 7608 22310 7655 22362
rect 7655 22310 7660 22362
rect 7472 22246 7477 22298
rect 7477 22246 7524 22298
rect 7540 22246 7592 22298
rect 7608 22246 7655 22298
rect 7655 22246 7660 22298
rect 7472 22182 7477 22234
rect 7477 22182 7524 22234
rect 7540 22182 7592 22234
rect 7608 22182 7655 22234
rect 7655 22182 7660 22234
rect 7472 22118 7477 22170
rect 7477 22118 7524 22170
rect 7540 22118 7592 22170
rect 7608 22118 7655 22170
rect 7655 22118 7660 22170
rect 7472 22054 7477 22106
rect 7477 22054 7524 22106
rect 7540 22054 7592 22106
rect 7608 22054 7655 22106
rect 7655 22054 7660 22106
rect 7472 21990 7477 22042
rect 7477 21990 7524 22042
rect 7540 21990 7592 22042
rect 7608 21990 7655 22042
rect 7655 21990 7660 22042
rect 7472 21926 7477 21978
rect 7477 21926 7524 21978
rect 7540 21926 7592 21978
rect 7608 21926 7655 21978
rect 7655 21926 7660 21978
rect 7472 21862 7477 21914
rect 7477 21862 7524 21914
rect 7540 21862 7592 21914
rect 7608 21862 7655 21914
rect 7655 21862 7660 21914
rect 7472 21798 7477 21850
rect 7477 21798 7524 21850
rect 7540 21798 7592 21850
rect 7608 21798 7655 21850
rect 7655 21798 7660 21850
rect 7472 21734 7477 21786
rect 7477 21734 7524 21786
rect 7540 21734 7592 21786
rect 7608 21734 7655 21786
rect 7655 21734 7660 21786
rect 7472 21670 7477 21722
rect 7477 21670 7524 21722
rect 7540 21670 7592 21722
rect 7608 21670 7655 21722
rect 7655 21670 7660 21722
rect 7472 21606 7477 21658
rect 7477 21606 7524 21658
rect 7540 21606 7592 21658
rect 7608 21606 7655 21658
rect 7655 21606 7660 21658
rect 7472 21542 7477 21594
rect 7477 21542 7524 21594
rect 7540 21542 7592 21594
rect 7608 21542 7655 21594
rect 7655 21542 7660 21594
rect 7472 21477 7477 21529
rect 7477 21477 7524 21529
rect 7540 21477 7592 21529
rect 7608 21477 7655 21529
rect 7655 21477 7660 21529
rect 7472 21412 7477 21464
rect 7477 21412 7524 21464
rect 7540 21412 7592 21464
rect 7608 21412 7655 21464
rect 7655 21412 7660 21464
rect 7472 21347 7477 21399
rect 7477 21347 7524 21399
rect 7540 21347 7592 21399
rect 7608 21347 7655 21399
rect 7655 21347 7660 21399
rect 7472 21282 7477 21334
rect 7477 21282 7524 21334
rect 7540 21282 7592 21334
rect 7608 21282 7655 21334
rect 7655 21282 7660 21334
rect 7472 21217 7477 21269
rect 7477 21217 7524 21269
rect 7540 21217 7592 21269
rect 7608 21217 7655 21269
rect 7655 21217 7660 21269
rect 7472 21152 7477 21204
rect 7477 21152 7524 21204
rect 7540 21152 7592 21204
rect 7608 21152 7655 21204
rect 7655 21152 7660 21204
rect 7472 21087 7477 21139
rect 7477 21087 7524 21139
rect 7540 21087 7592 21139
rect 7608 21087 7655 21139
rect 7655 21087 7660 21139
rect 7472 21022 7477 21074
rect 7477 21022 7524 21074
rect 7540 21022 7592 21074
rect 7608 21022 7655 21074
rect 7655 21022 7660 21074
rect 7472 20957 7477 21009
rect 7477 20957 7524 21009
rect 7540 20957 7592 21009
rect 7608 20957 7655 21009
rect 7655 20957 7660 21009
rect 7472 20892 7477 20944
rect 7477 20892 7524 20944
rect 7540 20892 7592 20944
rect 7608 20892 7655 20944
rect 7655 20892 7660 20944
rect 7472 20827 7477 20879
rect 7477 20827 7524 20879
rect 7540 20827 7592 20879
rect 7608 20827 7655 20879
rect 7655 20827 7660 20879
rect 7472 20762 7477 20814
rect 7477 20762 7524 20814
rect 7540 20762 7592 20814
rect 7608 20762 7655 20814
rect 7655 20762 7660 20814
rect 7472 17838 7477 17890
rect 7477 17838 7524 17890
rect 7540 17838 7592 17890
rect 7608 17838 7655 17890
rect 7655 17838 7660 17890
rect 7472 17774 7477 17826
rect 7477 17774 7524 17826
rect 7540 17774 7592 17826
rect 7608 17774 7655 17826
rect 7655 17774 7660 17826
rect 7472 17710 7477 17762
rect 7477 17710 7524 17762
rect 7540 17710 7592 17762
rect 7608 17710 7655 17762
rect 7655 17710 7660 17762
rect 7472 17646 7477 17698
rect 7477 17646 7524 17698
rect 7540 17646 7592 17698
rect 7608 17646 7655 17698
rect 7655 17646 7660 17698
rect 7472 17582 7477 17634
rect 7477 17582 7524 17634
rect 7540 17582 7592 17634
rect 7608 17582 7655 17634
rect 7655 17582 7660 17634
rect 7472 17518 7477 17570
rect 7477 17518 7524 17570
rect 7540 17518 7592 17570
rect 7608 17518 7655 17570
rect 7655 17518 7660 17570
rect 7472 17454 7477 17506
rect 7477 17454 7524 17506
rect 7540 17454 7592 17506
rect 7608 17454 7655 17506
rect 7655 17454 7660 17506
rect 7472 17390 7477 17442
rect 7477 17390 7524 17442
rect 7540 17390 7592 17442
rect 7608 17390 7655 17442
rect 7655 17390 7660 17442
rect 7472 17326 7477 17378
rect 7477 17326 7524 17378
rect 7540 17326 7592 17378
rect 7608 17326 7655 17378
rect 7655 17326 7660 17378
rect 7472 17262 7477 17314
rect 7477 17262 7524 17314
rect 7540 17262 7592 17314
rect 7608 17262 7655 17314
rect 7655 17262 7660 17314
rect 7472 17198 7477 17250
rect 7477 17198 7524 17250
rect 7540 17198 7592 17250
rect 7608 17198 7655 17250
rect 7655 17198 7660 17250
rect 7472 17134 7477 17186
rect 7477 17134 7524 17186
rect 7540 17134 7592 17186
rect 7608 17134 7655 17186
rect 7655 17134 7660 17186
rect 7472 17070 7477 17122
rect 7477 17070 7524 17122
rect 7540 17070 7592 17122
rect 7608 17070 7655 17122
rect 7655 17070 7660 17122
rect 7472 17006 7477 17058
rect 7477 17006 7524 17058
rect 7540 17006 7592 17058
rect 7608 17006 7655 17058
rect 7655 17006 7660 17058
rect 7472 16942 7477 16994
rect 7477 16942 7524 16994
rect 7540 16942 7592 16994
rect 7608 16942 7655 16994
rect 7655 16942 7660 16994
rect 7472 16877 7477 16929
rect 7477 16877 7524 16929
rect 7540 16877 7592 16929
rect 7608 16877 7655 16929
rect 7655 16877 7660 16929
rect 7472 16812 7477 16864
rect 7477 16812 7524 16864
rect 7540 16812 7592 16864
rect 7608 16812 7655 16864
rect 7655 16812 7660 16864
rect 7472 16747 7477 16799
rect 7477 16747 7524 16799
rect 7540 16747 7592 16799
rect 7608 16747 7655 16799
rect 7655 16747 7660 16799
rect 7472 16682 7477 16734
rect 7477 16682 7524 16734
rect 7540 16682 7592 16734
rect 7608 16682 7655 16734
rect 7655 16682 7660 16734
rect 7472 16617 7477 16669
rect 7477 16617 7524 16669
rect 7540 16617 7592 16669
rect 7608 16617 7655 16669
rect 7655 16617 7660 16669
rect 7472 16552 7477 16604
rect 7477 16552 7524 16604
rect 7540 16552 7592 16604
rect 7608 16552 7655 16604
rect 7655 16552 7660 16604
rect 7472 16487 7477 16539
rect 7477 16487 7524 16539
rect 7540 16487 7592 16539
rect 7608 16487 7655 16539
rect 7655 16487 7660 16539
rect 7472 16422 7477 16474
rect 7477 16422 7524 16474
rect 7540 16422 7592 16474
rect 7608 16422 7655 16474
rect 7655 16422 7660 16474
rect 7472 16357 7477 16409
rect 7477 16357 7524 16409
rect 7540 16357 7592 16409
rect 7608 16357 7655 16409
rect 7655 16357 7660 16409
rect 7472 16292 7477 16344
rect 7477 16292 7524 16344
rect 7540 16292 7592 16344
rect 7608 16292 7655 16344
rect 7655 16292 7660 16344
rect 7472 16227 7477 16279
rect 7477 16227 7524 16279
rect 7540 16227 7592 16279
rect 7608 16227 7655 16279
rect 7655 16227 7660 16279
rect 7472 16162 7477 16214
rect 7477 16162 7524 16214
rect 7540 16162 7592 16214
rect 7608 16162 7655 16214
rect 7655 16162 7660 16214
rect 7472 13238 7477 13290
rect 7477 13238 7524 13290
rect 7540 13238 7592 13290
rect 7608 13238 7655 13290
rect 7655 13238 7660 13290
rect 7472 13174 7477 13226
rect 7477 13174 7524 13226
rect 7540 13174 7592 13226
rect 7608 13174 7655 13226
rect 7655 13174 7660 13226
rect 7472 13110 7477 13162
rect 7477 13110 7524 13162
rect 7540 13110 7592 13162
rect 7608 13110 7655 13162
rect 7655 13110 7660 13162
rect 7472 13046 7477 13098
rect 7477 13046 7524 13098
rect 7540 13046 7592 13098
rect 7608 13046 7655 13098
rect 7655 13046 7660 13098
rect 7472 12982 7477 13034
rect 7477 12982 7524 13034
rect 7540 12982 7592 13034
rect 7608 12982 7655 13034
rect 7655 12982 7660 13034
rect 7472 12918 7477 12970
rect 7477 12918 7524 12970
rect 7540 12918 7592 12970
rect 7608 12918 7655 12970
rect 7655 12918 7660 12970
rect 7472 12854 7477 12906
rect 7477 12854 7524 12906
rect 7540 12854 7592 12906
rect 7608 12854 7655 12906
rect 7655 12854 7660 12906
rect 7472 12790 7477 12842
rect 7477 12790 7524 12842
rect 7540 12790 7592 12842
rect 7608 12790 7655 12842
rect 7655 12790 7660 12842
rect 7472 12726 7477 12778
rect 7477 12726 7524 12778
rect 7540 12726 7592 12778
rect 7608 12726 7655 12778
rect 7655 12726 7660 12778
rect 7472 12662 7477 12714
rect 7477 12662 7524 12714
rect 7540 12662 7592 12714
rect 7608 12662 7655 12714
rect 7655 12662 7660 12714
rect 7472 12598 7477 12650
rect 7477 12598 7524 12650
rect 7540 12598 7592 12650
rect 7608 12598 7655 12650
rect 7655 12598 7660 12650
rect 7472 12534 7477 12586
rect 7477 12534 7524 12586
rect 7540 12534 7592 12586
rect 7608 12534 7655 12586
rect 7655 12534 7660 12586
rect 7472 12470 7477 12522
rect 7477 12470 7524 12522
rect 7540 12470 7592 12522
rect 7608 12470 7655 12522
rect 7655 12470 7660 12522
rect 7472 12406 7477 12458
rect 7477 12406 7524 12458
rect 7540 12406 7592 12458
rect 7608 12406 7655 12458
rect 7655 12406 7660 12458
rect 7472 12342 7477 12394
rect 7477 12342 7524 12394
rect 7540 12342 7592 12394
rect 7608 12342 7655 12394
rect 7655 12342 7660 12394
rect 7472 12277 7477 12329
rect 7477 12277 7524 12329
rect 7540 12277 7592 12329
rect 7608 12277 7655 12329
rect 7655 12277 7660 12329
rect 7472 12212 7477 12264
rect 7477 12212 7524 12264
rect 7540 12212 7592 12264
rect 7608 12212 7655 12264
rect 7655 12212 7660 12264
rect 7472 12147 7477 12199
rect 7477 12147 7524 12199
rect 7540 12147 7592 12199
rect 7608 12147 7655 12199
rect 7655 12147 7660 12199
rect 7472 12082 7477 12134
rect 7477 12082 7524 12134
rect 7540 12082 7592 12134
rect 7608 12082 7655 12134
rect 7655 12082 7660 12134
rect 7472 12017 7477 12069
rect 7477 12017 7524 12069
rect 7540 12017 7592 12069
rect 7608 12017 7655 12069
rect 7655 12017 7660 12069
rect 7472 11952 7477 12004
rect 7477 11952 7524 12004
rect 7540 11952 7592 12004
rect 7608 11952 7655 12004
rect 7655 11952 7660 12004
rect 7472 11887 7477 11939
rect 7477 11887 7524 11939
rect 7540 11887 7592 11939
rect 7608 11887 7655 11939
rect 7655 11887 7660 11939
rect 7472 11822 7477 11874
rect 7477 11822 7524 11874
rect 7540 11822 7592 11874
rect 7608 11822 7655 11874
rect 7655 11822 7660 11874
rect 7472 11757 7477 11809
rect 7477 11757 7524 11809
rect 7540 11757 7592 11809
rect 7608 11757 7655 11809
rect 7655 11757 7660 11809
rect 7472 11692 7477 11744
rect 7477 11692 7524 11744
rect 7540 11692 7592 11744
rect 7608 11692 7655 11744
rect 7655 11692 7660 11744
rect 7472 11627 7477 11679
rect 7477 11627 7524 11679
rect 7540 11627 7592 11679
rect 7608 11627 7655 11679
rect 7655 11627 7660 11679
rect 7472 11562 7477 11614
rect 7477 11562 7524 11614
rect 7540 11562 7592 11614
rect 7608 11562 7655 11614
rect 7655 11562 7660 11614
rect 7961 37945 8013 37997
rect 8039 37945 8091 37997
rect 7961 37877 8013 37929
rect 8039 37877 8091 37929
rect 7961 37809 8013 37861
rect 8039 37809 8091 37861
rect 7961 37741 8013 37793
rect 8039 37741 8091 37793
rect 7961 37673 8013 37725
rect 8039 37673 8091 37725
rect 7961 37605 8013 37657
rect 8039 37605 8091 37657
rect 7961 37537 8013 37589
rect 8039 37537 8091 37589
rect 7961 37469 8013 37521
rect 8039 37469 8091 37521
rect 7961 37401 8013 37453
rect 8039 37401 8091 37453
rect 7961 37333 8013 37385
rect 8039 37333 8091 37385
rect 7961 37266 8013 37318
rect 8039 37266 8091 37318
rect 7961 37199 8013 37251
rect 8039 37199 8091 37251
rect 7961 37132 8013 37184
rect 8039 37132 8091 37184
rect 7961 37065 8013 37117
rect 8039 37065 8091 37117
rect 7961 34173 8013 34225
rect 8039 34173 8091 34225
rect 7961 34109 8013 34161
rect 8039 34109 8091 34161
rect 7961 34045 8013 34097
rect 8039 34045 8091 34097
rect 7961 33981 8013 34033
rect 8039 33981 8091 34033
rect 7961 33917 8013 33969
rect 8039 33917 8091 33969
rect 7961 33853 8013 33905
rect 8039 33853 8091 33905
rect 7961 33789 8013 33841
rect 8039 33789 8091 33841
rect 7961 33725 8013 33777
rect 8039 33725 8091 33777
rect 7961 33661 8013 33713
rect 8039 33661 8091 33713
rect 7961 33597 8013 33649
rect 8039 33597 8091 33649
rect 7961 33533 8013 33585
rect 8039 33533 8091 33585
rect 7961 33469 8013 33521
rect 8039 33469 8091 33521
rect 7961 33405 8013 33457
rect 8039 33405 8091 33457
rect 7961 33341 8013 33393
rect 8039 33341 8091 33393
rect 7961 33277 8013 33329
rect 8039 33277 8091 33329
rect 7961 33212 8013 33264
rect 8039 33212 8091 33264
rect 7961 33147 8013 33199
rect 8039 33147 8091 33199
rect 7961 33082 8013 33134
rect 8039 33082 8091 33134
rect 7961 33017 8013 33069
rect 8039 33017 8091 33069
rect 7961 32952 8013 33004
rect 8039 32952 8091 33004
rect 7961 32887 8013 32939
rect 8039 32887 8091 32939
rect 7961 32822 8013 32874
rect 8039 32822 8091 32874
rect 7961 32757 8013 32809
rect 8039 32757 8091 32809
rect 7961 32692 8013 32744
rect 8039 32692 8091 32744
rect 7961 32627 8013 32679
rect 8039 32627 8091 32679
rect 7961 32562 8013 32614
rect 8039 32562 8091 32614
rect 7961 32497 8013 32549
rect 8039 32497 8091 32549
rect 7961 29573 8013 29625
rect 8039 29573 8091 29625
rect 7961 29509 8013 29561
rect 8039 29509 8091 29561
rect 7961 29445 8013 29497
rect 8039 29445 8091 29497
rect 7961 29381 8013 29433
rect 8039 29381 8091 29433
rect 7961 29317 8013 29369
rect 8039 29317 8091 29369
rect 7961 29253 8013 29305
rect 8039 29253 8091 29305
rect 7961 29189 8013 29241
rect 8039 29189 8091 29241
rect 7961 29125 8013 29177
rect 8039 29125 8091 29177
rect 7961 29061 8013 29113
rect 8039 29061 8091 29113
rect 7961 28997 8013 29049
rect 8039 28997 8091 29049
rect 7961 28933 8013 28985
rect 8039 28933 8091 28985
rect 7961 28869 8013 28921
rect 8039 28869 8091 28921
rect 7961 28805 8013 28857
rect 8039 28805 8091 28857
rect 7961 28741 8013 28793
rect 8039 28741 8091 28793
rect 7961 28677 8013 28729
rect 8039 28677 8091 28729
rect 7961 28612 8013 28664
rect 8039 28612 8091 28664
rect 7961 28547 8013 28599
rect 8039 28547 8091 28599
rect 7961 28482 8013 28534
rect 8039 28482 8091 28534
rect 7961 28417 8013 28469
rect 8039 28417 8091 28469
rect 7961 28352 8013 28404
rect 8039 28352 8091 28404
rect 7961 28287 8013 28339
rect 8039 28287 8091 28339
rect 7961 28222 8013 28274
rect 8039 28222 8091 28274
rect 7961 28157 8013 28209
rect 8039 28157 8091 28209
rect 7961 28092 8013 28144
rect 8039 28092 8091 28144
rect 7961 28027 8013 28079
rect 8039 28027 8091 28079
rect 7961 27962 8013 28014
rect 8039 27962 8091 28014
rect 7961 27897 8013 27949
rect 8039 27897 8091 27949
rect 7961 24973 8013 25025
rect 8039 24973 8091 25025
rect 7961 24909 8013 24961
rect 8039 24909 8091 24961
rect 7961 24845 8013 24897
rect 8039 24845 8091 24897
rect 7961 24781 8013 24833
rect 8039 24781 8091 24833
rect 7961 24717 8013 24769
rect 8039 24717 8091 24769
rect 7961 24653 8013 24705
rect 8039 24653 8091 24705
rect 7961 24589 8013 24641
rect 8039 24589 8091 24641
rect 7961 24525 8013 24577
rect 8039 24525 8091 24577
rect 7961 24461 8013 24513
rect 8039 24461 8091 24513
rect 7961 24397 8013 24449
rect 8039 24397 8091 24449
rect 7961 24333 8013 24385
rect 8039 24333 8091 24385
rect 7961 24269 8013 24321
rect 8039 24269 8091 24321
rect 7961 24205 8013 24257
rect 8039 24205 8091 24257
rect 7961 24141 8013 24193
rect 8039 24141 8091 24193
rect 7961 24077 8013 24129
rect 8039 24077 8091 24129
rect 7961 24012 8013 24064
rect 8039 24012 8091 24064
rect 7961 23947 8013 23999
rect 8039 23947 8091 23999
rect 7961 23882 8013 23934
rect 8039 23882 8091 23934
rect 7961 23817 8013 23869
rect 8039 23817 8091 23869
rect 7961 23752 8013 23804
rect 8039 23752 8091 23804
rect 7961 23687 8013 23739
rect 8039 23687 8091 23739
rect 7961 23622 8013 23674
rect 8039 23622 8091 23674
rect 7961 23557 8013 23609
rect 8039 23557 8091 23609
rect 7961 23492 8013 23544
rect 8039 23492 8091 23544
rect 7961 23427 8013 23479
rect 8039 23427 8091 23479
rect 7961 23362 8013 23414
rect 8039 23362 8091 23414
rect 7961 23297 8013 23349
rect 8039 23297 8091 23349
rect 7961 20373 8013 20425
rect 8039 20373 8091 20425
rect 7961 20309 8013 20361
rect 8039 20309 8091 20361
rect 7961 20245 8013 20297
rect 8039 20245 8091 20297
rect 7961 20181 8013 20233
rect 8039 20181 8091 20233
rect 7961 20117 8013 20169
rect 8039 20117 8091 20169
rect 7961 20053 8013 20105
rect 8039 20053 8091 20105
rect 7961 19989 8013 20041
rect 8039 19989 8091 20041
rect 7961 19925 8013 19977
rect 8039 19925 8091 19977
rect 7961 19861 8013 19913
rect 8039 19861 8091 19913
rect 7961 19797 8013 19849
rect 8039 19797 8091 19849
rect 7961 19733 8013 19785
rect 8039 19733 8091 19785
rect 7961 19669 8013 19721
rect 8039 19669 8091 19721
rect 7961 19605 8013 19657
rect 8039 19605 8091 19657
rect 7961 19541 8013 19593
rect 8039 19541 8091 19593
rect 7961 19477 8013 19529
rect 8039 19477 8091 19529
rect 7961 19412 8013 19464
rect 8039 19412 8091 19464
rect 7961 19347 8013 19399
rect 8039 19347 8091 19399
rect 7961 19282 8013 19334
rect 8039 19282 8091 19334
rect 7961 19217 8013 19269
rect 8039 19217 8091 19269
rect 7961 19152 8013 19204
rect 8039 19152 8091 19204
rect 7961 19087 8013 19139
rect 8039 19087 8091 19139
rect 7961 19022 8013 19074
rect 8039 19022 8091 19074
rect 7961 18957 8013 19009
rect 8039 18957 8091 19009
rect 7961 18892 8013 18944
rect 8039 18892 8091 18944
rect 7961 18827 8013 18879
rect 8039 18827 8091 18879
rect 7961 18762 8013 18814
rect 8039 18762 8091 18814
rect 7961 18697 8013 18749
rect 8039 18697 8091 18749
rect 7961 15773 8013 15825
rect 8039 15773 8091 15825
rect 7961 15709 8013 15761
rect 8039 15709 8091 15761
rect 7961 15645 8013 15697
rect 8039 15645 8091 15697
rect 7961 15581 8013 15633
rect 8039 15581 8091 15633
rect 7961 15517 8013 15569
rect 8039 15517 8091 15569
rect 7961 15453 8013 15505
rect 8039 15453 8091 15505
rect 7961 15389 8013 15441
rect 8039 15389 8091 15441
rect 7961 15325 8013 15377
rect 8039 15325 8091 15377
rect 7961 15261 8013 15313
rect 8039 15261 8091 15313
rect 7961 15197 8013 15249
rect 8039 15197 8091 15249
rect 7961 15133 8013 15185
rect 8039 15133 8091 15185
rect 7961 15069 8013 15121
rect 8039 15069 8091 15121
rect 7961 15005 8013 15057
rect 8039 15005 8091 15057
rect 7961 14941 8013 14993
rect 8039 14941 8091 14993
rect 7961 14877 8013 14929
rect 8039 14877 8091 14929
rect 7961 14812 8013 14864
rect 8039 14812 8091 14864
rect 7961 14747 8013 14799
rect 8039 14747 8091 14799
rect 7961 14682 8013 14734
rect 8039 14682 8091 14734
rect 7961 14617 8013 14669
rect 8039 14617 8091 14669
rect 7961 14552 8013 14604
rect 8039 14552 8091 14604
rect 7961 14487 8013 14539
rect 8039 14487 8091 14539
rect 7961 14422 8013 14474
rect 8039 14422 8091 14474
rect 7961 14357 8013 14409
rect 8039 14357 8091 14409
rect 7961 14292 8013 14344
rect 8039 14292 8091 14344
rect 7961 14227 8013 14279
rect 8039 14227 8091 14279
rect 7961 14162 8013 14214
rect 8039 14162 8091 14214
rect 7961 14097 8013 14149
rect 8039 14097 8091 14149
rect 7961 11173 8013 11225
rect 8039 11173 8091 11225
rect 7961 11109 8013 11161
rect 8039 11109 8091 11161
rect 7961 11045 8013 11097
rect 8039 11045 8091 11097
rect 7961 10981 8013 11033
rect 8039 10981 8091 11033
rect 7961 10917 8013 10969
rect 8039 10917 8091 10969
rect 7961 10853 8013 10905
rect 8039 10853 8091 10905
rect 7961 10789 8013 10841
rect 8039 10789 8091 10841
rect 7961 10725 8013 10777
rect 8039 10725 8091 10777
rect 7961 10661 8013 10713
rect 8039 10661 8091 10713
rect 7961 10597 8013 10649
rect 8039 10597 8091 10649
rect 7961 10533 8013 10585
rect 8039 10533 8091 10585
rect 7961 10469 8013 10521
rect 8039 10469 8091 10521
rect 7961 10405 8013 10457
rect 8039 10405 8091 10457
rect 7961 10341 8013 10393
rect 8039 10341 8091 10393
rect 7961 10277 8013 10329
rect 8039 10277 8091 10329
rect 7961 10212 8013 10264
rect 8039 10212 8091 10264
rect 7961 10147 8013 10199
rect 8039 10147 8091 10199
rect 7961 10082 8013 10134
rect 8039 10082 8091 10134
rect 7961 10017 8013 10069
rect 8039 10017 8091 10069
rect 7961 9952 8013 10004
rect 8039 9952 8091 10004
rect 7961 9887 8013 9939
rect 8039 9887 8091 9939
rect 7961 9822 8013 9874
rect 8039 9822 8091 9874
rect 7961 9757 8013 9809
rect 8039 9757 8091 9809
rect 7961 9692 8013 9744
rect 8039 9692 8091 9744
rect 7961 9627 8013 9679
rect 8039 9627 8091 9679
rect 7961 9562 8013 9614
rect 8039 9562 8091 9614
rect 7961 9497 8013 9549
rect 8039 9497 8091 9549
rect 8392 36238 8397 36290
rect 8397 36238 8444 36290
rect 8460 36238 8512 36290
rect 8528 36238 8575 36290
rect 8575 36238 8580 36290
rect 8392 36174 8397 36226
rect 8397 36174 8444 36226
rect 8460 36174 8512 36226
rect 8528 36174 8575 36226
rect 8575 36174 8580 36226
rect 8392 36110 8397 36162
rect 8397 36110 8444 36162
rect 8460 36110 8512 36162
rect 8528 36110 8575 36162
rect 8575 36110 8580 36162
rect 8392 36046 8397 36098
rect 8397 36046 8444 36098
rect 8460 36046 8512 36098
rect 8528 36046 8575 36098
rect 8575 36046 8580 36098
rect 8392 35982 8397 36034
rect 8397 35982 8444 36034
rect 8460 35982 8512 36034
rect 8528 35982 8575 36034
rect 8575 35982 8580 36034
rect 8392 35918 8397 35970
rect 8397 35918 8444 35970
rect 8460 35918 8512 35970
rect 8528 35918 8575 35970
rect 8575 35918 8580 35970
rect 8392 35854 8397 35906
rect 8397 35854 8444 35906
rect 8460 35854 8512 35906
rect 8528 35854 8575 35906
rect 8575 35854 8580 35906
rect 8392 35790 8397 35842
rect 8397 35790 8444 35842
rect 8460 35790 8512 35842
rect 8528 35790 8575 35842
rect 8575 35790 8580 35842
rect 8392 35726 8397 35778
rect 8397 35726 8444 35778
rect 8460 35726 8512 35778
rect 8528 35726 8575 35778
rect 8575 35726 8580 35778
rect 8392 35662 8397 35714
rect 8397 35662 8444 35714
rect 8460 35662 8512 35714
rect 8528 35662 8575 35714
rect 8575 35662 8580 35714
rect 8392 35598 8397 35650
rect 8397 35598 8444 35650
rect 8460 35598 8512 35650
rect 8528 35598 8575 35650
rect 8575 35598 8580 35650
rect 8392 35534 8397 35586
rect 8397 35534 8444 35586
rect 8460 35534 8512 35586
rect 8528 35534 8575 35586
rect 8575 35534 8580 35586
rect 8392 35470 8397 35522
rect 8397 35470 8444 35522
rect 8460 35470 8512 35522
rect 8528 35470 8575 35522
rect 8575 35470 8580 35522
rect 8392 35406 8397 35458
rect 8397 35406 8444 35458
rect 8460 35406 8512 35458
rect 8528 35406 8575 35458
rect 8575 35406 8580 35458
rect 8392 35342 8397 35394
rect 8397 35342 8444 35394
rect 8460 35342 8512 35394
rect 8528 35342 8575 35394
rect 8575 35342 8580 35394
rect 8392 35277 8397 35329
rect 8397 35277 8444 35329
rect 8460 35277 8512 35329
rect 8528 35277 8575 35329
rect 8575 35277 8580 35329
rect 8392 35212 8397 35264
rect 8397 35212 8444 35264
rect 8460 35212 8512 35264
rect 8528 35212 8575 35264
rect 8575 35212 8580 35264
rect 8392 35147 8397 35199
rect 8397 35147 8444 35199
rect 8460 35147 8512 35199
rect 8528 35147 8575 35199
rect 8575 35147 8580 35199
rect 8392 35082 8397 35134
rect 8397 35082 8444 35134
rect 8460 35082 8512 35134
rect 8528 35082 8575 35134
rect 8575 35082 8580 35134
rect 8392 35017 8397 35069
rect 8397 35017 8444 35069
rect 8460 35017 8512 35069
rect 8528 35017 8575 35069
rect 8575 35017 8580 35069
rect 8392 34952 8397 35004
rect 8397 34952 8444 35004
rect 8460 34952 8512 35004
rect 8528 34952 8575 35004
rect 8575 34952 8580 35004
rect 8392 34887 8397 34939
rect 8397 34887 8444 34939
rect 8460 34887 8512 34939
rect 8528 34887 8575 34939
rect 8575 34887 8580 34939
rect 8392 34822 8397 34874
rect 8397 34822 8444 34874
rect 8460 34822 8512 34874
rect 8528 34822 8575 34874
rect 8575 34822 8580 34874
rect 8392 34757 8397 34809
rect 8397 34757 8444 34809
rect 8460 34757 8512 34809
rect 8528 34757 8575 34809
rect 8575 34757 8580 34809
rect 8392 34692 8397 34744
rect 8397 34692 8444 34744
rect 8460 34692 8512 34744
rect 8528 34692 8575 34744
rect 8575 34692 8580 34744
rect 8392 34627 8397 34679
rect 8397 34627 8444 34679
rect 8460 34627 8512 34679
rect 8528 34627 8575 34679
rect 8575 34627 8580 34679
rect 8392 34562 8397 34614
rect 8397 34562 8444 34614
rect 8460 34562 8512 34614
rect 8528 34562 8575 34614
rect 8575 34562 8580 34614
rect 8392 31638 8397 31690
rect 8397 31638 8444 31690
rect 8460 31638 8512 31690
rect 8528 31638 8575 31690
rect 8575 31638 8580 31690
rect 8392 31574 8397 31626
rect 8397 31574 8444 31626
rect 8460 31574 8512 31626
rect 8528 31574 8575 31626
rect 8575 31574 8580 31626
rect 8392 31510 8397 31562
rect 8397 31510 8444 31562
rect 8460 31510 8512 31562
rect 8528 31510 8575 31562
rect 8575 31510 8580 31562
rect 8392 31446 8397 31498
rect 8397 31446 8444 31498
rect 8460 31446 8512 31498
rect 8528 31446 8575 31498
rect 8575 31446 8580 31498
rect 8392 31382 8397 31434
rect 8397 31382 8444 31434
rect 8460 31382 8512 31434
rect 8528 31382 8575 31434
rect 8575 31382 8580 31434
rect 8392 31318 8397 31370
rect 8397 31318 8444 31370
rect 8460 31318 8512 31370
rect 8528 31318 8575 31370
rect 8575 31318 8580 31370
rect 8392 31254 8397 31306
rect 8397 31254 8444 31306
rect 8460 31254 8512 31306
rect 8528 31254 8575 31306
rect 8575 31254 8580 31306
rect 8392 31190 8397 31242
rect 8397 31190 8444 31242
rect 8460 31190 8512 31242
rect 8528 31190 8575 31242
rect 8575 31190 8580 31242
rect 8392 31126 8397 31178
rect 8397 31126 8444 31178
rect 8460 31126 8512 31178
rect 8528 31126 8575 31178
rect 8575 31126 8580 31178
rect 8392 31062 8397 31114
rect 8397 31062 8444 31114
rect 8460 31062 8512 31114
rect 8528 31062 8575 31114
rect 8575 31062 8580 31114
rect 8392 30998 8397 31050
rect 8397 30998 8444 31050
rect 8460 30998 8512 31050
rect 8528 30998 8575 31050
rect 8575 30998 8580 31050
rect 8392 30934 8397 30986
rect 8397 30934 8444 30986
rect 8460 30934 8512 30986
rect 8528 30934 8575 30986
rect 8575 30934 8580 30986
rect 8392 30870 8397 30922
rect 8397 30870 8444 30922
rect 8460 30870 8512 30922
rect 8528 30870 8575 30922
rect 8575 30870 8580 30922
rect 8392 30806 8397 30858
rect 8397 30806 8444 30858
rect 8460 30806 8512 30858
rect 8528 30806 8575 30858
rect 8575 30806 8580 30858
rect 8392 30742 8397 30794
rect 8397 30742 8444 30794
rect 8460 30742 8512 30794
rect 8528 30742 8575 30794
rect 8575 30742 8580 30794
rect 8392 30677 8397 30729
rect 8397 30677 8444 30729
rect 8460 30677 8512 30729
rect 8528 30677 8575 30729
rect 8575 30677 8580 30729
rect 8392 30612 8397 30664
rect 8397 30612 8444 30664
rect 8460 30612 8512 30664
rect 8528 30612 8575 30664
rect 8575 30612 8580 30664
rect 8392 30547 8397 30599
rect 8397 30547 8444 30599
rect 8460 30547 8512 30599
rect 8528 30547 8575 30599
rect 8575 30547 8580 30599
rect 8392 30482 8397 30534
rect 8397 30482 8444 30534
rect 8460 30482 8512 30534
rect 8528 30482 8575 30534
rect 8575 30482 8580 30534
rect 8392 30417 8397 30469
rect 8397 30417 8444 30469
rect 8460 30417 8512 30469
rect 8528 30417 8575 30469
rect 8575 30417 8580 30469
rect 8392 30352 8397 30404
rect 8397 30352 8444 30404
rect 8460 30352 8512 30404
rect 8528 30352 8575 30404
rect 8575 30352 8580 30404
rect 8392 30287 8397 30339
rect 8397 30287 8444 30339
rect 8460 30287 8512 30339
rect 8528 30287 8575 30339
rect 8575 30287 8580 30339
rect 8392 30222 8397 30274
rect 8397 30222 8444 30274
rect 8460 30222 8512 30274
rect 8528 30222 8575 30274
rect 8575 30222 8580 30274
rect 8392 30157 8397 30209
rect 8397 30157 8444 30209
rect 8460 30157 8512 30209
rect 8528 30157 8575 30209
rect 8575 30157 8580 30209
rect 8392 30092 8397 30144
rect 8397 30092 8444 30144
rect 8460 30092 8512 30144
rect 8528 30092 8575 30144
rect 8575 30092 8580 30144
rect 8392 30027 8397 30079
rect 8397 30027 8444 30079
rect 8460 30027 8512 30079
rect 8528 30027 8575 30079
rect 8575 30027 8580 30079
rect 8392 29962 8397 30014
rect 8397 29962 8444 30014
rect 8460 29962 8512 30014
rect 8528 29962 8575 30014
rect 8575 29962 8580 30014
rect 8392 27038 8397 27090
rect 8397 27038 8444 27090
rect 8460 27038 8512 27090
rect 8528 27038 8575 27090
rect 8575 27038 8580 27090
rect 8392 26974 8397 27026
rect 8397 26974 8444 27026
rect 8460 26974 8512 27026
rect 8528 26974 8575 27026
rect 8575 26974 8580 27026
rect 8392 26910 8397 26962
rect 8397 26910 8444 26962
rect 8460 26910 8512 26962
rect 8528 26910 8575 26962
rect 8575 26910 8580 26962
rect 8392 26846 8397 26898
rect 8397 26846 8444 26898
rect 8460 26846 8512 26898
rect 8528 26846 8575 26898
rect 8575 26846 8580 26898
rect 8392 26782 8397 26834
rect 8397 26782 8444 26834
rect 8460 26782 8512 26834
rect 8528 26782 8575 26834
rect 8575 26782 8580 26834
rect 8392 26718 8397 26770
rect 8397 26718 8444 26770
rect 8460 26718 8512 26770
rect 8528 26718 8575 26770
rect 8575 26718 8580 26770
rect 8392 26654 8397 26706
rect 8397 26654 8444 26706
rect 8460 26654 8512 26706
rect 8528 26654 8575 26706
rect 8575 26654 8580 26706
rect 8392 26590 8397 26642
rect 8397 26590 8444 26642
rect 8460 26590 8512 26642
rect 8528 26590 8575 26642
rect 8575 26590 8580 26642
rect 8392 26526 8397 26578
rect 8397 26526 8444 26578
rect 8460 26526 8512 26578
rect 8528 26526 8575 26578
rect 8575 26526 8580 26578
rect 8392 26462 8397 26514
rect 8397 26462 8444 26514
rect 8460 26462 8512 26514
rect 8528 26462 8575 26514
rect 8575 26462 8580 26514
rect 8392 26398 8397 26450
rect 8397 26398 8444 26450
rect 8460 26398 8512 26450
rect 8528 26398 8575 26450
rect 8575 26398 8580 26450
rect 8392 26334 8397 26386
rect 8397 26334 8444 26386
rect 8460 26334 8512 26386
rect 8528 26334 8575 26386
rect 8575 26334 8580 26386
rect 8392 26270 8397 26322
rect 8397 26270 8444 26322
rect 8460 26270 8512 26322
rect 8528 26270 8575 26322
rect 8575 26270 8580 26322
rect 8392 26206 8397 26258
rect 8397 26206 8444 26258
rect 8460 26206 8512 26258
rect 8528 26206 8575 26258
rect 8575 26206 8580 26258
rect 8392 26142 8397 26194
rect 8397 26142 8444 26194
rect 8460 26142 8512 26194
rect 8528 26142 8575 26194
rect 8575 26142 8580 26194
rect 8392 26077 8397 26129
rect 8397 26077 8444 26129
rect 8460 26077 8512 26129
rect 8528 26077 8575 26129
rect 8575 26077 8580 26129
rect 8392 26012 8397 26064
rect 8397 26012 8444 26064
rect 8460 26012 8512 26064
rect 8528 26012 8575 26064
rect 8575 26012 8580 26064
rect 8392 25947 8397 25999
rect 8397 25947 8444 25999
rect 8460 25947 8512 25999
rect 8528 25947 8575 25999
rect 8575 25947 8580 25999
rect 8392 25882 8397 25934
rect 8397 25882 8444 25934
rect 8460 25882 8512 25934
rect 8528 25882 8575 25934
rect 8575 25882 8580 25934
rect 8392 25817 8397 25869
rect 8397 25817 8444 25869
rect 8460 25817 8512 25869
rect 8528 25817 8575 25869
rect 8575 25817 8580 25869
rect 8392 25752 8397 25804
rect 8397 25752 8444 25804
rect 8460 25752 8512 25804
rect 8528 25752 8575 25804
rect 8575 25752 8580 25804
rect 8392 25687 8397 25739
rect 8397 25687 8444 25739
rect 8460 25687 8512 25739
rect 8528 25687 8575 25739
rect 8575 25687 8580 25739
rect 8392 25622 8397 25674
rect 8397 25622 8444 25674
rect 8460 25622 8512 25674
rect 8528 25622 8575 25674
rect 8575 25622 8580 25674
rect 8392 25557 8397 25609
rect 8397 25557 8444 25609
rect 8460 25557 8512 25609
rect 8528 25557 8575 25609
rect 8575 25557 8580 25609
rect 8392 25492 8397 25544
rect 8397 25492 8444 25544
rect 8460 25492 8512 25544
rect 8528 25492 8575 25544
rect 8575 25492 8580 25544
rect 8392 25427 8397 25479
rect 8397 25427 8444 25479
rect 8460 25427 8512 25479
rect 8528 25427 8575 25479
rect 8575 25427 8580 25479
rect 8392 25362 8397 25414
rect 8397 25362 8444 25414
rect 8460 25362 8512 25414
rect 8528 25362 8575 25414
rect 8575 25362 8580 25414
rect 8392 22438 8397 22490
rect 8397 22438 8444 22490
rect 8460 22438 8512 22490
rect 8528 22438 8575 22490
rect 8575 22438 8580 22490
rect 8392 22374 8397 22426
rect 8397 22374 8444 22426
rect 8460 22374 8512 22426
rect 8528 22374 8575 22426
rect 8575 22374 8580 22426
rect 8392 22310 8397 22362
rect 8397 22310 8444 22362
rect 8460 22310 8512 22362
rect 8528 22310 8575 22362
rect 8575 22310 8580 22362
rect 8392 22246 8397 22298
rect 8397 22246 8444 22298
rect 8460 22246 8512 22298
rect 8528 22246 8575 22298
rect 8575 22246 8580 22298
rect 8392 22182 8397 22234
rect 8397 22182 8444 22234
rect 8460 22182 8512 22234
rect 8528 22182 8575 22234
rect 8575 22182 8580 22234
rect 8392 22118 8397 22170
rect 8397 22118 8444 22170
rect 8460 22118 8512 22170
rect 8528 22118 8575 22170
rect 8575 22118 8580 22170
rect 8392 22054 8397 22106
rect 8397 22054 8444 22106
rect 8460 22054 8512 22106
rect 8528 22054 8575 22106
rect 8575 22054 8580 22106
rect 8392 21990 8397 22042
rect 8397 21990 8444 22042
rect 8460 21990 8512 22042
rect 8528 21990 8575 22042
rect 8575 21990 8580 22042
rect 8392 21926 8397 21978
rect 8397 21926 8444 21978
rect 8460 21926 8512 21978
rect 8528 21926 8575 21978
rect 8575 21926 8580 21978
rect 8392 21862 8397 21914
rect 8397 21862 8444 21914
rect 8460 21862 8512 21914
rect 8528 21862 8575 21914
rect 8575 21862 8580 21914
rect 8392 21798 8397 21850
rect 8397 21798 8444 21850
rect 8460 21798 8512 21850
rect 8528 21798 8575 21850
rect 8575 21798 8580 21850
rect 8392 21734 8397 21786
rect 8397 21734 8444 21786
rect 8460 21734 8512 21786
rect 8528 21734 8575 21786
rect 8575 21734 8580 21786
rect 8392 21670 8397 21722
rect 8397 21670 8444 21722
rect 8460 21670 8512 21722
rect 8528 21670 8575 21722
rect 8575 21670 8580 21722
rect 8392 21606 8397 21658
rect 8397 21606 8444 21658
rect 8460 21606 8512 21658
rect 8528 21606 8575 21658
rect 8575 21606 8580 21658
rect 8392 21542 8397 21594
rect 8397 21542 8444 21594
rect 8460 21542 8512 21594
rect 8528 21542 8575 21594
rect 8575 21542 8580 21594
rect 8392 21477 8397 21529
rect 8397 21477 8444 21529
rect 8460 21477 8512 21529
rect 8528 21477 8575 21529
rect 8575 21477 8580 21529
rect 8392 21412 8397 21464
rect 8397 21412 8444 21464
rect 8460 21412 8512 21464
rect 8528 21412 8575 21464
rect 8575 21412 8580 21464
rect 8392 21347 8397 21399
rect 8397 21347 8444 21399
rect 8460 21347 8512 21399
rect 8528 21347 8575 21399
rect 8575 21347 8580 21399
rect 8392 21282 8397 21334
rect 8397 21282 8444 21334
rect 8460 21282 8512 21334
rect 8528 21282 8575 21334
rect 8575 21282 8580 21334
rect 8392 21217 8397 21269
rect 8397 21217 8444 21269
rect 8460 21217 8512 21269
rect 8528 21217 8575 21269
rect 8575 21217 8580 21269
rect 8392 21152 8397 21204
rect 8397 21152 8444 21204
rect 8460 21152 8512 21204
rect 8528 21152 8575 21204
rect 8575 21152 8580 21204
rect 8392 21087 8397 21139
rect 8397 21087 8444 21139
rect 8460 21087 8512 21139
rect 8528 21087 8575 21139
rect 8575 21087 8580 21139
rect 8392 21022 8397 21074
rect 8397 21022 8444 21074
rect 8460 21022 8512 21074
rect 8528 21022 8575 21074
rect 8575 21022 8580 21074
rect 8392 20957 8397 21009
rect 8397 20957 8444 21009
rect 8460 20957 8512 21009
rect 8528 20957 8575 21009
rect 8575 20957 8580 21009
rect 8392 20892 8397 20944
rect 8397 20892 8444 20944
rect 8460 20892 8512 20944
rect 8528 20892 8575 20944
rect 8575 20892 8580 20944
rect 8392 20827 8397 20879
rect 8397 20827 8444 20879
rect 8460 20827 8512 20879
rect 8528 20827 8575 20879
rect 8575 20827 8580 20879
rect 8392 20762 8397 20814
rect 8397 20762 8444 20814
rect 8460 20762 8512 20814
rect 8528 20762 8575 20814
rect 8575 20762 8580 20814
rect 8392 17838 8397 17890
rect 8397 17838 8444 17890
rect 8460 17838 8512 17890
rect 8528 17838 8575 17890
rect 8575 17838 8580 17890
rect 8392 17774 8397 17826
rect 8397 17774 8444 17826
rect 8460 17774 8512 17826
rect 8528 17774 8575 17826
rect 8575 17774 8580 17826
rect 8392 17710 8397 17762
rect 8397 17710 8444 17762
rect 8460 17710 8512 17762
rect 8528 17710 8575 17762
rect 8575 17710 8580 17762
rect 8392 17646 8397 17698
rect 8397 17646 8444 17698
rect 8460 17646 8512 17698
rect 8528 17646 8575 17698
rect 8575 17646 8580 17698
rect 8392 17582 8397 17634
rect 8397 17582 8444 17634
rect 8460 17582 8512 17634
rect 8528 17582 8575 17634
rect 8575 17582 8580 17634
rect 8392 17518 8397 17570
rect 8397 17518 8444 17570
rect 8460 17518 8512 17570
rect 8528 17518 8575 17570
rect 8575 17518 8580 17570
rect 8392 17454 8397 17506
rect 8397 17454 8444 17506
rect 8460 17454 8512 17506
rect 8528 17454 8575 17506
rect 8575 17454 8580 17506
rect 8392 17390 8397 17442
rect 8397 17390 8444 17442
rect 8460 17390 8512 17442
rect 8528 17390 8575 17442
rect 8575 17390 8580 17442
rect 8392 17326 8397 17378
rect 8397 17326 8444 17378
rect 8460 17326 8512 17378
rect 8528 17326 8575 17378
rect 8575 17326 8580 17378
rect 8392 17262 8397 17314
rect 8397 17262 8444 17314
rect 8460 17262 8512 17314
rect 8528 17262 8575 17314
rect 8575 17262 8580 17314
rect 8392 17198 8397 17250
rect 8397 17198 8444 17250
rect 8460 17198 8512 17250
rect 8528 17198 8575 17250
rect 8575 17198 8580 17250
rect 8392 17134 8397 17186
rect 8397 17134 8444 17186
rect 8460 17134 8512 17186
rect 8528 17134 8575 17186
rect 8575 17134 8580 17186
rect 8392 17070 8397 17122
rect 8397 17070 8444 17122
rect 8460 17070 8512 17122
rect 8528 17070 8575 17122
rect 8575 17070 8580 17122
rect 8392 17006 8397 17058
rect 8397 17006 8444 17058
rect 8460 17006 8512 17058
rect 8528 17006 8575 17058
rect 8575 17006 8580 17058
rect 8392 16942 8397 16994
rect 8397 16942 8444 16994
rect 8460 16942 8512 16994
rect 8528 16942 8575 16994
rect 8575 16942 8580 16994
rect 8392 16877 8397 16929
rect 8397 16877 8444 16929
rect 8460 16877 8512 16929
rect 8528 16877 8575 16929
rect 8575 16877 8580 16929
rect 8392 16812 8397 16864
rect 8397 16812 8444 16864
rect 8460 16812 8512 16864
rect 8528 16812 8575 16864
rect 8575 16812 8580 16864
rect 8392 16747 8397 16799
rect 8397 16747 8444 16799
rect 8460 16747 8512 16799
rect 8528 16747 8575 16799
rect 8575 16747 8580 16799
rect 8392 16682 8397 16734
rect 8397 16682 8444 16734
rect 8460 16682 8512 16734
rect 8528 16682 8575 16734
rect 8575 16682 8580 16734
rect 8392 16617 8397 16669
rect 8397 16617 8444 16669
rect 8460 16617 8512 16669
rect 8528 16617 8575 16669
rect 8575 16617 8580 16669
rect 8392 16552 8397 16604
rect 8397 16552 8444 16604
rect 8460 16552 8512 16604
rect 8528 16552 8575 16604
rect 8575 16552 8580 16604
rect 8392 16487 8397 16539
rect 8397 16487 8444 16539
rect 8460 16487 8512 16539
rect 8528 16487 8575 16539
rect 8575 16487 8580 16539
rect 8392 16422 8397 16474
rect 8397 16422 8444 16474
rect 8460 16422 8512 16474
rect 8528 16422 8575 16474
rect 8575 16422 8580 16474
rect 8392 16357 8397 16409
rect 8397 16357 8444 16409
rect 8460 16357 8512 16409
rect 8528 16357 8575 16409
rect 8575 16357 8580 16409
rect 8392 16292 8397 16344
rect 8397 16292 8444 16344
rect 8460 16292 8512 16344
rect 8528 16292 8575 16344
rect 8575 16292 8580 16344
rect 8392 16227 8397 16279
rect 8397 16227 8444 16279
rect 8460 16227 8512 16279
rect 8528 16227 8575 16279
rect 8575 16227 8580 16279
rect 8392 16162 8397 16214
rect 8397 16162 8444 16214
rect 8460 16162 8512 16214
rect 8528 16162 8575 16214
rect 8575 16162 8580 16214
rect 8392 13238 8397 13290
rect 8397 13238 8444 13290
rect 8460 13238 8512 13290
rect 8528 13238 8575 13290
rect 8575 13238 8580 13290
rect 8392 13174 8397 13226
rect 8397 13174 8444 13226
rect 8460 13174 8512 13226
rect 8528 13174 8575 13226
rect 8575 13174 8580 13226
rect 8392 13110 8397 13162
rect 8397 13110 8444 13162
rect 8460 13110 8512 13162
rect 8528 13110 8575 13162
rect 8575 13110 8580 13162
rect 8392 13046 8397 13098
rect 8397 13046 8444 13098
rect 8460 13046 8512 13098
rect 8528 13046 8575 13098
rect 8575 13046 8580 13098
rect 8392 12982 8397 13034
rect 8397 12982 8444 13034
rect 8460 12982 8512 13034
rect 8528 12982 8575 13034
rect 8575 12982 8580 13034
rect 8392 12918 8397 12970
rect 8397 12918 8444 12970
rect 8460 12918 8512 12970
rect 8528 12918 8575 12970
rect 8575 12918 8580 12970
rect 8392 12854 8397 12906
rect 8397 12854 8444 12906
rect 8460 12854 8512 12906
rect 8528 12854 8575 12906
rect 8575 12854 8580 12906
rect 8392 12790 8397 12842
rect 8397 12790 8444 12842
rect 8460 12790 8512 12842
rect 8528 12790 8575 12842
rect 8575 12790 8580 12842
rect 8392 12726 8397 12778
rect 8397 12726 8444 12778
rect 8460 12726 8512 12778
rect 8528 12726 8575 12778
rect 8575 12726 8580 12778
rect 8392 12662 8397 12714
rect 8397 12662 8444 12714
rect 8460 12662 8512 12714
rect 8528 12662 8575 12714
rect 8575 12662 8580 12714
rect 8392 12598 8397 12650
rect 8397 12598 8444 12650
rect 8460 12598 8512 12650
rect 8528 12598 8575 12650
rect 8575 12598 8580 12650
rect 8392 12534 8397 12586
rect 8397 12534 8444 12586
rect 8460 12534 8512 12586
rect 8528 12534 8575 12586
rect 8575 12534 8580 12586
rect 8392 12470 8397 12522
rect 8397 12470 8444 12522
rect 8460 12470 8512 12522
rect 8528 12470 8575 12522
rect 8575 12470 8580 12522
rect 8392 12406 8397 12458
rect 8397 12406 8444 12458
rect 8460 12406 8512 12458
rect 8528 12406 8575 12458
rect 8575 12406 8580 12458
rect 8392 12342 8397 12394
rect 8397 12342 8444 12394
rect 8460 12342 8512 12394
rect 8528 12342 8575 12394
rect 8575 12342 8580 12394
rect 8392 12277 8397 12329
rect 8397 12277 8444 12329
rect 8460 12277 8512 12329
rect 8528 12277 8575 12329
rect 8575 12277 8580 12329
rect 8392 12212 8397 12264
rect 8397 12212 8444 12264
rect 8460 12212 8512 12264
rect 8528 12212 8575 12264
rect 8575 12212 8580 12264
rect 8392 12147 8397 12199
rect 8397 12147 8444 12199
rect 8460 12147 8512 12199
rect 8528 12147 8575 12199
rect 8575 12147 8580 12199
rect 8392 12082 8397 12134
rect 8397 12082 8444 12134
rect 8460 12082 8512 12134
rect 8528 12082 8575 12134
rect 8575 12082 8580 12134
rect 8392 12017 8397 12069
rect 8397 12017 8444 12069
rect 8460 12017 8512 12069
rect 8528 12017 8575 12069
rect 8575 12017 8580 12069
rect 8392 11952 8397 12004
rect 8397 11952 8444 12004
rect 8460 11952 8512 12004
rect 8528 11952 8575 12004
rect 8575 11952 8580 12004
rect 8392 11887 8397 11939
rect 8397 11887 8444 11939
rect 8460 11887 8512 11939
rect 8528 11887 8575 11939
rect 8575 11887 8580 11939
rect 8392 11822 8397 11874
rect 8397 11822 8444 11874
rect 8460 11822 8512 11874
rect 8528 11822 8575 11874
rect 8575 11822 8580 11874
rect 8392 11757 8397 11809
rect 8397 11757 8444 11809
rect 8460 11757 8512 11809
rect 8528 11757 8575 11809
rect 8575 11757 8580 11809
rect 8392 11692 8397 11744
rect 8397 11692 8444 11744
rect 8460 11692 8512 11744
rect 8528 11692 8575 11744
rect 8575 11692 8580 11744
rect 8392 11627 8397 11679
rect 8397 11627 8444 11679
rect 8460 11627 8512 11679
rect 8528 11627 8575 11679
rect 8575 11627 8580 11679
rect 8392 11562 8397 11614
rect 8397 11562 8444 11614
rect 8460 11562 8512 11614
rect 8528 11562 8575 11614
rect 8575 11562 8580 11614
rect 8881 37945 8933 37997
rect 8959 37945 9011 37997
rect 8881 37877 8933 37929
rect 8959 37877 9011 37929
rect 8881 37809 8933 37861
rect 8959 37809 9011 37861
rect 8881 37741 8933 37793
rect 8959 37741 9011 37793
rect 8881 37673 8933 37725
rect 8959 37673 9011 37725
rect 8881 37605 8933 37657
rect 8959 37605 9011 37657
rect 8881 37537 8933 37589
rect 8959 37537 9011 37589
rect 8881 37469 8933 37521
rect 8959 37469 9011 37521
rect 8881 37401 8933 37453
rect 8959 37401 9011 37453
rect 8881 37333 8933 37385
rect 8959 37333 9011 37385
rect 8881 37266 8933 37318
rect 8959 37266 9011 37318
rect 8881 37199 8933 37251
rect 8959 37199 9011 37251
rect 8881 37132 8933 37184
rect 8959 37132 9011 37184
rect 8881 37065 8933 37117
rect 8959 37065 9011 37117
rect 8881 34173 8933 34225
rect 8959 34173 9011 34225
rect 8881 34109 8933 34161
rect 8959 34109 9011 34161
rect 8881 34045 8933 34097
rect 8959 34045 9011 34097
rect 8881 33981 8933 34033
rect 8959 33981 9011 34033
rect 8881 33917 8933 33969
rect 8959 33917 9011 33969
rect 8881 33853 8933 33905
rect 8959 33853 9011 33905
rect 8881 33789 8933 33841
rect 8959 33789 9011 33841
rect 8881 33725 8933 33777
rect 8959 33725 9011 33777
rect 8881 33661 8933 33713
rect 8959 33661 9011 33713
rect 8881 33597 8933 33649
rect 8959 33597 9011 33649
rect 8881 33533 8933 33585
rect 8959 33533 9011 33585
rect 8881 33469 8933 33521
rect 8959 33469 9011 33521
rect 8881 33405 8933 33457
rect 8959 33405 9011 33457
rect 8881 33341 8933 33393
rect 8959 33341 9011 33393
rect 8881 33277 8933 33329
rect 8959 33277 9011 33329
rect 8881 33212 8933 33264
rect 8959 33212 9011 33264
rect 8881 33147 8933 33199
rect 8959 33147 9011 33199
rect 8881 33082 8933 33134
rect 8959 33082 9011 33134
rect 8881 33017 8933 33069
rect 8959 33017 9011 33069
rect 8881 32952 8933 33004
rect 8959 32952 9011 33004
rect 8881 32887 8933 32939
rect 8959 32887 9011 32939
rect 8881 32822 8933 32874
rect 8959 32822 9011 32874
rect 8881 32757 8933 32809
rect 8959 32757 9011 32809
rect 8881 32692 8933 32744
rect 8959 32692 9011 32744
rect 8881 32627 8933 32679
rect 8959 32627 9011 32679
rect 8881 32562 8933 32614
rect 8959 32562 9011 32614
rect 8881 32497 8933 32549
rect 8959 32497 9011 32549
rect 8881 29573 8933 29625
rect 8959 29573 9011 29625
rect 8881 29509 8933 29561
rect 8959 29509 9011 29561
rect 8881 29445 8933 29497
rect 8959 29445 9011 29497
rect 8881 29381 8933 29433
rect 8959 29381 9011 29433
rect 8881 29317 8933 29369
rect 8959 29317 9011 29369
rect 8881 29253 8933 29305
rect 8959 29253 9011 29305
rect 8881 29189 8933 29241
rect 8959 29189 9011 29241
rect 8881 29125 8933 29177
rect 8959 29125 9011 29177
rect 8881 29061 8933 29113
rect 8959 29061 9011 29113
rect 8881 28997 8933 29049
rect 8959 28997 9011 29049
rect 8881 28933 8933 28985
rect 8959 28933 9011 28985
rect 8881 28869 8933 28921
rect 8959 28869 9011 28921
rect 8881 28805 8933 28857
rect 8959 28805 9011 28857
rect 8881 28741 8933 28793
rect 8959 28741 9011 28793
rect 8881 28677 8933 28729
rect 8959 28677 9011 28729
rect 8881 28612 8933 28664
rect 8959 28612 9011 28664
rect 8881 28547 8933 28599
rect 8959 28547 9011 28599
rect 8881 28482 8933 28534
rect 8959 28482 9011 28534
rect 8881 28417 8933 28469
rect 8959 28417 9011 28469
rect 8881 28352 8933 28404
rect 8959 28352 9011 28404
rect 8881 28287 8933 28339
rect 8959 28287 9011 28339
rect 8881 28222 8933 28274
rect 8959 28222 9011 28274
rect 8881 28157 8933 28209
rect 8959 28157 9011 28209
rect 8881 28092 8933 28144
rect 8959 28092 9011 28144
rect 8881 28027 8933 28079
rect 8959 28027 9011 28079
rect 8881 27962 8933 28014
rect 8959 27962 9011 28014
rect 8881 27897 8933 27949
rect 8959 27897 9011 27949
rect 8881 24973 8933 25025
rect 8959 24973 9011 25025
rect 8881 24909 8933 24961
rect 8959 24909 9011 24961
rect 8881 24845 8933 24897
rect 8959 24845 9011 24897
rect 8881 24781 8933 24833
rect 8959 24781 9011 24833
rect 8881 24717 8933 24769
rect 8959 24717 9011 24769
rect 8881 24653 8933 24705
rect 8959 24653 9011 24705
rect 8881 24589 8933 24641
rect 8959 24589 9011 24641
rect 8881 24525 8933 24577
rect 8959 24525 9011 24577
rect 8881 24461 8933 24513
rect 8959 24461 9011 24513
rect 8881 24397 8933 24449
rect 8959 24397 9011 24449
rect 8881 24333 8933 24385
rect 8959 24333 9011 24385
rect 8881 24269 8933 24321
rect 8959 24269 9011 24321
rect 8881 24205 8933 24257
rect 8959 24205 9011 24257
rect 8881 24141 8933 24193
rect 8959 24141 9011 24193
rect 8881 24077 8933 24129
rect 8959 24077 9011 24129
rect 8881 24012 8933 24064
rect 8959 24012 9011 24064
rect 8881 23947 8933 23999
rect 8959 23947 9011 23999
rect 8881 23882 8933 23934
rect 8959 23882 9011 23934
rect 8881 23817 8933 23869
rect 8959 23817 9011 23869
rect 8881 23752 8933 23804
rect 8959 23752 9011 23804
rect 8881 23687 8933 23739
rect 8959 23687 9011 23739
rect 8881 23622 8933 23674
rect 8959 23622 9011 23674
rect 8881 23557 8933 23609
rect 8959 23557 9011 23609
rect 8881 23492 8933 23544
rect 8959 23492 9011 23544
rect 8881 23427 8933 23479
rect 8959 23427 9011 23479
rect 8881 23362 8933 23414
rect 8959 23362 9011 23414
rect 8881 23297 8933 23349
rect 8959 23297 9011 23349
rect 8881 20373 8933 20425
rect 8959 20373 9011 20425
rect 8881 20309 8933 20361
rect 8959 20309 9011 20361
rect 8881 20245 8933 20297
rect 8959 20245 9011 20297
rect 8881 20181 8933 20233
rect 8959 20181 9011 20233
rect 8881 20117 8933 20169
rect 8959 20117 9011 20169
rect 8881 20053 8933 20105
rect 8959 20053 9011 20105
rect 8881 19989 8933 20041
rect 8959 19989 9011 20041
rect 8881 19925 8933 19977
rect 8959 19925 9011 19977
rect 8881 19861 8933 19913
rect 8959 19861 9011 19913
rect 8881 19797 8933 19849
rect 8959 19797 9011 19849
rect 8881 19733 8933 19785
rect 8959 19733 9011 19785
rect 8881 19669 8933 19721
rect 8959 19669 9011 19721
rect 8881 19605 8933 19657
rect 8959 19605 9011 19657
rect 8881 19541 8933 19593
rect 8959 19541 9011 19593
rect 8881 19477 8933 19529
rect 8959 19477 9011 19529
rect 8881 19412 8933 19464
rect 8959 19412 9011 19464
rect 8881 19347 8933 19399
rect 8959 19347 9011 19399
rect 8881 19282 8933 19334
rect 8959 19282 9011 19334
rect 8881 19217 8933 19269
rect 8959 19217 9011 19269
rect 8881 19152 8933 19204
rect 8959 19152 9011 19204
rect 8881 19087 8933 19139
rect 8959 19087 9011 19139
rect 8881 19022 8933 19074
rect 8959 19022 9011 19074
rect 8881 18957 8933 19009
rect 8959 18957 9011 19009
rect 8881 18892 8933 18944
rect 8959 18892 9011 18944
rect 8881 18827 8933 18879
rect 8959 18827 9011 18879
rect 8881 18762 8933 18814
rect 8959 18762 9011 18814
rect 8881 18697 8933 18749
rect 8959 18697 9011 18749
rect 8881 15773 8933 15825
rect 8959 15773 9011 15825
rect 8881 15709 8933 15761
rect 8959 15709 9011 15761
rect 8881 15645 8933 15697
rect 8959 15645 9011 15697
rect 8881 15581 8933 15633
rect 8959 15581 9011 15633
rect 8881 15517 8933 15569
rect 8959 15517 9011 15569
rect 8881 15453 8933 15505
rect 8959 15453 9011 15505
rect 8881 15389 8933 15441
rect 8959 15389 9011 15441
rect 8881 15325 8933 15377
rect 8959 15325 9011 15377
rect 8881 15261 8933 15313
rect 8959 15261 9011 15313
rect 8881 15197 8933 15249
rect 8959 15197 9011 15249
rect 8881 15133 8933 15185
rect 8959 15133 9011 15185
rect 8881 15069 8933 15121
rect 8959 15069 9011 15121
rect 8881 15005 8933 15057
rect 8959 15005 9011 15057
rect 8881 14941 8933 14993
rect 8959 14941 9011 14993
rect 8881 14877 8933 14929
rect 8959 14877 9011 14929
rect 8881 14812 8933 14864
rect 8959 14812 9011 14864
rect 8881 14747 8933 14799
rect 8959 14747 9011 14799
rect 8881 14682 8933 14734
rect 8959 14682 9011 14734
rect 8881 14617 8933 14669
rect 8959 14617 9011 14669
rect 8881 14552 8933 14604
rect 8959 14552 9011 14604
rect 8881 14487 8933 14539
rect 8959 14487 9011 14539
rect 8881 14422 8933 14474
rect 8959 14422 9011 14474
rect 8881 14357 8933 14409
rect 8959 14357 9011 14409
rect 8881 14292 8933 14344
rect 8959 14292 9011 14344
rect 8881 14227 8933 14279
rect 8959 14227 9011 14279
rect 8881 14162 8933 14214
rect 8959 14162 9011 14214
rect 8881 14097 8933 14149
rect 8959 14097 9011 14149
rect 8881 11173 8933 11225
rect 8959 11173 9011 11225
rect 8881 11109 8933 11161
rect 8959 11109 9011 11161
rect 8881 11045 8933 11097
rect 8959 11045 9011 11097
rect 8881 10981 8933 11033
rect 8959 10981 9011 11033
rect 8881 10917 8933 10969
rect 8959 10917 9011 10969
rect 8881 10853 8933 10905
rect 8959 10853 9011 10905
rect 8881 10789 8933 10841
rect 8959 10789 9011 10841
rect 8881 10725 8933 10777
rect 8959 10725 9011 10777
rect 8881 10661 8933 10713
rect 8959 10661 9011 10713
rect 8881 10597 8933 10649
rect 8959 10597 9011 10649
rect 8881 10533 8933 10585
rect 8959 10533 9011 10585
rect 8881 10469 8933 10521
rect 8959 10469 9011 10521
rect 8881 10405 8933 10457
rect 8959 10405 9011 10457
rect 8881 10341 8933 10393
rect 8959 10341 9011 10393
rect 8881 10277 8933 10329
rect 8959 10277 9011 10329
rect 8881 10212 8933 10264
rect 8959 10212 9011 10264
rect 8881 10147 8933 10199
rect 8959 10147 9011 10199
rect 8881 10082 8933 10134
rect 8959 10082 9011 10134
rect 8881 10017 8933 10069
rect 8959 10017 9011 10069
rect 8881 9952 8933 10004
rect 8959 9952 9011 10004
rect 8881 9887 8933 9939
rect 8959 9887 9011 9939
rect 8881 9822 8933 9874
rect 8959 9822 9011 9874
rect 8881 9757 8933 9809
rect 8959 9757 9011 9809
rect 8881 9692 8933 9744
rect 8959 9692 9011 9744
rect 8881 9627 8933 9679
rect 8959 9627 9011 9679
rect 8881 9562 8933 9614
rect 8959 9562 9011 9614
rect 8881 9497 8933 9549
rect 8959 9497 9011 9549
rect 9312 36238 9317 36290
rect 9317 36238 9364 36290
rect 9380 36238 9432 36290
rect 9448 36238 9495 36290
rect 9495 36238 9500 36290
rect 9312 36174 9317 36226
rect 9317 36174 9364 36226
rect 9380 36174 9432 36226
rect 9448 36174 9495 36226
rect 9495 36174 9500 36226
rect 9312 36110 9317 36162
rect 9317 36110 9364 36162
rect 9380 36110 9432 36162
rect 9448 36110 9495 36162
rect 9495 36110 9500 36162
rect 9312 36046 9317 36098
rect 9317 36046 9364 36098
rect 9380 36046 9432 36098
rect 9448 36046 9495 36098
rect 9495 36046 9500 36098
rect 9312 35982 9317 36034
rect 9317 35982 9364 36034
rect 9380 35982 9432 36034
rect 9448 35982 9495 36034
rect 9495 35982 9500 36034
rect 9312 35918 9317 35970
rect 9317 35918 9364 35970
rect 9380 35918 9432 35970
rect 9448 35918 9495 35970
rect 9495 35918 9500 35970
rect 9312 35854 9317 35906
rect 9317 35854 9364 35906
rect 9380 35854 9432 35906
rect 9448 35854 9495 35906
rect 9495 35854 9500 35906
rect 9312 35790 9317 35842
rect 9317 35790 9364 35842
rect 9380 35790 9432 35842
rect 9448 35790 9495 35842
rect 9495 35790 9500 35842
rect 9312 35726 9317 35778
rect 9317 35726 9364 35778
rect 9380 35726 9432 35778
rect 9448 35726 9495 35778
rect 9495 35726 9500 35778
rect 9312 35662 9317 35714
rect 9317 35662 9364 35714
rect 9380 35662 9432 35714
rect 9448 35662 9495 35714
rect 9495 35662 9500 35714
rect 9312 35598 9317 35650
rect 9317 35598 9364 35650
rect 9380 35598 9432 35650
rect 9448 35598 9495 35650
rect 9495 35598 9500 35650
rect 9312 35534 9317 35586
rect 9317 35534 9364 35586
rect 9380 35534 9432 35586
rect 9448 35534 9495 35586
rect 9495 35534 9500 35586
rect 9312 35470 9317 35522
rect 9317 35470 9364 35522
rect 9380 35470 9432 35522
rect 9448 35470 9495 35522
rect 9495 35470 9500 35522
rect 9312 35406 9317 35458
rect 9317 35406 9364 35458
rect 9380 35406 9432 35458
rect 9448 35406 9495 35458
rect 9495 35406 9500 35458
rect 9312 35342 9317 35394
rect 9317 35342 9364 35394
rect 9380 35342 9432 35394
rect 9448 35342 9495 35394
rect 9495 35342 9500 35394
rect 9312 35277 9317 35329
rect 9317 35277 9364 35329
rect 9380 35277 9432 35329
rect 9448 35277 9495 35329
rect 9495 35277 9500 35329
rect 9312 35212 9317 35264
rect 9317 35212 9364 35264
rect 9380 35212 9432 35264
rect 9448 35212 9495 35264
rect 9495 35212 9500 35264
rect 9312 35147 9317 35199
rect 9317 35147 9364 35199
rect 9380 35147 9432 35199
rect 9448 35147 9495 35199
rect 9495 35147 9500 35199
rect 9312 35082 9317 35134
rect 9317 35082 9364 35134
rect 9380 35082 9432 35134
rect 9448 35082 9495 35134
rect 9495 35082 9500 35134
rect 9312 35017 9317 35069
rect 9317 35017 9364 35069
rect 9380 35017 9432 35069
rect 9448 35017 9495 35069
rect 9495 35017 9500 35069
rect 9312 34952 9317 35004
rect 9317 34952 9364 35004
rect 9380 34952 9432 35004
rect 9448 34952 9495 35004
rect 9495 34952 9500 35004
rect 9312 34887 9317 34939
rect 9317 34887 9364 34939
rect 9380 34887 9432 34939
rect 9448 34887 9495 34939
rect 9495 34887 9500 34939
rect 9312 34822 9317 34874
rect 9317 34822 9364 34874
rect 9380 34822 9432 34874
rect 9448 34822 9495 34874
rect 9495 34822 9500 34874
rect 9312 34757 9317 34809
rect 9317 34757 9364 34809
rect 9380 34757 9432 34809
rect 9448 34757 9495 34809
rect 9495 34757 9500 34809
rect 9312 34692 9317 34744
rect 9317 34692 9364 34744
rect 9380 34692 9432 34744
rect 9448 34692 9495 34744
rect 9495 34692 9500 34744
rect 9312 34627 9317 34679
rect 9317 34627 9364 34679
rect 9380 34627 9432 34679
rect 9448 34627 9495 34679
rect 9495 34627 9500 34679
rect 9312 34562 9317 34614
rect 9317 34562 9364 34614
rect 9380 34562 9432 34614
rect 9448 34562 9495 34614
rect 9495 34562 9500 34614
rect 9312 31638 9317 31690
rect 9317 31638 9364 31690
rect 9380 31638 9432 31690
rect 9448 31638 9495 31690
rect 9495 31638 9500 31690
rect 9312 31574 9317 31626
rect 9317 31574 9364 31626
rect 9380 31574 9432 31626
rect 9448 31574 9495 31626
rect 9495 31574 9500 31626
rect 9312 31510 9317 31562
rect 9317 31510 9364 31562
rect 9380 31510 9432 31562
rect 9448 31510 9495 31562
rect 9495 31510 9500 31562
rect 9312 31446 9317 31498
rect 9317 31446 9364 31498
rect 9380 31446 9432 31498
rect 9448 31446 9495 31498
rect 9495 31446 9500 31498
rect 9312 31382 9317 31434
rect 9317 31382 9364 31434
rect 9380 31382 9432 31434
rect 9448 31382 9495 31434
rect 9495 31382 9500 31434
rect 9312 31318 9317 31370
rect 9317 31318 9364 31370
rect 9380 31318 9432 31370
rect 9448 31318 9495 31370
rect 9495 31318 9500 31370
rect 9312 31254 9317 31306
rect 9317 31254 9364 31306
rect 9380 31254 9432 31306
rect 9448 31254 9495 31306
rect 9495 31254 9500 31306
rect 9312 31190 9317 31242
rect 9317 31190 9364 31242
rect 9380 31190 9432 31242
rect 9448 31190 9495 31242
rect 9495 31190 9500 31242
rect 9312 31126 9317 31178
rect 9317 31126 9364 31178
rect 9380 31126 9432 31178
rect 9448 31126 9495 31178
rect 9495 31126 9500 31178
rect 9312 31062 9317 31114
rect 9317 31062 9364 31114
rect 9380 31062 9432 31114
rect 9448 31062 9495 31114
rect 9495 31062 9500 31114
rect 9312 30998 9317 31050
rect 9317 30998 9364 31050
rect 9380 30998 9432 31050
rect 9448 30998 9495 31050
rect 9495 30998 9500 31050
rect 9312 30934 9317 30986
rect 9317 30934 9364 30986
rect 9380 30934 9432 30986
rect 9448 30934 9495 30986
rect 9495 30934 9500 30986
rect 9312 30870 9317 30922
rect 9317 30870 9364 30922
rect 9380 30870 9432 30922
rect 9448 30870 9495 30922
rect 9495 30870 9500 30922
rect 9312 30806 9317 30858
rect 9317 30806 9364 30858
rect 9380 30806 9432 30858
rect 9448 30806 9495 30858
rect 9495 30806 9500 30858
rect 9312 30742 9317 30794
rect 9317 30742 9364 30794
rect 9380 30742 9432 30794
rect 9448 30742 9495 30794
rect 9495 30742 9500 30794
rect 9312 30677 9317 30729
rect 9317 30677 9364 30729
rect 9380 30677 9432 30729
rect 9448 30677 9495 30729
rect 9495 30677 9500 30729
rect 9312 30612 9317 30664
rect 9317 30612 9364 30664
rect 9380 30612 9432 30664
rect 9448 30612 9495 30664
rect 9495 30612 9500 30664
rect 9312 30547 9317 30599
rect 9317 30547 9364 30599
rect 9380 30547 9432 30599
rect 9448 30547 9495 30599
rect 9495 30547 9500 30599
rect 9312 30482 9317 30534
rect 9317 30482 9364 30534
rect 9380 30482 9432 30534
rect 9448 30482 9495 30534
rect 9495 30482 9500 30534
rect 9312 30417 9317 30469
rect 9317 30417 9364 30469
rect 9380 30417 9432 30469
rect 9448 30417 9495 30469
rect 9495 30417 9500 30469
rect 9312 30352 9317 30404
rect 9317 30352 9364 30404
rect 9380 30352 9432 30404
rect 9448 30352 9495 30404
rect 9495 30352 9500 30404
rect 9312 30287 9317 30339
rect 9317 30287 9364 30339
rect 9380 30287 9432 30339
rect 9448 30287 9495 30339
rect 9495 30287 9500 30339
rect 9312 30222 9317 30274
rect 9317 30222 9364 30274
rect 9380 30222 9432 30274
rect 9448 30222 9495 30274
rect 9495 30222 9500 30274
rect 9312 30157 9317 30209
rect 9317 30157 9364 30209
rect 9380 30157 9432 30209
rect 9448 30157 9495 30209
rect 9495 30157 9500 30209
rect 9312 30092 9317 30144
rect 9317 30092 9364 30144
rect 9380 30092 9432 30144
rect 9448 30092 9495 30144
rect 9495 30092 9500 30144
rect 9312 30027 9317 30079
rect 9317 30027 9364 30079
rect 9380 30027 9432 30079
rect 9448 30027 9495 30079
rect 9495 30027 9500 30079
rect 9312 29962 9317 30014
rect 9317 29962 9364 30014
rect 9380 29962 9432 30014
rect 9448 29962 9495 30014
rect 9495 29962 9500 30014
rect 9312 27038 9317 27090
rect 9317 27038 9364 27090
rect 9380 27038 9432 27090
rect 9448 27038 9495 27090
rect 9495 27038 9500 27090
rect 9312 26974 9317 27026
rect 9317 26974 9364 27026
rect 9380 26974 9432 27026
rect 9448 26974 9495 27026
rect 9495 26974 9500 27026
rect 9312 26910 9317 26962
rect 9317 26910 9364 26962
rect 9380 26910 9432 26962
rect 9448 26910 9495 26962
rect 9495 26910 9500 26962
rect 9312 26846 9317 26898
rect 9317 26846 9364 26898
rect 9380 26846 9432 26898
rect 9448 26846 9495 26898
rect 9495 26846 9500 26898
rect 9312 26782 9317 26834
rect 9317 26782 9364 26834
rect 9380 26782 9432 26834
rect 9448 26782 9495 26834
rect 9495 26782 9500 26834
rect 9312 26718 9317 26770
rect 9317 26718 9364 26770
rect 9380 26718 9432 26770
rect 9448 26718 9495 26770
rect 9495 26718 9500 26770
rect 9312 26654 9317 26706
rect 9317 26654 9364 26706
rect 9380 26654 9432 26706
rect 9448 26654 9495 26706
rect 9495 26654 9500 26706
rect 9312 26590 9317 26642
rect 9317 26590 9364 26642
rect 9380 26590 9432 26642
rect 9448 26590 9495 26642
rect 9495 26590 9500 26642
rect 9312 26526 9317 26578
rect 9317 26526 9364 26578
rect 9380 26526 9432 26578
rect 9448 26526 9495 26578
rect 9495 26526 9500 26578
rect 9312 26462 9317 26514
rect 9317 26462 9364 26514
rect 9380 26462 9432 26514
rect 9448 26462 9495 26514
rect 9495 26462 9500 26514
rect 9312 26398 9317 26450
rect 9317 26398 9364 26450
rect 9380 26398 9432 26450
rect 9448 26398 9495 26450
rect 9495 26398 9500 26450
rect 9312 26334 9317 26386
rect 9317 26334 9364 26386
rect 9380 26334 9432 26386
rect 9448 26334 9495 26386
rect 9495 26334 9500 26386
rect 9312 26270 9317 26322
rect 9317 26270 9364 26322
rect 9380 26270 9432 26322
rect 9448 26270 9495 26322
rect 9495 26270 9500 26322
rect 9312 26206 9317 26258
rect 9317 26206 9364 26258
rect 9380 26206 9432 26258
rect 9448 26206 9495 26258
rect 9495 26206 9500 26258
rect 9312 26142 9317 26194
rect 9317 26142 9364 26194
rect 9380 26142 9432 26194
rect 9448 26142 9495 26194
rect 9495 26142 9500 26194
rect 9312 26077 9317 26129
rect 9317 26077 9364 26129
rect 9380 26077 9432 26129
rect 9448 26077 9495 26129
rect 9495 26077 9500 26129
rect 9312 26012 9317 26064
rect 9317 26012 9364 26064
rect 9380 26012 9432 26064
rect 9448 26012 9495 26064
rect 9495 26012 9500 26064
rect 9312 25947 9317 25999
rect 9317 25947 9364 25999
rect 9380 25947 9432 25999
rect 9448 25947 9495 25999
rect 9495 25947 9500 25999
rect 9312 25882 9317 25934
rect 9317 25882 9364 25934
rect 9380 25882 9432 25934
rect 9448 25882 9495 25934
rect 9495 25882 9500 25934
rect 9312 25817 9317 25869
rect 9317 25817 9364 25869
rect 9380 25817 9432 25869
rect 9448 25817 9495 25869
rect 9495 25817 9500 25869
rect 9312 25752 9317 25804
rect 9317 25752 9364 25804
rect 9380 25752 9432 25804
rect 9448 25752 9495 25804
rect 9495 25752 9500 25804
rect 9312 25687 9317 25739
rect 9317 25687 9364 25739
rect 9380 25687 9432 25739
rect 9448 25687 9495 25739
rect 9495 25687 9500 25739
rect 9312 25622 9317 25674
rect 9317 25622 9364 25674
rect 9380 25622 9432 25674
rect 9448 25622 9495 25674
rect 9495 25622 9500 25674
rect 9312 25557 9317 25609
rect 9317 25557 9364 25609
rect 9380 25557 9432 25609
rect 9448 25557 9495 25609
rect 9495 25557 9500 25609
rect 9312 25492 9317 25544
rect 9317 25492 9364 25544
rect 9380 25492 9432 25544
rect 9448 25492 9495 25544
rect 9495 25492 9500 25544
rect 9312 25427 9317 25479
rect 9317 25427 9364 25479
rect 9380 25427 9432 25479
rect 9448 25427 9495 25479
rect 9495 25427 9500 25479
rect 9312 25362 9317 25414
rect 9317 25362 9364 25414
rect 9380 25362 9432 25414
rect 9448 25362 9495 25414
rect 9495 25362 9500 25414
rect 9312 22438 9317 22490
rect 9317 22438 9364 22490
rect 9380 22438 9432 22490
rect 9448 22438 9495 22490
rect 9495 22438 9500 22490
rect 9312 22374 9317 22426
rect 9317 22374 9364 22426
rect 9380 22374 9432 22426
rect 9448 22374 9495 22426
rect 9495 22374 9500 22426
rect 9312 22310 9317 22362
rect 9317 22310 9364 22362
rect 9380 22310 9432 22362
rect 9448 22310 9495 22362
rect 9495 22310 9500 22362
rect 9312 22246 9317 22298
rect 9317 22246 9364 22298
rect 9380 22246 9432 22298
rect 9448 22246 9495 22298
rect 9495 22246 9500 22298
rect 9312 22182 9317 22234
rect 9317 22182 9364 22234
rect 9380 22182 9432 22234
rect 9448 22182 9495 22234
rect 9495 22182 9500 22234
rect 9312 22118 9317 22170
rect 9317 22118 9364 22170
rect 9380 22118 9432 22170
rect 9448 22118 9495 22170
rect 9495 22118 9500 22170
rect 9312 22054 9317 22106
rect 9317 22054 9364 22106
rect 9380 22054 9432 22106
rect 9448 22054 9495 22106
rect 9495 22054 9500 22106
rect 9312 21990 9317 22042
rect 9317 21990 9364 22042
rect 9380 21990 9432 22042
rect 9448 21990 9495 22042
rect 9495 21990 9500 22042
rect 9312 21926 9317 21978
rect 9317 21926 9364 21978
rect 9380 21926 9432 21978
rect 9448 21926 9495 21978
rect 9495 21926 9500 21978
rect 9312 21862 9317 21914
rect 9317 21862 9364 21914
rect 9380 21862 9432 21914
rect 9448 21862 9495 21914
rect 9495 21862 9500 21914
rect 9312 21798 9317 21850
rect 9317 21798 9364 21850
rect 9380 21798 9432 21850
rect 9448 21798 9495 21850
rect 9495 21798 9500 21850
rect 9312 21734 9317 21786
rect 9317 21734 9364 21786
rect 9380 21734 9432 21786
rect 9448 21734 9495 21786
rect 9495 21734 9500 21786
rect 9312 21670 9317 21722
rect 9317 21670 9364 21722
rect 9380 21670 9432 21722
rect 9448 21670 9495 21722
rect 9495 21670 9500 21722
rect 9312 21606 9317 21658
rect 9317 21606 9364 21658
rect 9380 21606 9432 21658
rect 9448 21606 9495 21658
rect 9495 21606 9500 21658
rect 9312 21542 9317 21594
rect 9317 21542 9364 21594
rect 9380 21542 9432 21594
rect 9448 21542 9495 21594
rect 9495 21542 9500 21594
rect 9312 21477 9317 21529
rect 9317 21477 9364 21529
rect 9380 21477 9432 21529
rect 9448 21477 9495 21529
rect 9495 21477 9500 21529
rect 9312 21412 9317 21464
rect 9317 21412 9364 21464
rect 9380 21412 9432 21464
rect 9448 21412 9495 21464
rect 9495 21412 9500 21464
rect 9312 21347 9317 21399
rect 9317 21347 9364 21399
rect 9380 21347 9432 21399
rect 9448 21347 9495 21399
rect 9495 21347 9500 21399
rect 9312 21282 9317 21334
rect 9317 21282 9364 21334
rect 9380 21282 9432 21334
rect 9448 21282 9495 21334
rect 9495 21282 9500 21334
rect 9312 21217 9317 21269
rect 9317 21217 9364 21269
rect 9380 21217 9432 21269
rect 9448 21217 9495 21269
rect 9495 21217 9500 21269
rect 9312 21152 9317 21204
rect 9317 21152 9364 21204
rect 9380 21152 9432 21204
rect 9448 21152 9495 21204
rect 9495 21152 9500 21204
rect 9312 21087 9317 21139
rect 9317 21087 9364 21139
rect 9380 21087 9432 21139
rect 9448 21087 9495 21139
rect 9495 21087 9500 21139
rect 9312 21022 9317 21074
rect 9317 21022 9364 21074
rect 9380 21022 9432 21074
rect 9448 21022 9495 21074
rect 9495 21022 9500 21074
rect 9312 20957 9317 21009
rect 9317 20957 9364 21009
rect 9380 20957 9432 21009
rect 9448 20957 9495 21009
rect 9495 20957 9500 21009
rect 9312 20892 9317 20944
rect 9317 20892 9364 20944
rect 9380 20892 9432 20944
rect 9448 20892 9495 20944
rect 9495 20892 9500 20944
rect 9312 20827 9317 20879
rect 9317 20827 9364 20879
rect 9380 20827 9432 20879
rect 9448 20827 9495 20879
rect 9495 20827 9500 20879
rect 9312 20762 9317 20814
rect 9317 20762 9364 20814
rect 9380 20762 9432 20814
rect 9448 20762 9495 20814
rect 9495 20762 9500 20814
rect 9312 17838 9317 17890
rect 9317 17838 9364 17890
rect 9380 17838 9432 17890
rect 9448 17838 9495 17890
rect 9495 17838 9500 17890
rect 9312 17774 9317 17826
rect 9317 17774 9364 17826
rect 9380 17774 9432 17826
rect 9448 17774 9495 17826
rect 9495 17774 9500 17826
rect 9312 17710 9317 17762
rect 9317 17710 9364 17762
rect 9380 17710 9432 17762
rect 9448 17710 9495 17762
rect 9495 17710 9500 17762
rect 9312 17646 9317 17698
rect 9317 17646 9364 17698
rect 9380 17646 9432 17698
rect 9448 17646 9495 17698
rect 9495 17646 9500 17698
rect 9312 17582 9317 17634
rect 9317 17582 9364 17634
rect 9380 17582 9432 17634
rect 9448 17582 9495 17634
rect 9495 17582 9500 17634
rect 9312 17518 9317 17570
rect 9317 17518 9364 17570
rect 9380 17518 9432 17570
rect 9448 17518 9495 17570
rect 9495 17518 9500 17570
rect 9312 17454 9317 17506
rect 9317 17454 9364 17506
rect 9380 17454 9432 17506
rect 9448 17454 9495 17506
rect 9495 17454 9500 17506
rect 9312 17390 9317 17442
rect 9317 17390 9364 17442
rect 9380 17390 9432 17442
rect 9448 17390 9495 17442
rect 9495 17390 9500 17442
rect 9312 17326 9317 17378
rect 9317 17326 9364 17378
rect 9380 17326 9432 17378
rect 9448 17326 9495 17378
rect 9495 17326 9500 17378
rect 9312 17262 9317 17314
rect 9317 17262 9364 17314
rect 9380 17262 9432 17314
rect 9448 17262 9495 17314
rect 9495 17262 9500 17314
rect 9312 17198 9317 17250
rect 9317 17198 9364 17250
rect 9380 17198 9432 17250
rect 9448 17198 9495 17250
rect 9495 17198 9500 17250
rect 9312 17134 9317 17186
rect 9317 17134 9364 17186
rect 9380 17134 9432 17186
rect 9448 17134 9495 17186
rect 9495 17134 9500 17186
rect 9312 17070 9317 17122
rect 9317 17070 9364 17122
rect 9380 17070 9432 17122
rect 9448 17070 9495 17122
rect 9495 17070 9500 17122
rect 9312 17006 9317 17058
rect 9317 17006 9364 17058
rect 9380 17006 9432 17058
rect 9448 17006 9495 17058
rect 9495 17006 9500 17058
rect 9312 16942 9317 16994
rect 9317 16942 9364 16994
rect 9380 16942 9432 16994
rect 9448 16942 9495 16994
rect 9495 16942 9500 16994
rect 9312 16877 9317 16929
rect 9317 16877 9364 16929
rect 9380 16877 9432 16929
rect 9448 16877 9495 16929
rect 9495 16877 9500 16929
rect 9312 16812 9317 16864
rect 9317 16812 9364 16864
rect 9380 16812 9432 16864
rect 9448 16812 9495 16864
rect 9495 16812 9500 16864
rect 9312 16747 9317 16799
rect 9317 16747 9364 16799
rect 9380 16747 9432 16799
rect 9448 16747 9495 16799
rect 9495 16747 9500 16799
rect 9312 16682 9317 16734
rect 9317 16682 9364 16734
rect 9380 16682 9432 16734
rect 9448 16682 9495 16734
rect 9495 16682 9500 16734
rect 9312 16617 9317 16669
rect 9317 16617 9364 16669
rect 9380 16617 9432 16669
rect 9448 16617 9495 16669
rect 9495 16617 9500 16669
rect 9312 16552 9317 16604
rect 9317 16552 9364 16604
rect 9380 16552 9432 16604
rect 9448 16552 9495 16604
rect 9495 16552 9500 16604
rect 9312 16487 9317 16539
rect 9317 16487 9364 16539
rect 9380 16487 9432 16539
rect 9448 16487 9495 16539
rect 9495 16487 9500 16539
rect 9312 16422 9317 16474
rect 9317 16422 9364 16474
rect 9380 16422 9432 16474
rect 9448 16422 9495 16474
rect 9495 16422 9500 16474
rect 9312 16357 9317 16409
rect 9317 16357 9364 16409
rect 9380 16357 9432 16409
rect 9448 16357 9495 16409
rect 9495 16357 9500 16409
rect 9312 16292 9317 16344
rect 9317 16292 9364 16344
rect 9380 16292 9432 16344
rect 9448 16292 9495 16344
rect 9495 16292 9500 16344
rect 9312 16227 9317 16279
rect 9317 16227 9364 16279
rect 9380 16227 9432 16279
rect 9448 16227 9495 16279
rect 9495 16227 9500 16279
rect 9312 16162 9317 16214
rect 9317 16162 9364 16214
rect 9380 16162 9432 16214
rect 9448 16162 9495 16214
rect 9495 16162 9500 16214
rect 9312 13238 9317 13290
rect 9317 13238 9364 13290
rect 9380 13238 9432 13290
rect 9448 13238 9495 13290
rect 9495 13238 9500 13290
rect 9312 13174 9317 13226
rect 9317 13174 9364 13226
rect 9380 13174 9432 13226
rect 9448 13174 9495 13226
rect 9495 13174 9500 13226
rect 9312 13110 9317 13162
rect 9317 13110 9364 13162
rect 9380 13110 9432 13162
rect 9448 13110 9495 13162
rect 9495 13110 9500 13162
rect 9312 13046 9317 13098
rect 9317 13046 9364 13098
rect 9380 13046 9432 13098
rect 9448 13046 9495 13098
rect 9495 13046 9500 13098
rect 9312 12982 9317 13034
rect 9317 12982 9364 13034
rect 9380 12982 9432 13034
rect 9448 12982 9495 13034
rect 9495 12982 9500 13034
rect 9312 12918 9317 12970
rect 9317 12918 9364 12970
rect 9380 12918 9432 12970
rect 9448 12918 9495 12970
rect 9495 12918 9500 12970
rect 9312 12854 9317 12906
rect 9317 12854 9364 12906
rect 9380 12854 9432 12906
rect 9448 12854 9495 12906
rect 9495 12854 9500 12906
rect 9312 12790 9317 12842
rect 9317 12790 9364 12842
rect 9380 12790 9432 12842
rect 9448 12790 9495 12842
rect 9495 12790 9500 12842
rect 9312 12726 9317 12778
rect 9317 12726 9364 12778
rect 9380 12726 9432 12778
rect 9448 12726 9495 12778
rect 9495 12726 9500 12778
rect 9312 12662 9317 12714
rect 9317 12662 9364 12714
rect 9380 12662 9432 12714
rect 9448 12662 9495 12714
rect 9495 12662 9500 12714
rect 9312 12598 9317 12650
rect 9317 12598 9364 12650
rect 9380 12598 9432 12650
rect 9448 12598 9495 12650
rect 9495 12598 9500 12650
rect 9312 12534 9317 12586
rect 9317 12534 9364 12586
rect 9380 12534 9432 12586
rect 9448 12534 9495 12586
rect 9495 12534 9500 12586
rect 9312 12470 9317 12522
rect 9317 12470 9364 12522
rect 9380 12470 9432 12522
rect 9448 12470 9495 12522
rect 9495 12470 9500 12522
rect 9312 12406 9317 12458
rect 9317 12406 9364 12458
rect 9380 12406 9432 12458
rect 9448 12406 9495 12458
rect 9495 12406 9500 12458
rect 9312 12342 9317 12394
rect 9317 12342 9364 12394
rect 9380 12342 9432 12394
rect 9448 12342 9495 12394
rect 9495 12342 9500 12394
rect 9312 12277 9317 12329
rect 9317 12277 9364 12329
rect 9380 12277 9432 12329
rect 9448 12277 9495 12329
rect 9495 12277 9500 12329
rect 9312 12212 9317 12264
rect 9317 12212 9364 12264
rect 9380 12212 9432 12264
rect 9448 12212 9495 12264
rect 9495 12212 9500 12264
rect 9312 12147 9317 12199
rect 9317 12147 9364 12199
rect 9380 12147 9432 12199
rect 9448 12147 9495 12199
rect 9495 12147 9500 12199
rect 9312 12082 9317 12134
rect 9317 12082 9364 12134
rect 9380 12082 9432 12134
rect 9448 12082 9495 12134
rect 9495 12082 9500 12134
rect 9312 12017 9317 12069
rect 9317 12017 9364 12069
rect 9380 12017 9432 12069
rect 9448 12017 9495 12069
rect 9495 12017 9500 12069
rect 9312 11952 9317 12004
rect 9317 11952 9364 12004
rect 9380 11952 9432 12004
rect 9448 11952 9495 12004
rect 9495 11952 9500 12004
rect 9312 11887 9317 11939
rect 9317 11887 9364 11939
rect 9380 11887 9432 11939
rect 9448 11887 9495 11939
rect 9495 11887 9500 11939
rect 9312 11822 9317 11874
rect 9317 11822 9364 11874
rect 9380 11822 9432 11874
rect 9448 11822 9495 11874
rect 9495 11822 9500 11874
rect 9312 11757 9317 11809
rect 9317 11757 9364 11809
rect 9380 11757 9432 11809
rect 9448 11757 9495 11809
rect 9495 11757 9500 11809
rect 9312 11692 9317 11744
rect 9317 11692 9364 11744
rect 9380 11692 9432 11744
rect 9448 11692 9495 11744
rect 9495 11692 9500 11744
rect 9312 11627 9317 11679
rect 9317 11627 9364 11679
rect 9380 11627 9432 11679
rect 9448 11627 9495 11679
rect 9495 11627 9500 11679
rect 9312 11562 9317 11614
rect 9317 11562 9364 11614
rect 9380 11562 9432 11614
rect 9448 11562 9495 11614
rect 9495 11562 9500 11614
rect 9801 37945 9853 37997
rect 9879 37945 9931 37997
rect 9801 37877 9853 37929
rect 9879 37877 9931 37929
rect 9801 37809 9853 37861
rect 9879 37809 9931 37861
rect 9801 37741 9853 37793
rect 9879 37741 9931 37793
rect 9801 37673 9853 37725
rect 9879 37673 9931 37725
rect 9801 37605 9853 37657
rect 9879 37605 9931 37657
rect 9801 37537 9853 37589
rect 9879 37537 9931 37589
rect 9801 37469 9853 37521
rect 9879 37469 9931 37521
rect 9801 37401 9853 37453
rect 9879 37401 9931 37453
rect 9801 37333 9853 37385
rect 9879 37333 9931 37385
rect 9801 37266 9853 37318
rect 9879 37266 9931 37318
rect 9801 37199 9853 37251
rect 9879 37199 9931 37251
rect 9801 37132 9853 37184
rect 9879 37132 9931 37184
rect 9801 37065 9853 37117
rect 9879 37065 9931 37117
rect 9801 34173 9853 34225
rect 9879 34173 9931 34225
rect 9801 34109 9853 34161
rect 9879 34109 9931 34161
rect 9801 34045 9853 34097
rect 9879 34045 9931 34097
rect 9801 33981 9853 34033
rect 9879 33981 9931 34033
rect 9801 33917 9853 33969
rect 9879 33917 9931 33969
rect 9801 33853 9853 33905
rect 9879 33853 9931 33905
rect 9801 33789 9853 33841
rect 9879 33789 9931 33841
rect 9801 33725 9853 33777
rect 9879 33725 9931 33777
rect 9801 33661 9853 33713
rect 9879 33661 9931 33713
rect 9801 33597 9853 33649
rect 9879 33597 9931 33649
rect 9801 33533 9853 33585
rect 9879 33533 9931 33585
rect 9801 33469 9853 33521
rect 9879 33469 9931 33521
rect 9801 33405 9853 33457
rect 9879 33405 9931 33457
rect 9801 33341 9853 33393
rect 9879 33341 9931 33393
rect 9801 33277 9853 33329
rect 9879 33277 9931 33329
rect 9801 33212 9853 33264
rect 9879 33212 9931 33264
rect 9801 33147 9853 33199
rect 9879 33147 9931 33199
rect 9801 33082 9853 33134
rect 9879 33082 9931 33134
rect 9801 33017 9853 33069
rect 9879 33017 9931 33069
rect 9801 32952 9853 33004
rect 9879 32952 9931 33004
rect 9801 32887 9853 32939
rect 9879 32887 9931 32939
rect 9801 32822 9853 32874
rect 9879 32822 9931 32874
rect 9801 32757 9853 32809
rect 9879 32757 9931 32809
rect 9801 32692 9853 32744
rect 9879 32692 9931 32744
rect 9801 32627 9853 32679
rect 9879 32627 9931 32679
rect 9801 32562 9853 32614
rect 9879 32562 9931 32614
rect 9801 32497 9853 32549
rect 9879 32497 9931 32549
rect 9801 29573 9853 29625
rect 9879 29573 9931 29625
rect 9801 29509 9853 29561
rect 9879 29509 9931 29561
rect 9801 29445 9853 29497
rect 9879 29445 9931 29497
rect 9801 29381 9853 29433
rect 9879 29381 9931 29433
rect 9801 29317 9853 29369
rect 9879 29317 9931 29369
rect 9801 29253 9853 29305
rect 9879 29253 9931 29305
rect 9801 29189 9853 29241
rect 9879 29189 9931 29241
rect 9801 29125 9853 29177
rect 9879 29125 9931 29177
rect 9801 29061 9853 29113
rect 9879 29061 9931 29113
rect 9801 28997 9853 29049
rect 9879 28997 9931 29049
rect 9801 28933 9853 28985
rect 9879 28933 9931 28985
rect 9801 28869 9853 28921
rect 9879 28869 9931 28921
rect 9801 28805 9853 28857
rect 9879 28805 9931 28857
rect 9801 28741 9853 28793
rect 9879 28741 9931 28793
rect 9801 28677 9853 28729
rect 9879 28677 9931 28729
rect 9801 28612 9853 28664
rect 9879 28612 9931 28664
rect 9801 28547 9853 28599
rect 9879 28547 9931 28599
rect 9801 28482 9853 28534
rect 9879 28482 9931 28534
rect 9801 28417 9853 28469
rect 9879 28417 9931 28469
rect 9801 28352 9853 28404
rect 9879 28352 9931 28404
rect 9801 28287 9853 28339
rect 9879 28287 9931 28339
rect 9801 28222 9853 28274
rect 9879 28222 9931 28274
rect 9801 28157 9853 28209
rect 9879 28157 9931 28209
rect 9801 28092 9853 28144
rect 9879 28092 9931 28144
rect 9801 28027 9853 28079
rect 9879 28027 9931 28079
rect 9801 27962 9853 28014
rect 9879 27962 9931 28014
rect 9801 27897 9853 27949
rect 9879 27897 9931 27949
rect 9801 24973 9853 25025
rect 9879 24973 9931 25025
rect 9801 24909 9853 24961
rect 9879 24909 9931 24961
rect 9801 24845 9853 24897
rect 9879 24845 9931 24897
rect 9801 24781 9853 24833
rect 9879 24781 9931 24833
rect 9801 24717 9853 24769
rect 9879 24717 9931 24769
rect 9801 24653 9853 24705
rect 9879 24653 9931 24705
rect 9801 24589 9853 24641
rect 9879 24589 9931 24641
rect 9801 24525 9853 24577
rect 9879 24525 9931 24577
rect 9801 24461 9853 24513
rect 9879 24461 9931 24513
rect 9801 24397 9853 24449
rect 9879 24397 9931 24449
rect 9801 24333 9853 24385
rect 9879 24333 9931 24385
rect 9801 24269 9853 24321
rect 9879 24269 9931 24321
rect 9801 24205 9853 24257
rect 9879 24205 9931 24257
rect 9801 24141 9853 24193
rect 9879 24141 9931 24193
rect 9801 24077 9853 24129
rect 9879 24077 9931 24129
rect 9801 24012 9853 24064
rect 9879 24012 9931 24064
rect 9801 23947 9853 23999
rect 9879 23947 9931 23999
rect 9801 23882 9853 23934
rect 9879 23882 9931 23934
rect 9801 23817 9853 23869
rect 9879 23817 9931 23869
rect 9801 23752 9853 23804
rect 9879 23752 9931 23804
rect 9801 23687 9853 23739
rect 9879 23687 9931 23739
rect 9801 23622 9853 23674
rect 9879 23622 9931 23674
rect 9801 23557 9853 23609
rect 9879 23557 9931 23609
rect 9801 23492 9853 23544
rect 9879 23492 9931 23544
rect 9801 23427 9853 23479
rect 9879 23427 9931 23479
rect 9801 23362 9853 23414
rect 9879 23362 9931 23414
rect 9801 23297 9853 23349
rect 9879 23297 9931 23349
rect 9801 20373 9853 20425
rect 9879 20373 9931 20425
rect 9801 20309 9853 20361
rect 9879 20309 9931 20361
rect 9801 20245 9853 20297
rect 9879 20245 9931 20297
rect 9801 20181 9853 20233
rect 9879 20181 9931 20233
rect 9801 20117 9853 20169
rect 9879 20117 9931 20169
rect 9801 20053 9853 20105
rect 9879 20053 9931 20105
rect 9801 19989 9853 20041
rect 9879 19989 9931 20041
rect 9801 19925 9853 19977
rect 9879 19925 9931 19977
rect 9801 19861 9853 19913
rect 9879 19861 9931 19913
rect 9801 19797 9853 19849
rect 9879 19797 9931 19849
rect 9801 19733 9853 19785
rect 9879 19733 9931 19785
rect 9801 19669 9853 19721
rect 9879 19669 9931 19721
rect 9801 19605 9853 19657
rect 9879 19605 9931 19657
rect 9801 19541 9853 19593
rect 9879 19541 9931 19593
rect 9801 19477 9853 19529
rect 9879 19477 9931 19529
rect 9801 19412 9853 19464
rect 9879 19412 9931 19464
rect 9801 19347 9853 19399
rect 9879 19347 9931 19399
rect 9801 19282 9853 19334
rect 9879 19282 9931 19334
rect 9801 19217 9853 19269
rect 9879 19217 9931 19269
rect 9801 19152 9853 19204
rect 9879 19152 9931 19204
rect 9801 19087 9853 19139
rect 9879 19087 9931 19139
rect 9801 19022 9853 19074
rect 9879 19022 9931 19074
rect 9801 18957 9853 19009
rect 9879 18957 9931 19009
rect 9801 18892 9853 18944
rect 9879 18892 9931 18944
rect 9801 18827 9853 18879
rect 9879 18827 9931 18879
rect 9801 18762 9853 18814
rect 9879 18762 9931 18814
rect 9801 18697 9853 18749
rect 9879 18697 9931 18749
rect 9801 15773 9853 15825
rect 9879 15773 9931 15825
rect 9801 15709 9853 15761
rect 9879 15709 9931 15761
rect 9801 15645 9853 15697
rect 9879 15645 9931 15697
rect 9801 15581 9853 15633
rect 9879 15581 9931 15633
rect 9801 15517 9853 15569
rect 9879 15517 9931 15569
rect 9801 15453 9853 15505
rect 9879 15453 9931 15505
rect 9801 15389 9853 15441
rect 9879 15389 9931 15441
rect 9801 15325 9853 15377
rect 9879 15325 9931 15377
rect 9801 15261 9853 15313
rect 9879 15261 9931 15313
rect 9801 15197 9853 15249
rect 9879 15197 9931 15249
rect 9801 15133 9853 15185
rect 9879 15133 9931 15185
rect 9801 15069 9853 15121
rect 9879 15069 9931 15121
rect 9801 15005 9853 15057
rect 9879 15005 9931 15057
rect 9801 14941 9853 14993
rect 9879 14941 9931 14993
rect 9801 14877 9853 14929
rect 9879 14877 9931 14929
rect 9801 14812 9853 14864
rect 9879 14812 9931 14864
rect 9801 14747 9853 14799
rect 9879 14747 9931 14799
rect 9801 14682 9853 14734
rect 9879 14682 9931 14734
rect 9801 14617 9853 14669
rect 9879 14617 9931 14669
rect 9801 14552 9853 14604
rect 9879 14552 9931 14604
rect 9801 14487 9853 14539
rect 9879 14487 9931 14539
rect 9801 14422 9853 14474
rect 9879 14422 9931 14474
rect 9801 14357 9853 14409
rect 9879 14357 9931 14409
rect 9801 14292 9853 14344
rect 9879 14292 9931 14344
rect 9801 14227 9853 14279
rect 9879 14227 9931 14279
rect 9801 14162 9853 14214
rect 9879 14162 9931 14214
rect 9801 14097 9853 14149
rect 9879 14097 9931 14149
rect 9801 11173 9853 11225
rect 9879 11173 9931 11225
rect 9801 11109 9853 11161
rect 9879 11109 9931 11161
rect 9801 11045 9853 11097
rect 9879 11045 9931 11097
rect 9801 10981 9853 11033
rect 9879 10981 9931 11033
rect 9801 10917 9853 10969
rect 9879 10917 9931 10969
rect 9801 10853 9853 10905
rect 9879 10853 9931 10905
rect 9801 10789 9853 10841
rect 9879 10789 9931 10841
rect 9801 10725 9853 10777
rect 9879 10725 9931 10777
rect 9801 10661 9853 10713
rect 9879 10661 9931 10713
rect 9801 10597 9853 10649
rect 9879 10597 9931 10649
rect 9801 10533 9853 10585
rect 9879 10533 9931 10585
rect 9801 10469 9853 10521
rect 9879 10469 9931 10521
rect 9801 10405 9853 10457
rect 9879 10405 9931 10457
rect 9801 10341 9853 10393
rect 9879 10341 9931 10393
rect 9801 10277 9853 10329
rect 9879 10277 9931 10329
rect 9801 10212 9853 10264
rect 9879 10212 9931 10264
rect 9801 10147 9853 10199
rect 9879 10147 9931 10199
rect 9801 10082 9853 10134
rect 9879 10082 9931 10134
rect 9801 10017 9853 10069
rect 9879 10017 9931 10069
rect 9801 9952 9853 10004
rect 9879 9952 9931 10004
rect 9801 9887 9853 9939
rect 9879 9887 9931 9939
rect 9801 9822 9853 9874
rect 9879 9822 9931 9874
rect 9801 9757 9853 9809
rect 9879 9757 9931 9809
rect 9801 9692 9853 9744
rect 9879 9692 9931 9744
rect 9801 9627 9853 9679
rect 9879 9627 9931 9679
rect 9801 9562 9853 9614
rect 9879 9562 9931 9614
rect 9801 9497 9853 9549
rect 9879 9497 9931 9549
rect 10232 36238 10237 36290
rect 10237 36238 10284 36290
rect 10300 36238 10352 36290
rect 10368 36238 10415 36290
rect 10415 36238 10420 36290
rect 10232 36174 10237 36226
rect 10237 36174 10284 36226
rect 10300 36174 10352 36226
rect 10368 36174 10415 36226
rect 10415 36174 10420 36226
rect 10232 36110 10237 36162
rect 10237 36110 10284 36162
rect 10300 36110 10352 36162
rect 10368 36110 10415 36162
rect 10415 36110 10420 36162
rect 10232 36046 10237 36098
rect 10237 36046 10284 36098
rect 10300 36046 10352 36098
rect 10368 36046 10415 36098
rect 10415 36046 10420 36098
rect 10232 35982 10237 36034
rect 10237 35982 10284 36034
rect 10300 35982 10352 36034
rect 10368 35982 10415 36034
rect 10415 35982 10420 36034
rect 10232 35918 10237 35970
rect 10237 35918 10284 35970
rect 10300 35918 10352 35970
rect 10368 35918 10415 35970
rect 10415 35918 10420 35970
rect 10232 35854 10237 35906
rect 10237 35854 10284 35906
rect 10300 35854 10352 35906
rect 10368 35854 10415 35906
rect 10415 35854 10420 35906
rect 10232 35790 10237 35842
rect 10237 35790 10284 35842
rect 10300 35790 10352 35842
rect 10368 35790 10415 35842
rect 10415 35790 10420 35842
rect 10232 35726 10237 35778
rect 10237 35726 10284 35778
rect 10300 35726 10352 35778
rect 10368 35726 10415 35778
rect 10415 35726 10420 35778
rect 10232 35662 10237 35714
rect 10237 35662 10284 35714
rect 10300 35662 10352 35714
rect 10368 35662 10415 35714
rect 10415 35662 10420 35714
rect 10232 35598 10237 35650
rect 10237 35598 10284 35650
rect 10300 35598 10352 35650
rect 10368 35598 10415 35650
rect 10415 35598 10420 35650
rect 10232 35534 10237 35586
rect 10237 35534 10284 35586
rect 10300 35534 10352 35586
rect 10368 35534 10415 35586
rect 10415 35534 10420 35586
rect 10232 35470 10237 35522
rect 10237 35470 10284 35522
rect 10300 35470 10352 35522
rect 10368 35470 10415 35522
rect 10415 35470 10420 35522
rect 10232 35406 10237 35458
rect 10237 35406 10284 35458
rect 10300 35406 10352 35458
rect 10368 35406 10415 35458
rect 10415 35406 10420 35458
rect 10232 35342 10237 35394
rect 10237 35342 10284 35394
rect 10300 35342 10352 35394
rect 10368 35342 10415 35394
rect 10415 35342 10420 35394
rect 10232 35277 10237 35329
rect 10237 35277 10284 35329
rect 10300 35277 10352 35329
rect 10368 35277 10415 35329
rect 10415 35277 10420 35329
rect 10232 35212 10237 35264
rect 10237 35212 10284 35264
rect 10300 35212 10352 35264
rect 10368 35212 10415 35264
rect 10415 35212 10420 35264
rect 10232 35147 10237 35199
rect 10237 35147 10284 35199
rect 10300 35147 10352 35199
rect 10368 35147 10415 35199
rect 10415 35147 10420 35199
rect 10232 35082 10237 35134
rect 10237 35082 10284 35134
rect 10300 35082 10352 35134
rect 10368 35082 10415 35134
rect 10415 35082 10420 35134
rect 10232 35017 10237 35069
rect 10237 35017 10284 35069
rect 10300 35017 10352 35069
rect 10368 35017 10415 35069
rect 10415 35017 10420 35069
rect 10232 34952 10237 35004
rect 10237 34952 10284 35004
rect 10300 34952 10352 35004
rect 10368 34952 10415 35004
rect 10415 34952 10420 35004
rect 10232 34887 10237 34939
rect 10237 34887 10284 34939
rect 10300 34887 10352 34939
rect 10368 34887 10415 34939
rect 10415 34887 10420 34939
rect 10232 34822 10237 34874
rect 10237 34822 10284 34874
rect 10300 34822 10352 34874
rect 10368 34822 10415 34874
rect 10415 34822 10420 34874
rect 10232 34757 10237 34809
rect 10237 34757 10284 34809
rect 10300 34757 10352 34809
rect 10368 34757 10415 34809
rect 10415 34757 10420 34809
rect 10232 34692 10237 34744
rect 10237 34692 10284 34744
rect 10300 34692 10352 34744
rect 10368 34692 10415 34744
rect 10415 34692 10420 34744
rect 10232 34627 10237 34679
rect 10237 34627 10284 34679
rect 10300 34627 10352 34679
rect 10368 34627 10415 34679
rect 10415 34627 10420 34679
rect 10232 34562 10237 34614
rect 10237 34562 10284 34614
rect 10300 34562 10352 34614
rect 10368 34562 10415 34614
rect 10415 34562 10420 34614
rect 10232 31638 10237 31690
rect 10237 31638 10284 31690
rect 10300 31638 10352 31690
rect 10368 31638 10415 31690
rect 10415 31638 10420 31690
rect 10232 31574 10237 31626
rect 10237 31574 10284 31626
rect 10300 31574 10352 31626
rect 10368 31574 10415 31626
rect 10415 31574 10420 31626
rect 10232 31510 10237 31562
rect 10237 31510 10284 31562
rect 10300 31510 10352 31562
rect 10368 31510 10415 31562
rect 10415 31510 10420 31562
rect 10232 31446 10237 31498
rect 10237 31446 10284 31498
rect 10300 31446 10352 31498
rect 10368 31446 10415 31498
rect 10415 31446 10420 31498
rect 10232 31382 10237 31434
rect 10237 31382 10284 31434
rect 10300 31382 10352 31434
rect 10368 31382 10415 31434
rect 10415 31382 10420 31434
rect 10232 31318 10237 31370
rect 10237 31318 10284 31370
rect 10300 31318 10352 31370
rect 10368 31318 10415 31370
rect 10415 31318 10420 31370
rect 10232 31254 10237 31306
rect 10237 31254 10284 31306
rect 10300 31254 10352 31306
rect 10368 31254 10415 31306
rect 10415 31254 10420 31306
rect 10232 31190 10237 31242
rect 10237 31190 10284 31242
rect 10300 31190 10352 31242
rect 10368 31190 10415 31242
rect 10415 31190 10420 31242
rect 10232 31126 10237 31178
rect 10237 31126 10284 31178
rect 10300 31126 10352 31178
rect 10368 31126 10415 31178
rect 10415 31126 10420 31178
rect 10232 31062 10237 31114
rect 10237 31062 10284 31114
rect 10300 31062 10352 31114
rect 10368 31062 10415 31114
rect 10415 31062 10420 31114
rect 10232 30998 10237 31050
rect 10237 30998 10284 31050
rect 10300 30998 10352 31050
rect 10368 30998 10415 31050
rect 10415 30998 10420 31050
rect 10232 30934 10237 30986
rect 10237 30934 10284 30986
rect 10300 30934 10352 30986
rect 10368 30934 10415 30986
rect 10415 30934 10420 30986
rect 10232 30870 10237 30922
rect 10237 30870 10284 30922
rect 10300 30870 10352 30922
rect 10368 30870 10415 30922
rect 10415 30870 10420 30922
rect 10232 30806 10237 30858
rect 10237 30806 10284 30858
rect 10300 30806 10352 30858
rect 10368 30806 10415 30858
rect 10415 30806 10420 30858
rect 10232 30742 10237 30794
rect 10237 30742 10284 30794
rect 10300 30742 10352 30794
rect 10368 30742 10415 30794
rect 10415 30742 10420 30794
rect 10232 30677 10237 30729
rect 10237 30677 10284 30729
rect 10300 30677 10352 30729
rect 10368 30677 10415 30729
rect 10415 30677 10420 30729
rect 10232 30612 10237 30664
rect 10237 30612 10284 30664
rect 10300 30612 10352 30664
rect 10368 30612 10415 30664
rect 10415 30612 10420 30664
rect 10232 30547 10237 30599
rect 10237 30547 10284 30599
rect 10300 30547 10352 30599
rect 10368 30547 10415 30599
rect 10415 30547 10420 30599
rect 10232 30482 10237 30534
rect 10237 30482 10284 30534
rect 10300 30482 10352 30534
rect 10368 30482 10415 30534
rect 10415 30482 10420 30534
rect 10232 30417 10237 30469
rect 10237 30417 10284 30469
rect 10300 30417 10352 30469
rect 10368 30417 10415 30469
rect 10415 30417 10420 30469
rect 10232 30352 10237 30404
rect 10237 30352 10284 30404
rect 10300 30352 10352 30404
rect 10368 30352 10415 30404
rect 10415 30352 10420 30404
rect 10232 30287 10237 30339
rect 10237 30287 10284 30339
rect 10300 30287 10352 30339
rect 10368 30287 10415 30339
rect 10415 30287 10420 30339
rect 10232 30222 10237 30274
rect 10237 30222 10284 30274
rect 10300 30222 10352 30274
rect 10368 30222 10415 30274
rect 10415 30222 10420 30274
rect 10232 30157 10237 30209
rect 10237 30157 10284 30209
rect 10300 30157 10352 30209
rect 10368 30157 10415 30209
rect 10415 30157 10420 30209
rect 10232 30092 10237 30144
rect 10237 30092 10284 30144
rect 10300 30092 10352 30144
rect 10368 30092 10415 30144
rect 10415 30092 10420 30144
rect 10232 30027 10237 30079
rect 10237 30027 10284 30079
rect 10300 30027 10352 30079
rect 10368 30027 10415 30079
rect 10415 30027 10420 30079
rect 10232 29962 10237 30014
rect 10237 29962 10284 30014
rect 10300 29962 10352 30014
rect 10368 29962 10415 30014
rect 10415 29962 10420 30014
rect 10232 27038 10237 27090
rect 10237 27038 10284 27090
rect 10300 27038 10352 27090
rect 10368 27038 10415 27090
rect 10415 27038 10420 27090
rect 10232 26974 10237 27026
rect 10237 26974 10284 27026
rect 10300 26974 10352 27026
rect 10368 26974 10415 27026
rect 10415 26974 10420 27026
rect 10232 26910 10237 26962
rect 10237 26910 10284 26962
rect 10300 26910 10352 26962
rect 10368 26910 10415 26962
rect 10415 26910 10420 26962
rect 10232 26846 10237 26898
rect 10237 26846 10284 26898
rect 10300 26846 10352 26898
rect 10368 26846 10415 26898
rect 10415 26846 10420 26898
rect 10232 26782 10237 26834
rect 10237 26782 10284 26834
rect 10300 26782 10352 26834
rect 10368 26782 10415 26834
rect 10415 26782 10420 26834
rect 10232 26718 10237 26770
rect 10237 26718 10284 26770
rect 10300 26718 10352 26770
rect 10368 26718 10415 26770
rect 10415 26718 10420 26770
rect 10232 26654 10237 26706
rect 10237 26654 10284 26706
rect 10300 26654 10352 26706
rect 10368 26654 10415 26706
rect 10415 26654 10420 26706
rect 10232 26590 10237 26642
rect 10237 26590 10284 26642
rect 10300 26590 10352 26642
rect 10368 26590 10415 26642
rect 10415 26590 10420 26642
rect 10232 26526 10237 26578
rect 10237 26526 10284 26578
rect 10300 26526 10352 26578
rect 10368 26526 10415 26578
rect 10415 26526 10420 26578
rect 10232 26462 10237 26514
rect 10237 26462 10284 26514
rect 10300 26462 10352 26514
rect 10368 26462 10415 26514
rect 10415 26462 10420 26514
rect 10232 26398 10237 26450
rect 10237 26398 10284 26450
rect 10300 26398 10352 26450
rect 10368 26398 10415 26450
rect 10415 26398 10420 26450
rect 10232 26334 10237 26386
rect 10237 26334 10284 26386
rect 10300 26334 10352 26386
rect 10368 26334 10415 26386
rect 10415 26334 10420 26386
rect 10232 26270 10237 26322
rect 10237 26270 10284 26322
rect 10300 26270 10352 26322
rect 10368 26270 10415 26322
rect 10415 26270 10420 26322
rect 10232 26206 10237 26258
rect 10237 26206 10284 26258
rect 10300 26206 10352 26258
rect 10368 26206 10415 26258
rect 10415 26206 10420 26258
rect 10232 26142 10237 26194
rect 10237 26142 10284 26194
rect 10300 26142 10352 26194
rect 10368 26142 10415 26194
rect 10415 26142 10420 26194
rect 10232 26077 10237 26129
rect 10237 26077 10284 26129
rect 10300 26077 10352 26129
rect 10368 26077 10415 26129
rect 10415 26077 10420 26129
rect 10232 26012 10237 26064
rect 10237 26012 10284 26064
rect 10300 26012 10352 26064
rect 10368 26012 10415 26064
rect 10415 26012 10420 26064
rect 10232 25947 10237 25999
rect 10237 25947 10284 25999
rect 10300 25947 10352 25999
rect 10368 25947 10415 25999
rect 10415 25947 10420 25999
rect 10232 25882 10237 25934
rect 10237 25882 10284 25934
rect 10300 25882 10352 25934
rect 10368 25882 10415 25934
rect 10415 25882 10420 25934
rect 10232 25817 10237 25869
rect 10237 25817 10284 25869
rect 10300 25817 10352 25869
rect 10368 25817 10415 25869
rect 10415 25817 10420 25869
rect 10232 25752 10237 25804
rect 10237 25752 10284 25804
rect 10300 25752 10352 25804
rect 10368 25752 10415 25804
rect 10415 25752 10420 25804
rect 10232 25687 10237 25739
rect 10237 25687 10284 25739
rect 10300 25687 10352 25739
rect 10368 25687 10415 25739
rect 10415 25687 10420 25739
rect 10232 25622 10237 25674
rect 10237 25622 10284 25674
rect 10300 25622 10352 25674
rect 10368 25622 10415 25674
rect 10415 25622 10420 25674
rect 10232 25557 10237 25609
rect 10237 25557 10284 25609
rect 10300 25557 10352 25609
rect 10368 25557 10415 25609
rect 10415 25557 10420 25609
rect 10232 25492 10237 25544
rect 10237 25492 10284 25544
rect 10300 25492 10352 25544
rect 10368 25492 10415 25544
rect 10415 25492 10420 25544
rect 10232 25427 10237 25479
rect 10237 25427 10284 25479
rect 10300 25427 10352 25479
rect 10368 25427 10415 25479
rect 10415 25427 10420 25479
rect 10232 25362 10237 25414
rect 10237 25362 10284 25414
rect 10300 25362 10352 25414
rect 10368 25362 10415 25414
rect 10415 25362 10420 25414
rect 10232 22438 10237 22490
rect 10237 22438 10284 22490
rect 10300 22438 10352 22490
rect 10368 22438 10415 22490
rect 10415 22438 10420 22490
rect 10232 22374 10237 22426
rect 10237 22374 10284 22426
rect 10300 22374 10352 22426
rect 10368 22374 10415 22426
rect 10415 22374 10420 22426
rect 10232 22310 10237 22362
rect 10237 22310 10284 22362
rect 10300 22310 10352 22362
rect 10368 22310 10415 22362
rect 10415 22310 10420 22362
rect 10232 22246 10237 22298
rect 10237 22246 10284 22298
rect 10300 22246 10352 22298
rect 10368 22246 10415 22298
rect 10415 22246 10420 22298
rect 10232 22182 10237 22234
rect 10237 22182 10284 22234
rect 10300 22182 10352 22234
rect 10368 22182 10415 22234
rect 10415 22182 10420 22234
rect 10232 22118 10237 22170
rect 10237 22118 10284 22170
rect 10300 22118 10352 22170
rect 10368 22118 10415 22170
rect 10415 22118 10420 22170
rect 10232 22054 10237 22106
rect 10237 22054 10284 22106
rect 10300 22054 10352 22106
rect 10368 22054 10415 22106
rect 10415 22054 10420 22106
rect 10232 21990 10237 22042
rect 10237 21990 10284 22042
rect 10300 21990 10352 22042
rect 10368 21990 10415 22042
rect 10415 21990 10420 22042
rect 10232 21926 10237 21978
rect 10237 21926 10284 21978
rect 10300 21926 10352 21978
rect 10368 21926 10415 21978
rect 10415 21926 10420 21978
rect 10232 21862 10237 21914
rect 10237 21862 10284 21914
rect 10300 21862 10352 21914
rect 10368 21862 10415 21914
rect 10415 21862 10420 21914
rect 10232 21798 10237 21850
rect 10237 21798 10284 21850
rect 10300 21798 10352 21850
rect 10368 21798 10415 21850
rect 10415 21798 10420 21850
rect 10232 21734 10237 21786
rect 10237 21734 10284 21786
rect 10300 21734 10352 21786
rect 10368 21734 10415 21786
rect 10415 21734 10420 21786
rect 10232 21670 10237 21722
rect 10237 21670 10284 21722
rect 10300 21670 10352 21722
rect 10368 21670 10415 21722
rect 10415 21670 10420 21722
rect 10232 21606 10237 21658
rect 10237 21606 10284 21658
rect 10300 21606 10352 21658
rect 10368 21606 10415 21658
rect 10415 21606 10420 21658
rect 10232 21542 10237 21594
rect 10237 21542 10284 21594
rect 10300 21542 10352 21594
rect 10368 21542 10415 21594
rect 10415 21542 10420 21594
rect 10232 21477 10237 21529
rect 10237 21477 10284 21529
rect 10300 21477 10352 21529
rect 10368 21477 10415 21529
rect 10415 21477 10420 21529
rect 10232 21412 10237 21464
rect 10237 21412 10284 21464
rect 10300 21412 10352 21464
rect 10368 21412 10415 21464
rect 10415 21412 10420 21464
rect 10232 21347 10237 21399
rect 10237 21347 10284 21399
rect 10300 21347 10352 21399
rect 10368 21347 10415 21399
rect 10415 21347 10420 21399
rect 10232 21282 10237 21334
rect 10237 21282 10284 21334
rect 10300 21282 10352 21334
rect 10368 21282 10415 21334
rect 10415 21282 10420 21334
rect 10232 21217 10237 21269
rect 10237 21217 10284 21269
rect 10300 21217 10352 21269
rect 10368 21217 10415 21269
rect 10415 21217 10420 21269
rect 10232 21152 10237 21204
rect 10237 21152 10284 21204
rect 10300 21152 10352 21204
rect 10368 21152 10415 21204
rect 10415 21152 10420 21204
rect 10232 21087 10237 21139
rect 10237 21087 10284 21139
rect 10300 21087 10352 21139
rect 10368 21087 10415 21139
rect 10415 21087 10420 21139
rect 10232 21022 10237 21074
rect 10237 21022 10284 21074
rect 10300 21022 10352 21074
rect 10368 21022 10415 21074
rect 10415 21022 10420 21074
rect 10232 20957 10237 21009
rect 10237 20957 10284 21009
rect 10300 20957 10352 21009
rect 10368 20957 10415 21009
rect 10415 20957 10420 21009
rect 10232 20892 10237 20944
rect 10237 20892 10284 20944
rect 10300 20892 10352 20944
rect 10368 20892 10415 20944
rect 10415 20892 10420 20944
rect 10232 20827 10237 20879
rect 10237 20827 10284 20879
rect 10300 20827 10352 20879
rect 10368 20827 10415 20879
rect 10415 20827 10420 20879
rect 10232 20762 10237 20814
rect 10237 20762 10284 20814
rect 10300 20762 10352 20814
rect 10368 20762 10415 20814
rect 10415 20762 10420 20814
rect 10232 17838 10237 17890
rect 10237 17838 10284 17890
rect 10300 17838 10352 17890
rect 10368 17838 10415 17890
rect 10415 17838 10420 17890
rect 10232 17774 10237 17826
rect 10237 17774 10284 17826
rect 10300 17774 10352 17826
rect 10368 17774 10415 17826
rect 10415 17774 10420 17826
rect 10232 17710 10237 17762
rect 10237 17710 10284 17762
rect 10300 17710 10352 17762
rect 10368 17710 10415 17762
rect 10415 17710 10420 17762
rect 10232 17646 10237 17698
rect 10237 17646 10284 17698
rect 10300 17646 10352 17698
rect 10368 17646 10415 17698
rect 10415 17646 10420 17698
rect 10232 17582 10237 17634
rect 10237 17582 10284 17634
rect 10300 17582 10352 17634
rect 10368 17582 10415 17634
rect 10415 17582 10420 17634
rect 10232 17518 10237 17570
rect 10237 17518 10284 17570
rect 10300 17518 10352 17570
rect 10368 17518 10415 17570
rect 10415 17518 10420 17570
rect 10232 17454 10237 17506
rect 10237 17454 10284 17506
rect 10300 17454 10352 17506
rect 10368 17454 10415 17506
rect 10415 17454 10420 17506
rect 10232 17390 10237 17442
rect 10237 17390 10284 17442
rect 10300 17390 10352 17442
rect 10368 17390 10415 17442
rect 10415 17390 10420 17442
rect 10232 17326 10237 17378
rect 10237 17326 10284 17378
rect 10300 17326 10352 17378
rect 10368 17326 10415 17378
rect 10415 17326 10420 17378
rect 10232 17262 10237 17314
rect 10237 17262 10284 17314
rect 10300 17262 10352 17314
rect 10368 17262 10415 17314
rect 10415 17262 10420 17314
rect 10232 17198 10237 17250
rect 10237 17198 10284 17250
rect 10300 17198 10352 17250
rect 10368 17198 10415 17250
rect 10415 17198 10420 17250
rect 10232 17134 10237 17186
rect 10237 17134 10284 17186
rect 10300 17134 10352 17186
rect 10368 17134 10415 17186
rect 10415 17134 10420 17186
rect 10232 17070 10237 17122
rect 10237 17070 10284 17122
rect 10300 17070 10352 17122
rect 10368 17070 10415 17122
rect 10415 17070 10420 17122
rect 10232 17006 10237 17058
rect 10237 17006 10284 17058
rect 10300 17006 10352 17058
rect 10368 17006 10415 17058
rect 10415 17006 10420 17058
rect 10232 16942 10237 16994
rect 10237 16942 10284 16994
rect 10300 16942 10352 16994
rect 10368 16942 10415 16994
rect 10415 16942 10420 16994
rect 10232 16877 10237 16929
rect 10237 16877 10284 16929
rect 10300 16877 10352 16929
rect 10368 16877 10415 16929
rect 10415 16877 10420 16929
rect 10232 16812 10237 16864
rect 10237 16812 10284 16864
rect 10300 16812 10352 16864
rect 10368 16812 10415 16864
rect 10415 16812 10420 16864
rect 10232 16747 10237 16799
rect 10237 16747 10284 16799
rect 10300 16747 10352 16799
rect 10368 16747 10415 16799
rect 10415 16747 10420 16799
rect 10232 16682 10237 16734
rect 10237 16682 10284 16734
rect 10300 16682 10352 16734
rect 10368 16682 10415 16734
rect 10415 16682 10420 16734
rect 10232 16617 10237 16669
rect 10237 16617 10284 16669
rect 10300 16617 10352 16669
rect 10368 16617 10415 16669
rect 10415 16617 10420 16669
rect 10232 16552 10237 16604
rect 10237 16552 10284 16604
rect 10300 16552 10352 16604
rect 10368 16552 10415 16604
rect 10415 16552 10420 16604
rect 10232 16487 10237 16539
rect 10237 16487 10284 16539
rect 10300 16487 10352 16539
rect 10368 16487 10415 16539
rect 10415 16487 10420 16539
rect 10232 16422 10237 16474
rect 10237 16422 10284 16474
rect 10300 16422 10352 16474
rect 10368 16422 10415 16474
rect 10415 16422 10420 16474
rect 10232 16357 10237 16409
rect 10237 16357 10284 16409
rect 10300 16357 10352 16409
rect 10368 16357 10415 16409
rect 10415 16357 10420 16409
rect 10232 16292 10237 16344
rect 10237 16292 10284 16344
rect 10300 16292 10352 16344
rect 10368 16292 10415 16344
rect 10415 16292 10420 16344
rect 10232 16227 10237 16279
rect 10237 16227 10284 16279
rect 10300 16227 10352 16279
rect 10368 16227 10415 16279
rect 10415 16227 10420 16279
rect 10232 16162 10237 16214
rect 10237 16162 10284 16214
rect 10300 16162 10352 16214
rect 10368 16162 10415 16214
rect 10415 16162 10420 16214
rect 10232 13238 10237 13290
rect 10237 13238 10284 13290
rect 10300 13238 10352 13290
rect 10368 13238 10415 13290
rect 10415 13238 10420 13290
rect 10232 13174 10237 13226
rect 10237 13174 10284 13226
rect 10300 13174 10352 13226
rect 10368 13174 10415 13226
rect 10415 13174 10420 13226
rect 10232 13110 10237 13162
rect 10237 13110 10284 13162
rect 10300 13110 10352 13162
rect 10368 13110 10415 13162
rect 10415 13110 10420 13162
rect 10232 13046 10237 13098
rect 10237 13046 10284 13098
rect 10300 13046 10352 13098
rect 10368 13046 10415 13098
rect 10415 13046 10420 13098
rect 10232 12982 10237 13034
rect 10237 12982 10284 13034
rect 10300 12982 10352 13034
rect 10368 12982 10415 13034
rect 10415 12982 10420 13034
rect 10232 12918 10237 12970
rect 10237 12918 10284 12970
rect 10300 12918 10352 12970
rect 10368 12918 10415 12970
rect 10415 12918 10420 12970
rect 10232 12854 10237 12906
rect 10237 12854 10284 12906
rect 10300 12854 10352 12906
rect 10368 12854 10415 12906
rect 10415 12854 10420 12906
rect 10232 12790 10237 12842
rect 10237 12790 10284 12842
rect 10300 12790 10352 12842
rect 10368 12790 10415 12842
rect 10415 12790 10420 12842
rect 10232 12726 10237 12778
rect 10237 12726 10284 12778
rect 10300 12726 10352 12778
rect 10368 12726 10415 12778
rect 10415 12726 10420 12778
rect 10232 12662 10237 12714
rect 10237 12662 10284 12714
rect 10300 12662 10352 12714
rect 10368 12662 10415 12714
rect 10415 12662 10420 12714
rect 10232 12598 10237 12650
rect 10237 12598 10284 12650
rect 10300 12598 10352 12650
rect 10368 12598 10415 12650
rect 10415 12598 10420 12650
rect 10232 12534 10237 12586
rect 10237 12534 10284 12586
rect 10300 12534 10352 12586
rect 10368 12534 10415 12586
rect 10415 12534 10420 12586
rect 10232 12470 10237 12522
rect 10237 12470 10284 12522
rect 10300 12470 10352 12522
rect 10368 12470 10415 12522
rect 10415 12470 10420 12522
rect 10232 12406 10237 12458
rect 10237 12406 10284 12458
rect 10300 12406 10352 12458
rect 10368 12406 10415 12458
rect 10415 12406 10420 12458
rect 10232 12342 10237 12394
rect 10237 12342 10284 12394
rect 10300 12342 10352 12394
rect 10368 12342 10415 12394
rect 10415 12342 10420 12394
rect 10232 12277 10237 12329
rect 10237 12277 10284 12329
rect 10300 12277 10352 12329
rect 10368 12277 10415 12329
rect 10415 12277 10420 12329
rect 10232 12212 10237 12264
rect 10237 12212 10284 12264
rect 10300 12212 10352 12264
rect 10368 12212 10415 12264
rect 10415 12212 10420 12264
rect 10232 12147 10237 12199
rect 10237 12147 10284 12199
rect 10300 12147 10352 12199
rect 10368 12147 10415 12199
rect 10415 12147 10420 12199
rect 10232 12082 10237 12134
rect 10237 12082 10284 12134
rect 10300 12082 10352 12134
rect 10368 12082 10415 12134
rect 10415 12082 10420 12134
rect 10232 12017 10237 12069
rect 10237 12017 10284 12069
rect 10300 12017 10352 12069
rect 10368 12017 10415 12069
rect 10415 12017 10420 12069
rect 10232 11952 10237 12004
rect 10237 11952 10284 12004
rect 10300 11952 10352 12004
rect 10368 11952 10415 12004
rect 10415 11952 10420 12004
rect 10232 11887 10237 11939
rect 10237 11887 10284 11939
rect 10300 11887 10352 11939
rect 10368 11887 10415 11939
rect 10415 11887 10420 11939
rect 10232 11822 10237 11874
rect 10237 11822 10284 11874
rect 10300 11822 10352 11874
rect 10368 11822 10415 11874
rect 10415 11822 10420 11874
rect 10232 11757 10237 11809
rect 10237 11757 10284 11809
rect 10300 11757 10352 11809
rect 10368 11757 10415 11809
rect 10415 11757 10420 11809
rect 10232 11692 10237 11744
rect 10237 11692 10284 11744
rect 10300 11692 10352 11744
rect 10368 11692 10415 11744
rect 10415 11692 10420 11744
rect 10232 11627 10237 11679
rect 10237 11627 10284 11679
rect 10300 11627 10352 11679
rect 10368 11627 10415 11679
rect 10415 11627 10420 11679
rect 10232 11562 10237 11614
rect 10237 11562 10284 11614
rect 10300 11562 10352 11614
rect 10368 11562 10415 11614
rect 10415 11562 10420 11614
rect 10721 37945 10773 37997
rect 10799 37945 10851 37997
rect 10721 37877 10773 37929
rect 10799 37877 10851 37929
rect 10721 37809 10773 37861
rect 10799 37809 10851 37861
rect 10721 37741 10773 37793
rect 10799 37741 10851 37793
rect 10721 37673 10773 37725
rect 10799 37673 10851 37725
rect 10721 37605 10773 37657
rect 10799 37605 10851 37657
rect 10721 37537 10773 37589
rect 10799 37537 10851 37589
rect 10721 37469 10773 37521
rect 10799 37469 10851 37521
rect 10721 37401 10773 37453
rect 10799 37401 10851 37453
rect 10721 37333 10773 37385
rect 10799 37333 10851 37385
rect 10721 37266 10773 37318
rect 10799 37266 10851 37318
rect 10721 37199 10773 37251
rect 10799 37199 10851 37251
rect 10721 37132 10773 37184
rect 10799 37132 10851 37184
rect 10721 37065 10773 37117
rect 10799 37065 10851 37117
rect 10721 34173 10773 34225
rect 10799 34173 10851 34225
rect 10721 34109 10773 34161
rect 10799 34109 10851 34161
rect 10721 34045 10773 34097
rect 10799 34045 10851 34097
rect 10721 33981 10773 34033
rect 10799 33981 10851 34033
rect 10721 33917 10773 33969
rect 10799 33917 10851 33969
rect 10721 33853 10773 33905
rect 10799 33853 10851 33905
rect 10721 33789 10773 33841
rect 10799 33789 10851 33841
rect 10721 33725 10773 33777
rect 10799 33725 10851 33777
rect 10721 33661 10773 33713
rect 10799 33661 10851 33713
rect 10721 33597 10773 33649
rect 10799 33597 10851 33649
rect 10721 33533 10773 33585
rect 10799 33533 10851 33585
rect 10721 33469 10773 33521
rect 10799 33469 10851 33521
rect 10721 33405 10773 33457
rect 10799 33405 10851 33457
rect 10721 33341 10773 33393
rect 10799 33341 10851 33393
rect 10721 33277 10773 33329
rect 10799 33277 10851 33329
rect 10721 33212 10773 33264
rect 10799 33212 10851 33264
rect 10721 33147 10773 33199
rect 10799 33147 10851 33199
rect 10721 33082 10773 33134
rect 10799 33082 10851 33134
rect 10721 33017 10773 33069
rect 10799 33017 10851 33069
rect 10721 32952 10773 33004
rect 10799 32952 10851 33004
rect 10721 32887 10773 32939
rect 10799 32887 10851 32939
rect 10721 32822 10773 32874
rect 10799 32822 10851 32874
rect 10721 32757 10773 32809
rect 10799 32757 10851 32809
rect 10721 32692 10773 32744
rect 10799 32692 10851 32744
rect 10721 32627 10773 32679
rect 10799 32627 10851 32679
rect 10721 32562 10773 32614
rect 10799 32562 10851 32614
rect 10721 32497 10773 32549
rect 10799 32497 10851 32549
rect 10721 29573 10773 29625
rect 10799 29573 10851 29625
rect 10721 29509 10773 29561
rect 10799 29509 10851 29561
rect 10721 29445 10773 29497
rect 10799 29445 10851 29497
rect 10721 29381 10773 29433
rect 10799 29381 10851 29433
rect 10721 29317 10773 29369
rect 10799 29317 10851 29369
rect 10721 29253 10773 29305
rect 10799 29253 10851 29305
rect 10721 29189 10773 29241
rect 10799 29189 10851 29241
rect 10721 29125 10773 29177
rect 10799 29125 10851 29177
rect 10721 29061 10773 29113
rect 10799 29061 10851 29113
rect 10721 28997 10773 29049
rect 10799 28997 10851 29049
rect 10721 28933 10773 28985
rect 10799 28933 10851 28985
rect 10721 28869 10773 28921
rect 10799 28869 10851 28921
rect 10721 28805 10773 28857
rect 10799 28805 10851 28857
rect 10721 28741 10773 28793
rect 10799 28741 10851 28793
rect 10721 28677 10773 28729
rect 10799 28677 10851 28729
rect 10721 28612 10773 28664
rect 10799 28612 10851 28664
rect 10721 28547 10773 28599
rect 10799 28547 10851 28599
rect 10721 28482 10773 28534
rect 10799 28482 10851 28534
rect 10721 28417 10773 28469
rect 10799 28417 10851 28469
rect 10721 28352 10773 28404
rect 10799 28352 10851 28404
rect 10721 28287 10773 28339
rect 10799 28287 10851 28339
rect 10721 28222 10773 28274
rect 10799 28222 10851 28274
rect 10721 28157 10773 28209
rect 10799 28157 10851 28209
rect 10721 28092 10773 28144
rect 10799 28092 10851 28144
rect 10721 28027 10773 28079
rect 10799 28027 10851 28079
rect 10721 27962 10773 28014
rect 10799 27962 10851 28014
rect 10721 27897 10773 27949
rect 10799 27897 10851 27949
rect 10721 24973 10773 25025
rect 10799 24973 10851 25025
rect 10721 24909 10773 24961
rect 10799 24909 10851 24961
rect 10721 24845 10773 24897
rect 10799 24845 10851 24897
rect 10721 24781 10773 24833
rect 10799 24781 10851 24833
rect 10721 24717 10773 24769
rect 10799 24717 10851 24769
rect 10721 24653 10773 24705
rect 10799 24653 10851 24705
rect 10721 24589 10773 24641
rect 10799 24589 10851 24641
rect 10721 24525 10773 24577
rect 10799 24525 10851 24577
rect 10721 24461 10773 24513
rect 10799 24461 10851 24513
rect 10721 24397 10773 24449
rect 10799 24397 10851 24449
rect 10721 24333 10773 24385
rect 10799 24333 10851 24385
rect 10721 24269 10773 24321
rect 10799 24269 10851 24321
rect 10721 24205 10773 24257
rect 10799 24205 10851 24257
rect 10721 24141 10773 24193
rect 10799 24141 10851 24193
rect 10721 24077 10773 24129
rect 10799 24077 10851 24129
rect 10721 24012 10773 24064
rect 10799 24012 10851 24064
rect 10721 23947 10773 23999
rect 10799 23947 10851 23999
rect 10721 23882 10773 23934
rect 10799 23882 10851 23934
rect 10721 23817 10773 23869
rect 10799 23817 10851 23869
rect 10721 23752 10773 23804
rect 10799 23752 10851 23804
rect 10721 23687 10773 23739
rect 10799 23687 10851 23739
rect 10721 23622 10773 23674
rect 10799 23622 10851 23674
rect 10721 23557 10773 23609
rect 10799 23557 10851 23609
rect 10721 23492 10773 23544
rect 10799 23492 10851 23544
rect 10721 23427 10773 23479
rect 10799 23427 10851 23479
rect 10721 23362 10773 23414
rect 10799 23362 10851 23414
rect 10721 23297 10773 23349
rect 10799 23297 10851 23349
rect 10721 20373 10773 20425
rect 10799 20373 10851 20425
rect 10721 20309 10773 20361
rect 10799 20309 10851 20361
rect 10721 20245 10773 20297
rect 10799 20245 10851 20297
rect 10721 20181 10773 20233
rect 10799 20181 10851 20233
rect 10721 20117 10773 20169
rect 10799 20117 10851 20169
rect 10721 20053 10773 20105
rect 10799 20053 10851 20105
rect 10721 19989 10773 20041
rect 10799 19989 10851 20041
rect 10721 19925 10773 19977
rect 10799 19925 10851 19977
rect 10721 19861 10773 19913
rect 10799 19861 10851 19913
rect 10721 19797 10773 19849
rect 10799 19797 10851 19849
rect 10721 19733 10773 19785
rect 10799 19733 10851 19785
rect 10721 19669 10773 19721
rect 10799 19669 10851 19721
rect 10721 19605 10773 19657
rect 10799 19605 10851 19657
rect 10721 19541 10773 19593
rect 10799 19541 10851 19593
rect 10721 19477 10773 19529
rect 10799 19477 10851 19529
rect 10721 19412 10773 19464
rect 10799 19412 10851 19464
rect 10721 19347 10773 19399
rect 10799 19347 10851 19399
rect 10721 19282 10773 19334
rect 10799 19282 10851 19334
rect 10721 19217 10773 19269
rect 10799 19217 10851 19269
rect 10721 19152 10773 19204
rect 10799 19152 10851 19204
rect 10721 19087 10773 19139
rect 10799 19087 10851 19139
rect 10721 19022 10773 19074
rect 10799 19022 10851 19074
rect 10721 18957 10773 19009
rect 10799 18957 10851 19009
rect 10721 18892 10773 18944
rect 10799 18892 10851 18944
rect 10721 18827 10773 18879
rect 10799 18827 10851 18879
rect 10721 18762 10773 18814
rect 10799 18762 10851 18814
rect 10721 18697 10773 18749
rect 10799 18697 10851 18749
rect 10721 15773 10773 15825
rect 10799 15773 10851 15825
rect 10721 15709 10773 15761
rect 10799 15709 10851 15761
rect 10721 15645 10773 15697
rect 10799 15645 10851 15697
rect 10721 15581 10773 15633
rect 10799 15581 10851 15633
rect 10721 15517 10773 15569
rect 10799 15517 10851 15569
rect 10721 15453 10773 15505
rect 10799 15453 10851 15505
rect 10721 15389 10773 15441
rect 10799 15389 10851 15441
rect 10721 15325 10773 15377
rect 10799 15325 10851 15377
rect 10721 15261 10773 15313
rect 10799 15261 10851 15313
rect 10721 15197 10773 15249
rect 10799 15197 10851 15249
rect 10721 15133 10773 15185
rect 10799 15133 10851 15185
rect 10721 15069 10773 15121
rect 10799 15069 10851 15121
rect 10721 15005 10773 15057
rect 10799 15005 10851 15057
rect 10721 14941 10773 14993
rect 10799 14941 10851 14993
rect 10721 14877 10773 14929
rect 10799 14877 10851 14929
rect 10721 14812 10773 14864
rect 10799 14812 10851 14864
rect 10721 14747 10773 14799
rect 10799 14747 10851 14799
rect 10721 14682 10773 14734
rect 10799 14682 10851 14734
rect 10721 14617 10773 14669
rect 10799 14617 10851 14669
rect 10721 14552 10773 14604
rect 10799 14552 10851 14604
rect 10721 14487 10773 14539
rect 10799 14487 10851 14539
rect 10721 14422 10773 14474
rect 10799 14422 10851 14474
rect 10721 14357 10773 14409
rect 10799 14357 10851 14409
rect 10721 14292 10773 14344
rect 10799 14292 10851 14344
rect 10721 14227 10773 14279
rect 10799 14227 10851 14279
rect 10721 14162 10773 14214
rect 10799 14162 10851 14214
rect 10721 14097 10773 14149
rect 10799 14097 10851 14149
rect 10721 11173 10773 11225
rect 10799 11173 10851 11225
rect 10721 11109 10773 11161
rect 10799 11109 10851 11161
rect 10721 11045 10773 11097
rect 10799 11045 10851 11097
rect 10721 10981 10773 11033
rect 10799 10981 10851 11033
rect 10721 10917 10773 10969
rect 10799 10917 10851 10969
rect 10721 10853 10773 10905
rect 10799 10853 10851 10905
rect 10721 10789 10773 10841
rect 10799 10789 10851 10841
rect 10721 10725 10773 10777
rect 10799 10725 10851 10777
rect 10721 10661 10773 10713
rect 10799 10661 10851 10713
rect 10721 10597 10773 10649
rect 10799 10597 10851 10649
rect 10721 10533 10773 10585
rect 10799 10533 10851 10585
rect 10721 10469 10773 10521
rect 10799 10469 10851 10521
rect 10721 10405 10773 10457
rect 10799 10405 10851 10457
rect 10721 10341 10773 10393
rect 10799 10341 10851 10393
rect 10721 10277 10773 10329
rect 10799 10277 10851 10329
rect 10721 10212 10773 10264
rect 10799 10212 10851 10264
rect 10721 10147 10773 10199
rect 10799 10147 10851 10199
rect 10721 10082 10773 10134
rect 10799 10082 10851 10134
rect 10721 10017 10773 10069
rect 10799 10017 10851 10069
rect 10721 9952 10773 10004
rect 10799 9952 10851 10004
rect 10721 9887 10773 9939
rect 10799 9887 10851 9939
rect 10721 9822 10773 9874
rect 10799 9822 10851 9874
rect 10721 9757 10773 9809
rect 10799 9757 10851 9809
rect 10721 9692 10773 9744
rect 10799 9692 10851 9744
rect 10721 9627 10773 9679
rect 10799 9627 10851 9679
rect 10721 9562 10773 9614
rect 10799 9562 10851 9614
rect 10721 9497 10773 9549
rect 10799 9497 10851 9549
rect 12072 38957 12077 39009
rect 12077 38957 12124 39009
rect 12140 38957 12192 39009
rect 12208 38957 12255 39009
rect 12255 38957 12260 39009
rect 12072 38892 12077 38944
rect 12077 38892 12124 38944
rect 12140 38892 12192 38944
rect 12208 38892 12255 38944
rect 12255 38892 12260 38944
rect 12072 38827 12077 38879
rect 12077 38827 12124 38879
rect 12140 38827 12192 38879
rect 12208 38827 12255 38879
rect 12255 38827 12260 38879
rect 12072 38762 12077 38814
rect 12077 38762 12124 38814
rect 12140 38762 12192 38814
rect 12208 38762 12255 38814
rect 12255 38762 12260 38814
rect 12072 38697 12077 38749
rect 12077 38697 12124 38749
rect 12140 38697 12192 38749
rect 12208 38697 12255 38749
rect 12255 38697 12260 38749
rect 12072 38632 12077 38684
rect 12077 38632 12124 38684
rect 12140 38632 12192 38684
rect 12208 38632 12255 38684
rect 12255 38632 12260 38684
rect 12072 38567 12077 38619
rect 12077 38567 12124 38619
rect 12140 38567 12192 38619
rect 12208 38567 12255 38619
rect 12255 38567 12260 38619
rect 12072 38502 12077 38554
rect 12077 38502 12124 38554
rect 12140 38502 12192 38554
rect 12208 38502 12255 38554
rect 12255 38502 12260 38554
rect 12072 38451 12124 38490
rect 12072 38438 12077 38451
rect 12077 38438 12111 38451
rect 12111 38438 12124 38451
rect 12140 38451 12192 38490
rect 12140 38438 12149 38451
rect 12149 38438 12183 38451
rect 12183 38438 12192 38451
rect 12208 38451 12260 38490
rect 12208 38438 12221 38451
rect 12221 38438 12255 38451
rect 12255 38438 12260 38451
rect 12072 38417 12077 38426
rect 12077 38417 12111 38426
rect 12111 38417 12124 38426
rect 12072 38378 12124 38417
rect 12072 38374 12077 38378
rect 12077 38374 12111 38378
rect 12111 38374 12124 38378
rect 12140 38417 12149 38426
rect 12149 38417 12183 38426
rect 12183 38417 12192 38426
rect 12140 38378 12192 38417
rect 12140 38374 12149 38378
rect 12149 38374 12183 38378
rect 12183 38374 12192 38378
rect 12208 38417 12221 38426
rect 12221 38417 12255 38426
rect 12255 38417 12260 38426
rect 12208 38378 12260 38417
rect 12208 38374 12221 38378
rect 12221 38374 12255 38378
rect 12255 38374 12260 38378
rect 12072 38344 12077 38362
rect 12077 38344 12111 38362
rect 12111 38344 12124 38362
rect 12072 38310 12124 38344
rect 12140 38344 12149 38362
rect 12149 38344 12183 38362
rect 12183 38344 12192 38362
rect 12140 38310 12192 38344
rect 12208 38344 12221 38362
rect 12221 38344 12255 38362
rect 12255 38344 12260 38362
rect 12208 38310 12260 38344
rect 12072 38271 12077 38298
rect 12077 38271 12111 38298
rect 12111 38271 12124 38298
rect 12072 38246 12124 38271
rect 12140 38271 12149 38298
rect 12149 38271 12183 38298
rect 12183 38271 12192 38298
rect 12140 38246 12192 38271
rect 12208 38271 12221 38298
rect 12221 38271 12255 38298
rect 12255 38271 12260 38298
rect 12208 38246 12260 38271
rect 12072 38232 12124 38234
rect 12072 38198 12077 38232
rect 12077 38198 12111 38232
rect 12111 38198 12124 38232
rect 12072 38182 12124 38198
rect 12140 38232 12192 38234
rect 12140 38198 12149 38232
rect 12149 38198 12183 38232
rect 12183 38198 12192 38232
rect 12140 38182 12192 38198
rect 12208 38232 12260 38234
rect 12208 38198 12221 38232
rect 12221 38198 12255 38232
rect 12255 38198 12260 38232
rect 12208 38182 12260 38198
rect 12072 38159 12124 38170
rect 12072 38125 12077 38159
rect 12077 38125 12111 38159
rect 12111 38125 12124 38159
rect 12072 38118 12124 38125
rect 12140 38159 12192 38170
rect 12140 38125 12149 38159
rect 12149 38125 12183 38159
rect 12183 38125 12192 38159
rect 12140 38118 12192 38125
rect 12208 38159 12260 38170
rect 12208 38125 12221 38159
rect 12221 38125 12255 38159
rect 12255 38125 12260 38159
rect 12208 38118 12260 38125
rect 11152 36238 11157 36290
rect 11157 36238 11204 36290
rect 11220 36238 11272 36290
rect 11288 36238 11335 36290
rect 11335 36238 11340 36290
rect 11152 36174 11157 36226
rect 11157 36174 11204 36226
rect 11220 36174 11272 36226
rect 11288 36174 11335 36226
rect 11335 36174 11340 36226
rect 11152 36110 11157 36162
rect 11157 36110 11204 36162
rect 11220 36110 11272 36162
rect 11288 36110 11335 36162
rect 11335 36110 11340 36162
rect 11152 36046 11157 36098
rect 11157 36046 11204 36098
rect 11220 36046 11272 36098
rect 11288 36046 11335 36098
rect 11335 36046 11340 36098
rect 11152 35982 11157 36034
rect 11157 35982 11204 36034
rect 11220 35982 11272 36034
rect 11288 35982 11335 36034
rect 11335 35982 11340 36034
rect 11152 35918 11157 35970
rect 11157 35918 11204 35970
rect 11220 35918 11272 35970
rect 11288 35918 11335 35970
rect 11335 35918 11340 35970
rect 11152 35854 11157 35906
rect 11157 35854 11204 35906
rect 11220 35854 11272 35906
rect 11288 35854 11335 35906
rect 11335 35854 11340 35906
rect 11152 35790 11157 35842
rect 11157 35790 11204 35842
rect 11220 35790 11272 35842
rect 11288 35790 11335 35842
rect 11335 35790 11340 35842
rect 11152 35726 11157 35778
rect 11157 35726 11204 35778
rect 11220 35726 11272 35778
rect 11288 35726 11335 35778
rect 11335 35726 11340 35778
rect 11152 35662 11157 35714
rect 11157 35662 11204 35714
rect 11220 35662 11272 35714
rect 11288 35662 11335 35714
rect 11335 35662 11340 35714
rect 11152 35598 11157 35650
rect 11157 35598 11204 35650
rect 11220 35598 11272 35650
rect 11288 35598 11335 35650
rect 11335 35598 11340 35650
rect 11152 35534 11157 35586
rect 11157 35534 11204 35586
rect 11220 35534 11272 35586
rect 11288 35534 11335 35586
rect 11335 35534 11340 35586
rect 11152 35470 11157 35522
rect 11157 35470 11204 35522
rect 11220 35470 11272 35522
rect 11288 35470 11335 35522
rect 11335 35470 11340 35522
rect 11152 35406 11157 35458
rect 11157 35406 11204 35458
rect 11220 35406 11272 35458
rect 11288 35406 11335 35458
rect 11335 35406 11340 35458
rect 11152 35342 11157 35394
rect 11157 35342 11204 35394
rect 11220 35342 11272 35394
rect 11288 35342 11335 35394
rect 11335 35342 11340 35394
rect 11152 35277 11157 35329
rect 11157 35277 11204 35329
rect 11220 35277 11272 35329
rect 11288 35277 11335 35329
rect 11335 35277 11340 35329
rect 11152 35212 11157 35264
rect 11157 35212 11204 35264
rect 11220 35212 11272 35264
rect 11288 35212 11335 35264
rect 11335 35212 11340 35264
rect 11152 35147 11157 35199
rect 11157 35147 11204 35199
rect 11220 35147 11272 35199
rect 11288 35147 11335 35199
rect 11335 35147 11340 35199
rect 11152 35082 11157 35134
rect 11157 35082 11204 35134
rect 11220 35082 11272 35134
rect 11288 35082 11335 35134
rect 11335 35082 11340 35134
rect 11152 35017 11157 35069
rect 11157 35017 11204 35069
rect 11220 35017 11272 35069
rect 11288 35017 11335 35069
rect 11335 35017 11340 35069
rect 11152 34952 11157 35004
rect 11157 34952 11204 35004
rect 11220 34952 11272 35004
rect 11288 34952 11335 35004
rect 11335 34952 11340 35004
rect 11152 34887 11157 34939
rect 11157 34887 11204 34939
rect 11220 34887 11272 34939
rect 11288 34887 11335 34939
rect 11335 34887 11340 34939
rect 11152 34822 11157 34874
rect 11157 34822 11204 34874
rect 11220 34822 11272 34874
rect 11288 34822 11335 34874
rect 11335 34822 11340 34874
rect 11152 34757 11157 34809
rect 11157 34757 11204 34809
rect 11220 34757 11272 34809
rect 11288 34757 11335 34809
rect 11335 34757 11340 34809
rect 11152 34692 11157 34744
rect 11157 34692 11204 34744
rect 11220 34692 11272 34744
rect 11288 34692 11335 34744
rect 11335 34692 11340 34744
rect 11152 34627 11157 34679
rect 11157 34627 11204 34679
rect 11220 34627 11272 34679
rect 11288 34627 11335 34679
rect 11335 34627 11340 34679
rect 11152 34562 11157 34614
rect 11157 34562 11204 34614
rect 11220 34562 11272 34614
rect 11288 34562 11335 34614
rect 11335 34562 11340 34614
rect 11152 31638 11157 31690
rect 11157 31638 11204 31690
rect 11220 31638 11272 31690
rect 11288 31638 11335 31690
rect 11335 31638 11340 31690
rect 11152 31574 11157 31626
rect 11157 31574 11204 31626
rect 11220 31574 11272 31626
rect 11288 31574 11335 31626
rect 11335 31574 11340 31626
rect 11152 31510 11157 31562
rect 11157 31510 11204 31562
rect 11220 31510 11272 31562
rect 11288 31510 11335 31562
rect 11335 31510 11340 31562
rect 11152 31446 11157 31498
rect 11157 31446 11204 31498
rect 11220 31446 11272 31498
rect 11288 31446 11335 31498
rect 11335 31446 11340 31498
rect 11152 31382 11157 31434
rect 11157 31382 11204 31434
rect 11220 31382 11272 31434
rect 11288 31382 11335 31434
rect 11335 31382 11340 31434
rect 11152 31318 11157 31370
rect 11157 31318 11204 31370
rect 11220 31318 11272 31370
rect 11288 31318 11335 31370
rect 11335 31318 11340 31370
rect 11152 31254 11157 31306
rect 11157 31254 11204 31306
rect 11220 31254 11272 31306
rect 11288 31254 11335 31306
rect 11335 31254 11340 31306
rect 11152 31190 11157 31242
rect 11157 31190 11204 31242
rect 11220 31190 11272 31242
rect 11288 31190 11335 31242
rect 11335 31190 11340 31242
rect 11152 31126 11157 31178
rect 11157 31126 11204 31178
rect 11220 31126 11272 31178
rect 11288 31126 11335 31178
rect 11335 31126 11340 31178
rect 11152 31062 11157 31114
rect 11157 31062 11204 31114
rect 11220 31062 11272 31114
rect 11288 31062 11335 31114
rect 11335 31062 11340 31114
rect 11152 30998 11157 31050
rect 11157 30998 11204 31050
rect 11220 30998 11272 31050
rect 11288 30998 11335 31050
rect 11335 30998 11340 31050
rect 11152 30934 11157 30986
rect 11157 30934 11204 30986
rect 11220 30934 11272 30986
rect 11288 30934 11335 30986
rect 11335 30934 11340 30986
rect 11152 30870 11157 30922
rect 11157 30870 11204 30922
rect 11220 30870 11272 30922
rect 11288 30870 11335 30922
rect 11335 30870 11340 30922
rect 11152 30806 11157 30858
rect 11157 30806 11204 30858
rect 11220 30806 11272 30858
rect 11288 30806 11335 30858
rect 11335 30806 11340 30858
rect 11152 30742 11157 30794
rect 11157 30742 11204 30794
rect 11220 30742 11272 30794
rect 11288 30742 11335 30794
rect 11335 30742 11340 30794
rect 11152 30677 11157 30729
rect 11157 30677 11204 30729
rect 11220 30677 11272 30729
rect 11288 30677 11335 30729
rect 11335 30677 11340 30729
rect 11152 30612 11157 30664
rect 11157 30612 11204 30664
rect 11220 30612 11272 30664
rect 11288 30612 11335 30664
rect 11335 30612 11340 30664
rect 11152 30547 11157 30599
rect 11157 30547 11204 30599
rect 11220 30547 11272 30599
rect 11288 30547 11335 30599
rect 11335 30547 11340 30599
rect 11152 30482 11157 30534
rect 11157 30482 11204 30534
rect 11220 30482 11272 30534
rect 11288 30482 11335 30534
rect 11335 30482 11340 30534
rect 11152 30417 11157 30469
rect 11157 30417 11204 30469
rect 11220 30417 11272 30469
rect 11288 30417 11335 30469
rect 11335 30417 11340 30469
rect 11152 30352 11157 30404
rect 11157 30352 11204 30404
rect 11220 30352 11272 30404
rect 11288 30352 11335 30404
rect 11335 30352 11340 30404
rect 11152 30287 11157 30339
rect 11157 30287 11204 30339
rect 11220 30287 11272 30339
rect 11288 30287 11335 30339
rect 11335 30287 11340 30339
rect 11152 30222 11157 30274
rect 11157 30222 11204 30274
rect 11220 30222 11272 30274
rect 11288 30222 11335 30274
rect 11335 30222 11340 30274
rect 11152 30157 11157 30209
rect 11157 30157 11204 30209
rect 11220 30157 11272 30209
rect 11288 30157 11335 30209
rect 11335 30157 11340 30209
rect 11152 30092 11157 30144
rect 11157 30092 11204 30144
rect 11220 30092 11272 30144
rect 11288 30092 11335 30144
rect 11335 30092 11340 30144
rect 11152 30027 11157 30079
rect 11157 30027 11204 30079
rect 11220 30027 11272 30079
rect 11288 30027 11335 30079
rect 11335 30027 11340 30079
rect 11152 29962 11157 30014
rect 11157 29962 11204 30014
rect 11220 29962 11272 30014
rect 11288 29962 11335 30014
rect 11335 29962 11340 30014
rect 11152 27038 11157 27090
rect 11157 27038 11204 27090
rect 11220 27038 11272 27090
rect 11288 27038 11335 27090
rect 11335 27038 11340 27090
rect 11152 26974 11157 27026
rect 11157 26974 11204 27026
rect 11220 26974 11272 27026
rect 11288 26974 11335 27026
rect 11335 26974 11340 27026
rect 11152 26910 11157 26962
rect 11157 26910 11204 26962
rect 11220 26910 11272 26962
rect 11288 26910 11335 26962
rect 11335 26910 11340 26962
rect 11152 26846 11157 26898
rect 11157 26846 11204 26898
rect 11220 26846 11272 26898
rect 11288 26846 11335 26898
rect 11335 26846 11340 26898
rect 11152 26782 11157 26834
rect 11157 26782 11204 26834
rect 11220 26782 11272 26834
rect 11288 26782 11335 26834
rect 11335 26782 11340 26834
rect 11152 26718 11157 26770
rect 11157 26718 11204 26770
rect 11220 26718 11272 26770
rect 11288 26718 11335 26770
rect 11335 26718 11340 26770
rect 11152 26654 11157 26706
rect 11157 26654 11204 26706
rect 11220 26654 11272 26706
rect 11288 26654 11335 26706
rect 11335 26654 11340 26706
rect 11152 26590 11157 26642
rect 11157 26590 11204 26642
rect 11220 26590 11272 26642
rect 11288 26590 11335 26642
rect 11335 26590 11340 26642
rect 11152 26526 11157 26578
rect 11157 26526 11204 26578
rect 11220 26526 11272 26578
rect 11288 26526 11335 26578
rect 11335 26526 11340 26578
rect 11152 26462 11157 26514
rect 11157 26462 11204 26514
rect 11220 26462 11272 26514
rect 11288 26462 11335 26514
rect 11335 26462 11340 26514
rect 11152 26398 11157 26450
rect 11157 26398 11204 26450
rect 11220 26398 11272 26450
rect 11288 26398 11335 26450
rect 11335 26398 11340 26450
rect 11152 26334 11157 26386
rect 11157 26334 11204 26386
rect 11220 26334 11272 26386
rect 11288 26334 11335 26386
rect 11335 26334 11340 26386
rect 11152 26270 11157 26322
rect 11157 26270 11204 26322
rect 11220 26270 11272 26322
rect 11288 26270 11335 26322
rect 11335 26270 11340 26322
rect 11152 26206 11157 26258
rect 11157 26206 11204 26258
rect 11220 26206 11272 26258
rect 11288 26206 11335 26258
rect 11335 26206 11340 26258
rect 11152 26142 11157 26194
rect 11157 26142 11204 26194
rect 11220 26142 11272 26194
rect 11288 26142 11335 26194
rect 11335 26142 11340 26194
rect 11152 26077 11157 26129
rect 11157 26077 11204 26129
rect 11220 26077 11272 26129
rect 11288 26077 11335 26129
rect 11335 26077 11340 26129
rect 11152 26012 11157 26064
rect 11157 26012 11204 26064
rect 11220 26012 11272 26064
rect 11288 26012 11335 26064
rect 11335 26012 11340 26064
rect 11152 25947 11157 25999
rect 11157 25947 11204 25999
rect 11220 25947 11272 25999
rect 11288 25947 11335 25999
rect 11335 25947 11340 25999
rect 11152 25882 11157 25934
rect 11157 25882 11204 25934
rect 11220 25882 11272 25934
rect 11288 25882 11335 25934
rect 11335 25882 11340 25934
rect 11152 25817 11157 25869
rect 11157 25817 11204 25869
rect 11220 25817 11272 25869
rect 11288 25817 11335 25869
rect 11335 25817 11340 25869
rect 11152 25752 11157 25804
rect 11157 25752 11204 25804
rect 11220 25752 11272 25804
rect 11288 25752 11335 25804
rect 11335 25752 11340 25804
rect 11152 25687 11157 25739
rect 11157 25687 11204 25739
rect 11220 25687 11272 25739
rect 11288 25687 11335 25739
rect 11335 25687 11340 25739
rect 11152 25622 11157 25674
rect 11157 25622 11204 25674
rect 11220 25622 11272 25674
rect 11288 25622 11335 25674
rect 11335 25622 11340 25674
rect 11152 25557 11157 25609
rect 11157 25557 11204 25609
rect 11220 25557 11272 25609
rect 11288 25557 11335 25609
rect 11335 25557 11340 25609
rect 11152 25492 11157 25544
rect 11157 25492 11204 25544
rect 11220 25492 11272 25544
rect 11288 25492 11335 25544
rect 11335 25492 11340 25544
rect 11152 25427 11157 25479
rect 11157 25427 11204 25479
rect 11220 25427 11272 25479
rect 11288 25427 11335 25479
rect 11335 25427 11340 25479
rect 11152 25362 11157 25414
rect 11157 25362 11204 25414
rect 11220 25362 11272 25414
rect 11288 25362 11335 25414
rect 11335 25362 11340 25414
rect 11152 22438 11157 22490
rect 11157 22438 11204 22490
rect 11220 22438 11272 22490
rect 11288 22438 11335 22490
rect 11335 22438 11340 22490
rect 11152 22374 11157 22426
rect 11157 22374 11204 22426
rect 11220 22374 11272 22426
rect 11288 22374 11335 22426
rect 11335 22374 11340 22426
rect 11152 22310 11157 22362
rect 11157 22310 11204 22362
rect 11220 22310 11272 22362
rect 11288 22310 11335 22362
rect 11335 22310 11340 22362
rect 11152 22246 11157 22298
rect 11157 22246 11204 22298
rect 11220 22246 11272 22298
rect 11288 22246 11335 22298
rect 11335 22246 11340 22298
rect 11152 22182 11157 22234
rect 11157 22182 11204 22234
rect 11220 22182 11272 22234
rect 11288 22182 11335 22234
rect 11335 22182 11340 22234
rect 11152 22118 11157 22170
rect 11157 22118 11204 22170
rect 11220 22118 11272 22170
rect 11288 22118 11335 22170
rect 11335 22118 11340 22170
rect 11152 22054 11157 22106
rect 11157 22054 11204 22106
rect 11220 22054 11272 22106
rect 11288 22054 11335 22106
rect 11335 22054 11340 22106
rect 11152 21990 11157 22042
rect 11157 21990 11204 22042
rect 11220 21990 11272 22042
rect 11288 21990 11335 22042
rect 11335 21990 11340 22042
rect 11152 21926 11157 21978
rect 11157 21926 11204 21978
rect 11220 21926 11272 21978
rect 11288 21926 11335 21978
rect 11335 21926 11340 21978
rect 11152 21862 11157 21914
rect 11157 21862 11204 21914
rect 11220 21862 11272 21914
rect 11288 21862 11335 21914
rect 11335 21862 11340 21914
rect 11152 21798 11157 21850
rect 11157 21798 11204 21850
rect 11220 21798 11272 21850
rect 11288 21798 11335 21850
rect 11335 21798 11340 21850
rect 11152 21734 11157 21786
rect 11157 21734 11204 21786
rect 11220 21734 11272 21786
rect 11288 21734 11335 21786
rect 11335 21734 11340 21786
rect 11152 21670 11157 21722
rect 11157 21670 11204 21722
rect 11220 21670 11272 21722
rect 11288 21670 11335 21722
rect 11335 21670 11340 21722
rect 11152 21606 11157 21658
rect 11157 21606 11204 21658
rect 11220 21606 11272 21658
rect 11288 21606 11335 21658
rect 11335 21606 11340 21658
rect 11152 21542 11157 21594
rect 11157 21542 11204 21594
rect 11220 21542 11272 21594
rect 11288 21542 11335 21594
rect 11335 21542 11340 21594
rect 11152 21477 11157 21529
rect 11157 21477 11204 21529
rect 11220 21477 11272 21529
rect 11288 21477 11335 21529
rect 11335 21477 11340 21529
rect 11152 21412 11157 21464
rect 11157 21412 11204 21464
rect 11220 21412 11272 21464
rect 11288 21412 11335 21464
rect 11335 21412 11340 21464
rect 11152 21347 11157 21399
rect 11157 21347 11204 21399
rect 11220 21347 11272 21399
rect 11288 21347 11335 21399
rect 11335 21347 11340 21399
rect 11152 21282 11157 21334
rect 11157 21282 11204 21334
rect 11220 21282 11272 21334
rect 11288 21282 11335 21334
rect 11335 21282 11340 21334
rect 11152 21217 11157 21269
rect 11157 21217 11204 21269
rect 11220 21217 11272 21269
rect 11288 21217 11335 21269
rect 11335 21217 11340 21269
rect 11152 21152 11157 21204
rect 11157 21152 11204 21204
rect 11220 21152 11272 21204
rect 11288 21152 11335 21204
rect 11335 21152 11340 21204
rect 11152 21087 11157 21139
rect 11157 21087 11204 21139
rect 11220 21087 11272 21139
rect 11288 21087 11335 21139
rect 11335 21087 11340 21139
rect 11152 21022 11157 21074
rect 11157 21022 11204 21074
rect 11220 21022 11272 21074
rect 11288 21022 11335 21074
rect 11335 21022 11340 21074
rect 11152 20957 11157 21009
rect 11157 20957 11204 21009
rect 11220 20957 11272 21009
rect 11288 20957 11335 21009
rect 11335 20957 11340 21009
rect 11152 20892 11157 20944
rect 11157 20892 11204 20944
rect 11220 20892 11272 20944
rect 11288 20892 11335 20944
rect 11335 20892 11340 20944
rect 11152 20827 11157 20879
rect 11157 20827 11204 20879
rect 11220 20827 11272 20879
rect 11288 20827 11335 20879
rect 11335 20827 11340 20879
rect 11152 20762 11157 20814
rect 11157 20762 11204 20814
rect 11220 20762 11272 20814
rect 11288 20762 11335 20814
rect 11335 20762 11340 20814
rect 11152 17838 11157 17890
rect 11157 17838 11204 17890
rect 11220 17838 11272 17890
rect 11288 17838 11335 17890
rect 11335 17838 11340 17890
rect 11152 17774 11157 17826
rect 11157 17774 11204 17826
rect 11220 17774 11272 17826
rect 11288 17774 11335 17826
rect 11335 17774 11340 17826
rect 11152 17710 11157 17762
rect 11157 17710 11204 17762
rect 11220 17710 11272 17762
rect 11288 17710 11335 17762
rect 11335 17710 11340 17762
rect 11152 17646 11157 17698
rect 11157 17646 11204 17698
rect 11220 17646 11272 17698
rect 11288 17646 11335 17698
rect 11335 17646 11340 17698
rect 11152 17582 11157 17634
rect 11157 17582 11204 17634
rect 11220 17582 11272 17634
rect 11288 17582 11335 17634
rect 11335 17582 11340 17634
rect 11152 17518 11157 17570
rect 11157 17518 11204 17570
rect 11220 17518 11272 17570
rect 11288 17518 11335 17570
rect 11335 17518 11340 17570
rect 11152 17454 11157 17506
rect 11157 17454 11204 17506
rect 11220 17454 11272 17506
rect 11288 17454 11335 17506
rect 11335 17454 11340 17506
rect 11152 17390 11157 17442
rect 11157 17390 11204 17442
rect 11220 17390 11272 17442
rect 11288 17390 11335 17442
rect 11335 17390 11340 17442
rect 11152 17326 11157 17378
rect 11157 17326 11204 17378
rect 11220 17326 11272 17378
rect 11288 17326 11335 17378
rect 11335 17326 11340 17378
rect 11152 17262 11157 17314
rect 11157 17262 11204 17314
rect 11220 17262 11272 17314
rect 11288 17262 11335 17314
rect 11335 17262 11340 17314
rect 11152 17198 11157 17250
rect 11157 17198 11204 17250
rect 11220 17198 11272 17250
rect 11288 17198 11335 17250
rect 11335 17198 11340 17250
rect 11152 17134 11157 17186
rect 11157 17134 11204 17186
rect 11220 17134 11272 17186
rect 11288 17134 11335 17186
rect 11335 17134 11340 17186
rect 11152 17070 11157 17122
rect 11157 17070 11204 17122
rect 11220 17070 11272 17122
rect 11288 17070 11335 17122
rect 11335 17070 11340 17122
rect 11152 17006 11157 17058
rect 11157 17006 11204 17058
rect 11220 17006 11272 17058
rect 11288 17006 11335 17058
rect 11335 17006 11340 17058
rect 11152 16942 11157 16994
rect 11157 16942 11204 16994
rect 11220 16942 11272 16994
rect 11288 16942 11335 16994
rect 11335 16942 11340 16994
rect 11152 16877 11157 16929
rect 11157 16877 11204 16929
rect 11220 16877 11272 16929
rect 11288 16877 11335 16929
rect 11335 16877 11340 16929
rect 11152 16812 11157 16864
rect 11157 16812 11204 16864
rect 11220 16812 11272 16864
rect 11288 16812 11335 16864
rect 11335 16812 11340 16864
rect 11152 16747 11157 16799
rect 11157 16747 11204 16799
rect 11220 16747 11272 16799
rect 11288 16747 11335 16799
rect 11335 16747 11340 16799
rect 11152 16682 11157 16734
rect 11157 16682 11204 16734
rect 11220 16682 11272 16734
rect 11288 16682 11335 16734
rect 11335 16682 11340 16734
rect 11152 16617 11157 16669
rect 11157 16617 11204 16669
rect 11220 16617 11272 16669
rect 11288 16617 11335 16669
rect 11335 16617 11340 16669
rect 11152 16552 11157 16604
rect 11157 16552 11204 16604
rect 11220 16552 11272 16604
rect 11288 16552 11335 16604
rect 11335 16552 11340 16604
rect 11152 16487 11157 16539
rect 11157 16487 11204 16539
rect 11220 16487 11272 16539
rect 11288 16487 11335 16539
rect 11335 16487 11340 16539
rect 11152 16422 11157 16474
rect 11157 16422 11204 16474
rect 11220 16422 11272 16474
rect 11288 16422 11335 16474
rect 11335 16422 11340 16474
rect 11152 16357 11157 16409
rect 11157 16357 11204 16409
rect 11220 16357 11272 16409
rect 11288 16357 11335 16409
rect 11335 16357 11340 16409
rect 11152 16292 11157 16344
rect 11157 16292 11204 16344
rect 11220 16292 11272 16344
rect 11288 16292 11335 16344
rect 11335 16292 11340 16344
rect 11152 16227 11157 16279
rect 11157 16227 11204 16279
rect 11220 16227 11272 16279
rect 11288 16227 11335 16279
rect 11335 16227 11340 16279
rect 11152 16162 11157 16214
rect 11157 16162 11204 16214
rect 11220 16162 11272 16214
rect 11288 16162 11335 16214
rect 11335 16162 11340 16214
rect 11152 13238 11157 13290
rect 11157 13238 11204 13290
rect 11220 13238 11272 13290
rect 11288 13238 11335 13290
rect 11335 13238 11340 13290
rect 11152 13174 11157 13226
rect 11157 13174 11204 13226
rect 11220 13174 11272 13226
rect 11288 13174 11335 13226
rect 11335 13174 11340 13226
rect 11152 13110 11157 13162
rect 11157 13110 11204 13162
rect 11220 13110 11272 13162
rect 11288 13110 11335 13162
rect 11335 13110 11340 13162
rect 11152 13046 11157 13098
rect 11157 13046 11204 13098
rect 11220 13046 11272 13098
rect 11288 13046 11335 13098
rect 11335 13046 11340 13098
rect 11152 12982 11157 13034
rect 11157 12982 11204 13034
rect 11220 12982 11272 13034
rect 11288 12982 11335 13034
rect 11335 12982 11340 13034
rect 11152 12918 11157 12970
rect 11157 12918 11204 12970
rect 11220 12918 11272 12970
rect 11288 12918 11335 12970
rect 11335 12918 11340 12970
rect 11152 12854 11157 12906
rect 11157 12854 11204 12906
rect 11220 12854 11272 12906
rect 11288 12854 11335 12906
rect 11335 12854 11340 12906
rect 11152 12790 11157 12842
rect 11157 12790 11204 12842
rect 11220 12790 11272 12842
rect 11288 12790 11335 12842
rect 11335 12790 11340 12842
rect 11152 12726 11157 12778
rect 11157 12726 11204 12778
rect 11220 12726 11272 12778
rect 11288 12726 11335 12778
rect 11335 12726 11340 12778
rect 11152 12662 11157 12714
rect 11157 12662 11204 12714
rect 11220 12662 11272 12714
rect 11288 12662 11335 12714
rect 11335 12662 11340 12714
rect 11152 12598 11157 12650
rect 11157 12598 11204 12650
rect 11220 12598 11272 12650
rect 11288 12598 11335 12650
rect 11335 12598 11340 12650
rect 11152 12534 11157 12586
rect 11157 12534 11204 12586
rect 11220 12534 11272 12586
rect 11288 12534 11335 12586
rect 11335 12534 11340 12586
rect 11152 12470 11157 12522
rect 11157 12470 11204 12522
rect 11220 12470 11272 12522
rect 11288 12470 11335 12522
rect 11335 12470 11340 12522
rect 11152 12406 11157 12458
rect 11157 12406 11204 12458
rect 11220 12406 11272 12458
rect 11288 12406 11335 12458
rect 11335 12406 11340 12458
rect 11152 12342 11157 12394
rect 11157 12342 11204 12394
rect 11220 12342 11272 12394
rect 11288 12342 11335 12394
rect 11335 12342 11340 12394
rect 11152 12277 11157 12329
rect 11157 12277 11204 12329
rect 11220 12277 11272 12329
rect 11288 12277 11335 12329
rect 11335 12277 11340 12329
rect 11152 12212 11157 12264
rect 11157 12212 11204 12264
rect 11220 12212 11272 12264
rect 11288 12212 11335 12264
rect 11335 12212 11340 12264
rect 11152 12147 11157 12199
rect 11157 12147 11204 12199
rect 11220 12147 11272 12199
rect 11288 12147 11335 12199
rect 11335 12147 11340 12199
rect 11152 12082 11157 12134
rect 11157 12082 11204 12134
rect 11220 12082 11272 12134
rect 11288 12082 11335 12134
rect 11335 12082 11340 12134
rect 11152 12017 11157 12069
rect 11157 12017 11204 12069
rect 11220 12017 11272 12069
rect 11288 12017 11335 12069
rect 11335 12017 11340 12069
rect 11152 11952 11157 12004
rect 11157 11952 11204 12004
rect 11220 11952 11272 12004
rect 11288 11952 11335 12004
rect 11335 11952 11340 12004
rect 11152 11887 11157 11939
rect 11157 11887 11204 11939
rect 11220 11887 11272 11939
rect 11288 11887 11335 11939
rect 11335 11887 11340 11939
rect 11152 11822 11157 11874
rect 11157 11822 11204 11874
rect 11220 11822 11272 11874
rect 11288 11822 11335 11874
rect 11335 11822 11340 11874
rect 11152 11757 11157 11809
rect 11157 11757 11204 11809
rect 11220 11757 11272 11809
rect 11288 11757 11335 11809
rect 11335 11757 11340 11809
rect 11152 11692 11157 11744
rect 11157 11692 11204 11744
rect 11220 11692 11272 11744
rect 11288 11692 11335 11744
rect 11335 11692 11340 11744
rect 11152 11627 11157 11679
rect 11157 11627 11204 11679
rect 11220 11627 11272 11679
rect 11288 11627 11335 11679
rect 11335 11627 11340 11679
rect 11152 11562 11157 11614
rect 11157 11562 11204 11614
rect 11220 11562 11272 11614
rect 11288 11562 11335 11614
rect 11335 11562 11340 11614
rect 11641 37945 11693 37997
rect 11719 37945 11771 37997
rect 11641 37877 11693 37929
rect 11719 37877 11771 37929
rect 11641 37809 11693 37861
rect 11719 37809 11771 37861
rect 11641 37741 11693 37793
rect 11719 37741 11771 37793
rect 11641 37673 11693 37725
rect 11719 37673 11771 37725
rect 11641 37605 11693 37657
rect 11719 37605 11771 37657
rect 11641 37537 11693 37589
rect 11719 37537 11771 37589
rect 11641 37469 11693 37521
rect 11719 37469 11771 37521
rect 11641 37401 11693 37453
rect 11719 37401 11771 37453
rect 11641 37333 11693 37385
rect 11719 37333 11771 37385
rect 11641 37266 11693 37318
rect 11719 37266 11771 37318
rect 11641 37199 11693 37251
rect 11719 37199 11771 37251
rect 11641 37132 11693 37184
rect 11719 37132 11771 37184
rect 11641 37065 11693 37117
rect 11719 37065 11771 37117
rect 11641 34173 11693 34225
rect 11719 34173 11771 34225
rect 11641 34109 11693 34161
rect 11719 34109 11771 34161
rect 11641 34045 11693 34097
rect 11719 34045 11771 34097
rect 11641 33981 11693 34033
rect 11719 33981 11771 34033
rect 11641 33917 11693 33969
rect 11719 33917 11771 33969
rect 11641 33853 11693 33905
rect 11719 33853 11771 33905
rect 11641 33789 11693 33841
rect 11719 33789 11771 33841
rect 11641 33725 11693 33777
rect 11719 33725 11771 33777
rect 11641 33661 11693 33713
rect 11719 33661 11771 33713
rect 11641 33597 11693 33649
rect 11719 33597 11771 33649
rect 11641 33533 11693 33585
rect 11719 33533 11771 33585
rect 11641 33469 11693 33521
rect 11719 33469 11771 33521
rect 11641 33405 11693 33457
rect 11719 33405 11771 33457
rect 11641 33341 11693 33393
rect 11719 33341 11771 33393
rect 11641 33277 11693 33329
rect 11719 33277 11771 33329
rect 11641 33212 11693 33264
rect 11719 33212 11771 33264
rect 11641 33147 11693 33199
rect 11719 33147 11771 33199
rect 11641 33082 11693 33134
rect 11719 33082 11771 33134
rect 11641 33017 11693 33069
rect 11719 33017 11771 33069
rect 11641 32952 11693 33004
rect 11719 32952 11771 33004
rect 11641 32887 11693 32939
rect 11719 32887 11771 32939
rect 11641 32822 11693 32874
rect 11719 32822 11771 32874
rect 11641 32757 11693 32809
rect 11719 32757 11771 32809
rect 11641 32692 11693 32744
rect 11719 32692 11771 32744
rect 11641 32627 11693 32679
rect 11719 32627 11771 32679
rect 11641 32562 11693 32614
rect 11719 32562 11771 32614
rect 11641 32497 11693 32549
rect 11719 32497 11771 32549
rect 11641 29573 11693 29625
rect 11719 29573 11771 29625
rect 11641 29509 11693 29561
rect 11719 29509 11771 29561
rect 11641 29445 11693 29497
rect 11719 29445 11771 29497
rect 11641 29381 11693 29433
rect 11719 29381 11771 29433
rect 11641 29317 11693 29369
rect 11719 29317 11771 29369
rect 11641 29253 11693 29305
rect 11719 29253 11771 29305
rect 11641 29189 11693 29241
rect 11719 29189 11771 29241
rect 11641 29125 11693 29177
rect 11719 29125 11771 29177
rect 11641 29061 11693 29113
rect 11719 29061 11771 29113
rect 11641 28997 11693 29049
rect 11719 28997 11771 29049
rect 11641 28933 11693 28985
rect 11719 28933 11771 28985
rect 11641 28869 11693 28921
rect 11719 28869 11771 28921
rect 11641 28805 11693 28857
rect 11719 28805 11771 28857
rect 11641 28741 11693 28793
rect 11719 28741 11771 28793
rect 11641 28677 11693 28729
rect 11719 28677 11771 28729
rect 11641 28612 11693 28664
rect 11719 28612 11771 28664
rect 11641 28547 11693 28599
rect 11719 28547 11771 28599
rect 11641 28482 11693 28534
rect 11719 28482 11771 28534
rect 11641 28417 11693 28469
rect 11719 28417 11771 28469
rect 11641 28352 11693 28404
rect 11719 28352 11771 28404
rect 11641 28287 11693 28339
rect 11719 28287 11771 28339
rect 11641 28222 11693 28274
rect 11719 28222 11771 28274
rect 11641 28157 11693 28209
rect 11719 28157 11771 28209
rect 11641 28092 11693 28144
rect 11719 28092 11771 28144
rect 11641 28027 11693 28079
rect 11719 28027 11771 28079
rect 11641 27962 11693 28014
rect 11719 27962 11771 28014
rect 11641 27897 11693 27949
rect 11719 27897 11771 27949
rect 11641 24973 11693 25025
rect 11719 24973 11771 25025
rect 11641 24909 11693 24961
rect 11719 24909 11771 24961
rect 11641 24845 11693 24897
rect 11719 24845 11771 24897
rect 11641 24781 11693 24833
rect 11719 24781 11771 24833
rect 11641 24717 11693 24769
rect 11719 24717 11771 24769
rect 11641 24653 11693 24705
rect 11719 24653 11771 24705
rect 11641 24589 11693 24641
rect 11719 24589 11771 24641
rect 11641 24525 11693 24577
rect 11719 24525 11771 24577
rect 11641 24461 11693 24513
rect 11719 24461 11771 24513
rect 11641 24397 11693 24449
rect 11719 24397 11771 24449
rect 11641 24333 11693 24385
rect 11719 24333 11771 24385
rect 11641 24269 11693 24321
rect 11719 24269 11771 24321
rect 11641 24205 11693 24257
rect 11719 24205 11771 24257
rect 11641 24141 11693 24193
rect 11719 24141 11771 24193
rect 11641 24077 11693 24129
rect 11719 24077 11771 24129
rect 11641 24012 11693 24064
rect 11719 24012 11771 24064
rect 11641 23947 11693 23999
rect 11719 23947 11771 23999
rect 11641 23882 11693 23934
rect 11719 23882 11771 23934
rect 11641 23817 11693 23869
rect 11719 23817 11771 23869
rect 11641 23752 11693 23804
rect 11719 23752 11771 23804
rect 11641 23687 11693 23739
rect 11719 23687 11771 23739
rect 11641 23622 11693 23674
rect 11719 23622 11771 23674
rect 11641 23557 11693 23609
rect 11719 23557 11771 23609
rect 11641 23492 11693 23544
rect 11719 23492 11771 23544
rect 11641 23427 11693 23479
rect 11719 23427 11771 23479
rect 11641 23362 11693 23414
rect 11719 23362 11771 23414
rect 11641 23297 11693 23349
rect 11719 23297 11771 23349
rect 11641 20373 11693 20425
rect 11719 20373 11771 20425
rect 11641 20309 11693 20361
rect 11719 20309 11771 20361
rect 11641 20245 11693 20297
rect 11719 20245 11771 20297
rect 11641 20181 11693 20233
rect 11719 20181 11771 20233
rect 11641 20117 11693 20169
rect 11719 20117 11771 20169
rect 11641 20053 11693 20105
rect 11719 20053 11771 20105
rect 11641 19989 11693 20041
rect 11719 19989 11771 20041
rect 11641 19925 11693 19977
rect 11719 19925 11771 19977
rect 11641 19861 11693 19913
rect 11719 19861 11771 19913
rect 11641 19797 11693 19849
rect 11719 19797 11771 19849
rect 11641 19733 11693 19785
rect 11719 19733 11771 19785
rect 11641 19669 11693 19721
rect 11719 19669 11771 19721
rect 11641 19605 11693 19657
rect 11719 19605 11771 19657
rect 11641 19541 11693 19593
rect 11719 19541 11771 19593
rect 11641 19477 11693 19529
rect 11719 19477 11771 19529
rect 11641 19412 11693 19464
rect 11719 19412 11771 19464
rect 11641 19347 11693 19399
rect 11719 19347 11771 19399
rect 11641 19282 11693 19334
rect 11719 19282 11771 19334
rect 11641 19217 11693 19269
rect 11719 19217 11771 19269
rect 11641 19152 11693 19204
rect 11719 19152 11771 19204
rect 11641 19087 11693 19139
rect 11719 19087 11771 19139
rect 11641 19022 11693 19074
rect 11719 19022 11771 19074
rect 11641 18957 11693 19009
rect 11719 18957 11771 19009
rect 11641 18892 11693 18944
rect 11719 18892 11771 18944
rect 11641 18827 11693 18879
rect 11719 18827 11771 18879
rect 11641 18762 11693 18814
rect 11719 18762 11771 18814
rect 11641 18697 11693 18749
rect 11719 18697 11771 18749
rect 11641 15773 11693 15825
rect 11719 15773 11771 15825
rect 11641 15709 11693 15761
rect 11719 15709 11771 15761
rect 11641 15645 11693 15697
rect 11719 15645 11771 15697
rect 11641 15581 11693 15633
rect 11719 15581 11771 15633
rect 11641 15517 11693 15569
rect 11719 15517 11771 15569
rect 11641 15453 11693 15505
rect 11719 15453 11771 15505
rect 11641 15389 11693 15441
rect 11719 15389 11771 15441
rect 11641 15325 11693 15377
rect 11719 15325 11771 15377
rect 11641 15261 11693 15313
rect 11719 15261 11771 15313
rect 11641 15197 11693 15249
rect 11719 15197 11771 15249
rect 11641 15133 11693 15185
rect 11719 15133 11771 15185
rect 11641 15069 11693 15121
rect 11719 15069 11771 15121
rect 11641 15005 11693 15057
rect 11719 15005 11771 15057
rect 11641 14941 11693 14993
rect 11719 14941 11771 14993
rect 11641 14877 11693 14929
rect 11719 14877 11771 14929
rect 11641 14812 11693 14864
rect 11719 14812 11771 14864
rect 11641 14747 11693 14799
rect 11719 14747 11771 14799
rect 11641 14682 11693 14734
rect 11719 14682 11771 14734
rect 11641 14617 11693 14669
rect 11719 14617 11771 14669
rect 11641 14552 11693 14604
rect 11719 14552 11771 14604
rect 11641 14487 11693 14539
rect 11719 14487 11771 14539
rect 11641 14422 11693 14474
rect 11719 14422 11771 14474
rect 11641 14357 11693 14409
rect 11719 14357 11771 14409
rect 11641 14292 11693 14344
rect 11719 14292 11771 14344
rect 11641 14227 11693 14279
rect 11719 14227 11771 14279
rect 11641 14162 11693 14214
rect 11719 14162 11771 14214
rect 11641 14097 11693 14149
rect 11719 14097 11771 14149
rect 11641 11173 11693 11225
rect 11719 11173 11771 11225
rect 11641 11109 11693 11161
rect 11719 11109 11771 11161
rect 11641 11045 11693 11097
rect 11719 11045 11771 11097
rect 11641 10981 11693 11033
rect 11719 10981 11771 11033
rect 11641 10917 11693 10969
rect 11719 10917 11771 10969
rect 11641 10853 11693 10905
rect 11719 10853 11771 10905
rect 11641 10789 11693 10841
rect 11719 10789 11771 10841
rect 11641 10725 11693 10777
rect 11719 10725 11771 10777
rect 11641 10661 11693 10713
rect 11719 10661 11771 10713
rect 11641 10597 11693 10649
rect 11719 10597 11771 10649
rect 11641 10533 11693 10585
rect 11719 10533 11771 10585
rect 11641 10469 11693 10521
rect 11719 10469 11771 10521
rect 11641 10405 11693 10457
rect 11719 10405 11771 10457
rect 11641 10341 11693 10393
rect 11719 10341 11771 10393
rect 11641 10277 11693 10329
rect 11719 10277 11771 10329
rect 11641 10212 11693 10264
rect 11719 10212 11771 10264
rect 11641 10147 11693 10199
rect 11719 10147 11771 10199
rect 11641 10082 11693 10134
rect 11719 10082 11771 10134
rect 11641 10017 11693 10069
rect 11719 10017 11771 10069
rect 11641 9952 11693 10004
rect 11719 9952 11771 10004
rect 11641 9887 11693 9939
rect 11719 9887 11771 9939
rect 11641 9822 11693 9874
rect 11719 9822 11771 9874
rect 11641 9757 11693 9809
rect 11719 9757 11771 9809
rect 11641 9692 11693 9744
rect 11719 9692 11771 9744
rect 11641 9627 11693 9679
rect 11719 9627 11771 9679
rect 11641 9562 11693 9614
rect 11719 9562 11771 9614
rect 11641 9497 11693 9549
rect 11719 9497 11771 9549
rect 12992 38957 12997 39009
rect 12997 38957 13044 39009
rect 13060 38957 13112 39009
rect 13128 38957 13175 39009
rect 13175 38957 13180 39009
rect 12992 38893 12997 38945
rect 12997 38893 13044 38945
rect 13060 38893 13112 38945
rect 13128 38893 13175 38945
rect 13175 38893 13180 38945
rect 12992 38829 12997 38881
rect 12997 38829 13044 38881
rect 13060 38829 13112 38881
rect 13128 38829 13175 38881
rect 13175 38829 13180 38881
rect 12992 38765 12997 38817
rect 12997 38765 13044 38817
rect 13060 38765 13112 38817
rect 13128 38765 13175 38817
rect 13175 38765 13180 38817
rect 12992 38701 12997 38753
rect 12997 38701 13044 38753
rect 13060 38701 13112 38753
rect 13128 38701 13175 38753
rect 13175 38701 13180 38753
rect 12992 38637 12997 38689
rect 12997 38637 13044 38689
rect 13060 38637 13112 38689
rect 13128 38637 13175 38689
rect 13175 38637 13180 38689
rect 12992 38573 12997 38625
rect 12997 38573 13044 38625
rect 13060 38573 13112 38625
rect 13128 38573 13175 38625
rect 13175 38573 13180 38625
rect 12992 38508 12997 38560
rect 12997 38508 13044 38560
rect 13060 38508 13112 38560
rect 13128 38508 13175 38560
rect 13175 38508 13180 38560
rect 12992 38490 12997 38495
rect 12997 38490 13044 38495
rect 13060 38490 13112 38495
rect 13128 38490 13175 38495
rect 13175 38490 13180 38495
rect 12992 38451 13044 38490
rect 12992 38443 12997 38451
rect 12997 38443 13031 38451
rect 13031 38443 13044 38451
rect 13060 38451 13112 38490
rect 13060 38443 13069 38451
rect 13069 38443 13103 38451
rect 13103 38443 13112 38451
rect 13128 38451 13180 38490
rect 13128 38443 13141 38451
rect 13141 38443 13175 38451
rect 13175 38443 13180 38451
rect 12992 38417 12997 38430
rect 12997 38417 13031 38430
rect 13031 38417 13044 38430
rect 12992 38378 13044 38417
rect 13060 38417 13069 38430
rect 13069 38417 13103 38430
rect 13103 38417 13112 38430
rect 13060 38378 13112 38417
rect 13128 38417 13141 38430
rect 13141 38417 13175 38430
rect 13175 38417 13180 38430
rect 13128 38378 13180 38417
rect 12992 38344 12997 38365
rect 12997 38344 13031 38365
rect 13031 38344 13044 38365
rect 12992 38313 13044 38344
rect 13060 38344 13069 38365
rect 13069 38344 13103 38365
rect 13103 38344 13112 38365
rect 13060 38313 13112 38344
rect 13128 38344 13141 38365
rect 13141 38344 13175 38365
rect 13175 38344 13180 38365
rect 13128 38313 13180 38344
rect 12992 38271 12997 38300
rect 12997 38271 13031 38300
rect 13031 38271 13044 38300
rect 12992 38248 13044 38271
rect 13060 38271 13069 38300
rect 13069 38271 13103 38300
rect 13103 38271 13112 38300
rect 13060 38248 13112 38271
rect 13128 38271 13141 38300
rect 13141 38271 13175 38300
rect 13175 38271 13180 38300
rect 13128 38248 13180 38271
rect 12992 38232 13044 38235
rect 12992 38198 12997 38232
rect 12997 38198 13031 38232
rect 13031 38198 13044 38232
rect 12992 38183 13044 38198
rect 13060 38232 13112 38235
rect 13060 38198 13069 38232
rect 13069 38198 13103 38232
rect 13103 38198 13112 38232
rect 13060 38183 13112 38198
rect 13128 38232 13180 38235
rect 13128 38198 13141 38232
rect 13141 38198 13175 38232
rect 13175 38198 13180 38232
rect 13128 38183 13180 38198
rect 12992 38159 13044 38170
rect 12992 38125 12997 38159
rect 12997 38125 13031 38159
rect 13031 38125 13044 38159
rect 12992 38118 13044 38125
rect 13060 38159 13112 38170
rect 13060 38125 13069 38159
rect 13069 38125 13103 38159
rect 13103 38125 13112 38159
rect 13060 38118 13112 38125
rect 13128 38159 13180 38170
rect 13128 38125 13141 38159
rect 13141 38125 13175 38159
rect 13175 38125 13180 38159
rect 13128 38118 13180 38125
rect 12561 37945 12613 37997
rect 12639 37945 12691 37997
rect 12561 37877 12613 37929
rect 12639 37877 12691 37929
rect 12561 37809 12613 37861
rect 12639 37809 12691 37861
rect 12561 37741 12613 37793
rect 12639 37741 12691 37793
rect 12561 37673 12613 37725
rect 12639 37673 12691 37725
rect 12561 37605 12613 37657
rect 12639 37605 12691 37657
rect 12561 37537 12613 37589
rect 12639 37537 12691 37589
rect 12561 37469 12613 37521
rect 12639 37469 12691 37521
rect 12561 37401 12613 37453
rect 12639 37401 12691 37453
rect 12561 37333 12613 37385
rect 12639 37333 12691 37385
rect 12561 37266 12613 37318
rect 12639 37266 12691 37318
rect 12561 37199 12613 37251
rect 12639 37199 12691 37251
rect 12561 37132 12613 37184
rect 12639 37132 12691 37184
rect 12561 37065 12613 37117
rect 12639 37065 12691 37117
rect 12561 34173 12613 34225
rect 12639 34173 12691 34225
rect 12561 34109 12613 34161
rect 12639 34109 12691 34161
rect 12561 34045 12613 34097
rect 12639 34045 12691 34097
rect 12561 33981 12613 34033
rect 12639 33981 12691 34033
rect 12561 33917 12613 33969
rect 12639 33917 12691 33969
rect 12561 33853 12613 33905
rect 12639 33853 12691 33905
rect 12561 33789 12613 33841
rect 12639 33789 12691 33841
rect 12561 33725 12613 33777
rect 12639 33725 12691 33777
rect 12561 33661 12613 33713
rect 12639 33661 12691 33713
rect 12561 33597 12613 33649
rect 12639 33597 12691 33649
rect 12561 33533 12613 33585
rect 12639 33533 12691 33585
rect 12561 33469 12613 33521
rect 12639 33469 12691 33521
rect 12561 33405 12613 33457
rect 12639 33405 12691 33457
rect 12561 33341 12613 33393
rect 12639 33341 12691 33393
rect 12561 33277 12613 33329
rect 12639 33277 12691 33329
rect 12561 33212 12613 33264
rect 12639 33212 12691 33264
rect 12561 33147 12613 33199
rect 12639 33147 12691 33199
rect 12561 33082 12613 33134
rect 12639 33082 12691 33134
rect 12561 33017 12613 33069
rect 12639 33017 12691 33069
rect 12561 32952 12613 33004
rect 12639 32952 12691 33004
rect 12561 32887 12613 32939
rect 12639 32887 12691 32939
rect 12561 32822 12613 32874
rect 12639 32822 12691 32874
rect 12561 32757 12613 32809
rect 12639 32757 12691 32809
rect 12561 32692 12613 32744
rect 12639 32692 12691 32744
rect 12561 32627 12613 32679
rect 12639 32627 12691 32679
rect 12561 32562 12613 32614
rect 12639 32562 12691 32614
rect 12561 32497 12613 32549
rect 12639 32497 12691 32549
rect 12561 29573 12613 29625
rect 12639 29573 12691 29625
rect 12561 29509 12613 29561
rect 12639 29509 12691 29561
rect 12561 29445 12613 29497
rect 12639 29445 12691 29497
rect 12561 29381 12613 29433
rect 12639 29381 12691 29433
rect 12561 29317 12613 29369
rect 12639 29317 12691 29369
rect 12561 29253 12613 29305
rect 12639 29253 12691 29305
rect 12561 29189 12613 29241
rect 12639 29189 12691 29241
rect 12561 29125 12613 29177
rect 12639 29125 12691 29177
rect 12561 29061 12613 29113
rect 12639 29061 12691 29113
rect 12561 28997 12613 29049
rect 12639 28997 12691 29049
rect 12561 28933 12613 28985
rect 12639 28933 12691 28985
rect 12561 28869 12613 28921
rect 12639 28869 12691 28921
rect 12561 28805 12613 28857
rect 12639 28805 12691 28857
rect 12561 28741 12613 28793
rect 12639 28741 12691 28793
rect 12561 28677 12613 28729
rect 12639 28677 12691 28729
rect 12561 28612 12613 28664
rect 12639 28612 12691 28664
rect 12561 28547 12613 28599
rect 12639 28547 12691 28599
rect 12561 28482 12613 28534
rect 12639 28482 12691 28534
rect 12561 28417 12613 28469
rect 12639 28417 12691 28469
rect 12561 28352 12613 28404
rect 12639 28352 12691 28404
rect 12561 28287 12613 28339
rect 12639 28287 12691 28339
rect 12561 28222 12613 28274
rect 12639 28222 12691 28274
rect 12561 28157 12613 28209
rect 12639 28157 12691 28209
rect 12561 28092 12613 28144
rect 12639 28092 12691 28144
rect 12561 28027 12613 28079
rect 12639 28027 12691 28079
rect 12561 27962 12613 28014
rect 12639 27962 12691 28014
rect 12561 27897 12613 27949
rect 12639 27897 12691 27949
rect 12561 24973 12613 25025
rect 12639 24973 12691 25025
rect 12561 24909 12613 24961
rect 12639 24909 12691 24961
rect 12561 24845 12613 24897
rect 12639 24845 12691 24897
rect 12561 24781 12613 24833
rect 12639 24781 12691 24833
rect 12561 24717 12613 24769
rect 12639 24717 12691 24769
rect 12561 24653 12613 24705
rect 12639 24653 12691 24705
rect 12561 24589 12613 24641
rect 12639 24589 12691 24641
rect 12561 24525 12613 24577
rect 12639 24525 12691 24577
rect 12561 24461 12613 24513
rect 12639 24461 12691 24513
rect 12561 24397 12613 24449
rect 12639 24397 12691 24449
rect 12561 24333 12613 24385
rect 12639 24333 12691 24385
rect 12561 24269 12613 24321
rect 12639 24269 12691 24321
rect 12561 24205 12613 24257
rect 12639 24205 12691 24257
rect 12561 24141 12613 24193
rect 12639 24141 12691 24193
rect 12561 24077 12613 24129
rect 12639 24077 12691 24129
rect 12561 24012 12613 24064
rect 12639 24012 12691 24064
rect 12561 23947 12613 23999
rect 12639 23947 12691 23999
rect 12561 23882 12613 23934
rect 12639 23882 12691 23934
rect 12561 23817 12613 23869
rect 12639 23817 12691 23869
rect 12561 23752 12613 23804
rect 12639 23752 12691 23804
rect 12561 23687 12613 23739
rect 12639 23687 12691 23739
rect 12561 23622 12613 23674
rect 12639 23622 12691 23674
rect 12561 23557 12613 23609
rect 12639 23557 12691 23609
rect 12561 23492 12613 23544
rect 12639 23492 12691 23544
rect 12561 23427 12613 23479
rect 12639 23427 12691 23479
rect 12561 23362 12613 23414
rect 12639 23362 12691 23414
rect 12561 23297 12613 23349
rect 12639 23297 12691 23349
rect 12561 20373 12613 20425
rect 12639 20373 12691 20425
rect 12561 20309 12613 20361
rect 12639 20309 12691 20361
rect 12561 20245 12613 20297
rect 12639 20245 12691 20297
rect 12561 20181 12613 20233
rect 12639 20181 12691 20233
rect 12561 20117 12613 20169
rect 12639 20117 12691 20169
rect 12561 20053 12613 20105
rect 12639 20053 12691 20105
rect 12561 19989 12613 20041
rect 12639 19989 12691 20041
rect 12561 19925 12613 19977
rect 12639 19925 12691 19977
rect 12561 19861 12613 19913
rect 12639 19861 12691 19913
rect 12561 19797 12613 19849
rect 12639 19797 12691 19849
rect 12561 19733 12613 19785
rect 12639 19733 12691 19785
rect 12561 19669 12613 19721
rect 12639 19669 12691 19721
rect 12561 19605 12613 19657
rect 12639 19605 12691 19657
rect 12561 19541 12613 19593
rect 12639 19541 12691 19593
rect 12561 19477 12613 19529
rect 12639 19477 12691 19529
rect 12561 19412 12613 19464
rect 12639 19412 12691 19464
rect 12561 19347 12613 19399
rect 12639 19347 12691 19399
rect 12561 19282 12613 19334
rect 12639 19282 12691 19334
rect 12561 19217 12613 19269
rect 12639 19217 12691 19269
rect 12561 19152 12613 19204
rect 12639 19152 12691 19204
rect 12561 19087 12613 19139
rect 12639 19087 12691 19139
rect 12561 19022 12613 19074
rect 12639 19022 12691 19074
rect 12561 18957 12613 19009
rect 12639 18957 12691 19009
rect 12561 18892 12613 18944
rect 12639 18892 12691 18944
rect 12561 18827 12613 18879
rect 12639 18827 12691 18879
rect 12561 18762 12613 18814
rect 12639 18762 12691 18814
rect 12561 18697 12613 18749
rect 12639 18697 12691 18749
rect 12561 15773 12613 15825
rect 12639 15773 12691 15825
rect 12561 15709 12613 15761
rect 12639 15709 12691 15761
rect 12561 15645 12613 15697
rect 12639 15645 12691 15697
rect 12561 15581 12613 15633
rect 12639 15581 12691 15633
rect 12561 15517 12613 15569
rect 12639 15517 12691 15569
rect 12561 15453 12613 15505
rect 12639 15453 12691 15505
rect 12561 15389 12613 15441
rect 12639 15389 12691 15441
rect 12561 15325 12613 15377
rect 12639 15325 12691 15377
rect 12561 15261 12613 15313
rect 12639 15261 12691 15313
rect 12561 15197 12613 15249
rect 12639 15197 12691 15249
rect 12561 15133 12613 15185
rect 12639 15133 12691 15185
rect 12561 15069 12613 15121
rect 12639 15069 12691 15121
rect 12561 15005 12613 15057
rect 12639 15005 12691 15057
rect 12561 14941 12613 14993
rect 12639 14941 12691 14993
rect 12561 14877 12613 14929
rect 12639 14877 12691 14929
rect 12561 14812 12613 14864
rect 12639 14812 12691 14864
rect 12561 14747 12613 14799
rect 12639 14747 12691 14799
rect 12561 14682 12613 14734
rect 12639 14682 12691 14734
rect 12561 14617 12613 14669
rect 12639 14617 12691 14669
rect 12561 14552 12613 14604
rect 12639 14552 12691 14604
rect 12561 14487 12613 14539
rect 12639 14487 12691 14539
rect 12561 14422 12613 14474
rect 12639 14422 12691 14474
rect 12561 14357 12613 14409
rect 12639 14357 12691 14409
rect 12561 14292 12613 14344
rect 12639 14292 12691 14344
rect 12561 14227 12613 14279
rect 12639 14227 12691 14279
rect 12561 14162 12613 14214
rect 12639 14162 12691 14214
rect 12561 14097 12613 14149
rect 12639 14097 12691 14149
rect 12561 11173 12613 11225
rect 12639 11173 12691 11225
rect 12561 11109 12613 11161
rect 12639 11109 12691 11161
rect 12561 11045 12613 11097
rect 12639 11045 12691 11097
rect 12561 10981 12613 11033
rect 12639 10981 12691 11033
rect 12561 10917 12613 10969
rect 12639 10917 12691 10969
rect 12561 10853 12613 10905
rect 12639 10853 12691 10905
rect 12561 10789 12613 10841
rect 12639 10789 12691 10841
rect 12561 10725 12613 10777
rect 12639 10725 12691 10777
rect 12561 10661 12613 10713
rect 12639 10661 12691 10713
rect 12561 10597 12613 10649
rect 12639 10597 12691 10649
rect 12561 10533 12613 10585
rect 12639 10533 12691 10585
rect 12561 10469 12613 10521
rect 12639 10469 12691 10521
rect 12561 10405 12613 10457
rect 12639 10405 12691 10457
rect 12561 10341 12613 10393
rect 12639 10341 12691 10393
rect 12561 10277 12613 10329
rect 12639 10277 12691 10329
rect 12561 10212 12613 10264
rect 12639 10212 12691 10264
rect 12561 10147 12613 10199
rect 12639 10147 12691 10199
rect 12561 10082 12613 10134
rect 12639 10082 12691 10134
rect 12561 10017 12613 10069
rect 12639 10017 12691 10069
rect 12561 9952 12613 10004
rect 12639 9952 12691 10004
rect 12561 9887 12613 9939
rect 12639 9887 12691 9939
rect 12561 9822 12613 9874
rect 12639 9822 12691 9874
rect 12561 9757 12613 9809
rect 12639 9757 12691 9809
rect 12561 9692 12613 9744
rect 12639 9692 12691 9744
rect 12561 9627 12613 9679
rect 12639 9627 12691 9679
rect 12561 9562 12613 9614
rect 12639 9562 12691 9614
rect 12561 9497 12613 9549
rect 12639 9497 12691 9549
rect 2233 9344 2285 9352
rect 2233 9310 2255 9344
rect 2255 9310 2285 9344
rect 2335 9343 2387 9352
rect 2233 9300 2285 9310
rect 2335 9309 2365 9343
rect 2365 9309 2387 9343
rect 2335 9300 2387 9309
rect 2233 9271 2285 9287
rect 2233 9237 2255 9271
rect 2255 9237 2285 9271
rect 2335 9270 2387 9287
rect 2233 9235 2285 9237
rect 2335 9235 2365 9270
rect 2365 9235 2387 9270
rect 2233 9198 2285 9222
rect 2335 9198 2365 9222
rect 2365 9198 2387 9222
rect 2233 9170 2255 9198
rect 2255 9170 2285 9198
rect 2335 9170 2387 9198
rect 2233 9105 2285 9157
rect 2335 9105 2387 9157
rect 11204 8879 11256 8881
rect 11204 8845 11219 8879
rect 11219 8845 11253 8879
rect 11253 8845 11256 8879
rect 11204 8829 11256 8845
rect 11274 8879 11326 8881
rect 11274 8845 11292 8879
rect 11292 8845 11326 8879
rect 11274 8829 11326 8845
rect 11344 8879 11396 8881
rect 11414 8879 11466 8881
rect 11483 8879 11535 8881
rect 11552 8879 11604 8881
rect 11621 8879 11673 8881
rect 11690 8879 11742 8881
rect 11759 8879 11811 8881
rect 11828 8879 11880 8881
rect 11897 8879 11949 8881
rect 11344 8845 11365 8879
rect 11365 8845 11396 8879
rect 11414 8845 11438 8879
rect 11438 8845 11466 8879
rect 11483 8845 11511 8879
rect 11511 8845 11535 8879
rect 11552 8845 11584 8879
rect 11584 8845 11604 8879
rect 11621 8845 11657 8879
rect 11657 8845 11673 8879
rect 11690 8845 11691 8879
rect 11691 8845 11730 8879
rect 11730 8845 11742 8879
rect 11759 8845 11764 8879
rect 11764 8845 11803 8879
rect 11803 8845 11811 8879
rect 11828 8845 11837 8879
rect 11837 8845 11876 8879
rect 11876 8845 11880 8879
rect 11897 8845 11910 8879
rect 11910 8845 11949 8879
rect 11344 8829 11396 8845
rect 11414 8829 11466 8845
rect 11483 8829 11535 8845
rect 11552 8829 11604 8845
rect 11621 8829 11673 8845
rect 11690 8829 11742 8845
rect 11759 8829 11811 8845
rect 11828 8829 11880 8845
rect 11897 8829 11949 8845
rect 11204 8735 11256 8759
rect 11204 8707 11218 8735
rect 11218 8707 11252 8735
rect 11252 8707 11256 8735
rect 11274 8735 11326 8759
rect 11274 8707 11291 8735
rect 11291 8707 11325 8735
rect 11325 8707 11326 8735
rect 11344 8735 11396 8759
rect 11414 8735 11466 8759
rect 11483 8735 11535 8759
rect 11552 8735 11604 8759
rect 11621 8735 11673 8759
rect 11690 8735 11742 8759
rect 11759 8735 11811 8759
rect 11828 8735 11880 8759
rect 11897 8735 11949 8759
rect 11344 8707 11364 8735
rect 11364 8707 11396 8735
rect 11414 8707 11437 8735
rect 11437 8707 11466 8735
rect 11483 8707 11510 8735
rect 11510 8707 11535 8735
rect 11552 8707 11583 8735
rect 11583 8707 11604 8735
rect 11621 8707 11656 8735
rect 11656 8707 11673 8735
rect 11690 8707 11729 8735
rect 11729 8707 11742 8735
rect 11759 8707 11763 8735
rect 11763 8707 11802 8735
rect 11802 8707 11811 8735
rect 11828 8707 11836 8735
rect 11836 8707 11875 8735
rect 11875 8707 11880 8735
rect 11897 8707 11909 8735
rect 11909 8707 11948 8735
rect 11948 8707 11949 8735
rect 11204 8465 11227 8495
rect 11227 8465 11256 8495
rect 11274 8465 11300 8495
rect 11300 8465 11326 8495
rect 11344 8465 11373 8495
rect 11373 8465 11396 8495
rect 11414 8465 11446 8495
rect 11446 8465 11466 8495
rect 11204 8443 11256 8465
rect 11274 8443 11326 8465
rect 11344 8443 11396 8465
rect 11414 8443 11466 8465
rect 11483 8465 11485 8495
rect 11485 8465 11519 8495
rect 11519 8465 11535 8495
rect 11483 8443 11535 8465
rect 11552 8465 11558 8495
rect 11558 8465 11592 8495
rect 11592 8465 11604 8495
rect 11552 8443 11604 8465
rect 11621 8465 11631 8495
rect 11631 8465 11665 8495
rect 11665 8465 11673 8495
rect 11621 8443 11673 8465
rect 11690 8465 11704 8495
rect 11704 8465 11738 8495
rect 11738 8465 11742 8495
rect 11690 8443 11742 8465
rect 11759 8465 11777 8495
rect 11777 8465 11811 8495
rect 11759 8443 11811 8465
rect 11828 8465 11850 8495
rect 11850 8465 11880 8495
rect 11897 8465 11923 8495
rect 11923 8465 11949 8495
rect 11828 8443 11880 8465
rect 11897 8443 11949 8465
rect 11204 8355 11256 8373
rect 11274 8355 11326 8373
rect 11344 8355 11396 8373
rect 11414 8355 11466 8373
rect 11204 8321 11226 8355
rect 11226 8321 11256 8355
rect 11274 8321 11299 8355
rect 11299 8321 11326 8355
rect 11344 8321 11372 8355
rect 11372 8321 11396 8355
rect 11414 8321 11445 8355
rect 11445 8321 11466 8355
rect 11483 8355 11535 8373
rect 11483 8321 11484 8355
rect 11484 8321 11518 8355
rect 11518 8321 11535 8355
rect 11552 8355 11604 8373
rect 11552 8321 11557 8355
rect 11557 8321 11591 8355
rect 11591 8321 11604 8355
rect 11621 8355 11673 8373
rect 11621 8321 11630 8355
rect 11630 8321 11664 8355
rect 11664 8321 11673 8355
rect 11690 8355 11742 8373
rect 11690 8321 11703 8355
rect 11703 8321 11737 8355
rect 11737 8321 11742 8355
rect 11759 8355 11811 8373
rect 11759 8321 11776 8355
rect 11776 8321 11810 8355
rect 11810 8321 11811 8355
rect 11828 8355 11880 8373
rect 11897 8355 11949 8373
rect 11828 8321 11849 8355
rect 11849 8321 11880 8355
rect 11897 8321 11922 8355
rect 11922 8321 11949 8355
rect 695 7883 698 7914
rect 698 7883 732 7914
rect 732 7883 747 7914
rect 695 7862 747 7883
rect 761 7883 771 7914
rect 771 7883 805 7914
rect 805 7883 813 7914
rect 761 7862 813 7883
rect 827 7883 844 7914
rect 844 7883 878 7914
rect 878 7883 879 7914
rect 827 7862 879 7883
rect 893 7883 917 7914
rect 917 7883 945 7914
rect 959 7883 990 7914
rect 990 7883 1011 7914
rect 1025 7883 1063 7914
rect 1063 7883 1077 7914
rect 1091 7883 1097 7914
rect 1097 7883 1136 7914
rect 1136 7883 1143 7914
rect 1157 7883 1170 7914
rect 1170 7883 1209 7914
rect 1223 7883 1243 7914
rect 1243 7883 1275 7914
rect 1289 7883 1316 7914
rect 1316 7883 1341 7914
rect 893 7862 945 7883
rect 959 7862 1011 7883
rect 1025 7862 1077 7883
rect 1091 7862 1143 7883
rect 1157 7862 1209 7883
rect 1223 7862 1275 7883
rect 1289 7862 1341 7883
rect 1355 7883 1389 7914
rect 1389 7883 1407 7914
rect 1355 7862 1407 7883
rect 1421 7883 1428 7914
rect 1428 7883 1462 7914
rect 1462 7883 1473 7914
rect 1421 7862 1473 7883
rect 1487 7883 1501 7914
rect 1501 7883 1535 7914
rect 1535 7883 1539 7914
rect 1487 7862 1539 7883
rect 1553 7883 1574 7914
rect 1574 7883 1605 7914
rect 1619 7883 1647 7914
rect 1647 7883 1671 7914
rect 1684 7883 1720 7914
rect 1720 7883 1736 7914
rect 1749 7883 1754 7914
rect 1754 7883 1793 7914
rect 1793 7883 1801 7914
rect 1814 7883 1827 7914
rect 1827 7883 1866 7914
rect 1879 7883 1900 7914
rect 1900 7883 1931 7914
rect 1944 7883 1973 7914
rect 1973 7883 1996 7914
rect 1553 7862 1605 7883
rect 1619 7862 1671 7883
rect 1684 7862 1736 7883
rect 1749 7862 1801 7883
rect 1814 7862 1866 7883
rect 1879 7862 1931 7883
rect 1944 7862 1996 7883
rect 2009 7883 2012 7914
rect 2012 7883 2046 7914
rect 2046 7883 2061 7914
rect 2009 7862 2061 7883
rect 2074 7883 2085 7914
rect 2085 7883 2119 7914
rect 2119 7883 2126 7914
rect 2074 7862 2126 7883
rect 2139 7883 2158 7914
rect 2158 7883 2191 7914
rect 2204 7883 2231 7914
rect 2231 7883 2256 7914
rect 2269 7883 2304 7914
rect 2304 7883 2321 7914
rect 2334 7883 2338 7914
rect 2338 7883 2377 7914
rect 2377 7883 2386 7914
rect 2399 7883 2411 7914
rect 2411 7883 2450 7914
rect 2450 7883 2451 7914
rect 2464 7883 2484 7914
rect 2484 7883 2516 7914
rect 2529 7883 2557 7914
rect 2557 7883 2581 7914
rect 2139 7862 2191 7883
rect 2204 7862 2256 7883
rect 2269 7862 2321 7883
rect 2334 7862 2386 7883
rect 2399 7862 2451 7883
rect 2464 7862 2516 7883
rect 2529 7862 2581 7883
rect 2594 7883 2596 7914
rect 2596 7883 2630 7914
rect 2630 7883 2646 7914
rect 2594 7862 2646 7883
rect 2659 7883 2669 7914
rect 2669 7883 2703 7914
rect 2703 7883 2711 7914
rect 2659 7862 2711 7883
rect 2724 7883 2742 7914
rect 2742 7883 2776 7914
rect 2724 7862 2776 7883
rect 2789 7883 2815 7914
rect 2815 7883 2841 7914
rect 2854 7883 2888 7914
rect 2888 7883 2906 7914
rect 2919 7883 2922 7914
rect 2922 7883 2961 7914
rect 2961 7883 2971 7914
rect 2984 7883 2995 7914
rect 2995 7883 3034 7914
rect 3034 7883 3036 7914
rect 3049 7883 3068 7914
rect 3068 7883 3101 7914
rect 3114 7883 3141 7914
rect 3141 7883 3166 7914
rect 2789 7862 2841 7883
rect 2854 7862 2906 7883
rect 2919 7862 2971 7883
rect 2984 7862 3036 7883
rect 3049 7862 3101 7883
rect 3114 7862 3166 7883
rect 3179 7883 3180 7914
rect 3180 7883 3214 7914
rect 3214 7883 3231 7914
rect 3179 7862 3231 7883
rect 3244 7883 3253 7914
rect 3253 7883 3287 7914
rect 3287 7883 3296 7914
rect 3244 7862 3296 7883
rect 3309 7883 3326 7914
rect 3326 7883 3360 7914
rect 3360 7883 3361 7914
rect 3309 7862 3361 7883
rect 3374 7883 3399 7914
rect 3399 7883 3426 7914
rect 3439 7883 3472 7914
rect 3472 7883 3491 7914
rect 3504 7883 3506 7914
rect 3506 7883 3545 7914
rect 3545 7883 3556 7914
rect 3569 7883 3579 7914
rect 3579 7883 3618 7914
rect 3618 7883 3621 7914
rect 3374 7862 3426 7883
rect 3439 7862 3491 7883
rect 3504 7862 3556 7883
rect 3569 7862 3621 7883
rect 631 7845 683 7850
rect 631 7798 683 7845
rect 631 7734 683 7786
rect 749 7773 801 7796
rect 814 7773 866 7796
rect 879 7773 931 7796
rect 944 7773 996 7796
rect 1009 7773 1061 7796
rect 1073 7773 1125 7796
rect 1137 7773 1189 7796
rect 749 7744 801 7773
rect 814 7744 843 7773
rect 843 7744 866 7773
rect 879 7744 916 7773
rect 916 7744 931 7773
rect 944 7744 950 7773
rect 950 7744 989 7773
rect 989 7744 996 7773
rect 1009 7744 1023 7773
rect 1023 7744 1061 7773
rect 1073 7744 1096 7773
rect 1096 7744 1125 7773
rect 1137 7744 1169 7773
rect 1169 7744 1189 7773
rect 1201 7773 1253 7796
rect 1201 7744 1208 7773
rect 1208 7744 1242 7773
rect 1242 7744 1253 7773
rect 1265 7773 1317 7796
rect 1265 7744 1281 7773
rect 1281 7744 1315 7773
rect 1315 7744 1317 7773
rect 1329 7773 1381 7796
rect 1393 7773 1445 7796
rect 1457 7773 1509 7796
rect 1521 7773 1573 7796
rect 1585 7773 1637 7796
rect 1649 7773 1701 7796
rect 1329 7744 1354 7773
rect 1354 7744 1381 7773
rect 1393 7744 1427 7773
rect 1427 7744 1445 7773
rect 1457 7744 1461 7773
rect 1461 7744 1500 7773
rect 1500 7744 1509 7773
rect 1521 7744 1534 7773
rect 1534 7744 1573 7773
rect 1585 7744 1607 7773
rect 1607 7744 1637 7773
rect 1649 7744 1680 7773
rect 1680 7744 1701 7773
rect 1713 7773 1765 7796
rect 1713 7744 1719 7773
rect 1719 7744 1753 7773
rect 1753 7744 1765 7773
rect 1777 7773 1829 7796
rect 1777 7744 1792 7773
rect 1792 7744 1826 7773
rect 1826 7744 1829 7773
rect 1841 7773 1893 7796
rect 1905 7773 1957 7796
rect 1969 7773 2021 7796
rect 2033 7773 2085 7796
rect 2097 7773 2149 7796
rect 2161 7773 2213 7796
rect 1841 7744 1865 7773
rect 1865 7744 1893 7773
rect 1905 7744 1938 7773
rect 1938 7744 1957 7773
rect 1969 7744 1972 7773
rect 1972 7744 2011 7773
rect 2011 7744 2021 7773
rect 2033 7744 2045 7773
rect 2045 7744 2084 7773
rect 2084 7744 2085 7773
rect 2097 7744 2118 7773
rect 2118 7744 2149 7773
rect 2161 7744 2191 7773
rect 2191 7744 2213 7773
rect 2225 7773 2277 7796
rect 2225 7744 2230 7773
rect 2230 7744 2264 7773
rect 2264 7744 2277 7773
rect 2289 7773 2341 7796
rect 2289 7744 2303 7773
rect 2303 7744 2337 7773
rect 2337 7744 2341 7773
rect 2353 7773 2405 7796
rect 2417 7773 2469 7796
rect 2481 7773 2533 7796
rect 2545 7773 2597 7796
rect 2609 7773 2661 7796
rect 2673 7773 2725 7796
rect 2353 7744 2376 7773
rect 2376 7744 2405 7773
rect 2417 7744 2449 7773
rect 2449 7744 2469 7773
rect 2481 7744 2483 7773
rect 2483 7744 2522 7773
rect 2522 7744 2533 7773
rect 2545 7744 2556 7773
rect 2556 7744 2595 7773
rect 2595 7744 2597 7773
rect 2609 7744 2629 7773
rect 2629 7744 2661 7773
rect 2673 7744 2702 7773
rect 2702 7744 2725 7773
rect 2737 7773 2789 7796
rect 2737 7744 2741 7773
rect 2741 7744 2775 7773
rect 2775 7744 2789 7773
rect 2801 7773 2853 7796
rect 2801 7744 2814 7773
rect 2814 7744 2848 7773
rect 2848 7744 2853 7773
rect 2865 7773 2917 7796
rect 2929 7773 2981 7796
rect 2993 7773 3045 7796
rect 3057 7773 3109 7796
rect 3121 7773 3173 7796
rect 3185 7773 3237 7796
rect 2865 7744 2887 7773
rect 2887 7744 2917 7773
rect 2929 7744 2960 7773
rect 2960 7744 2981 7773
rect 2993 7744 2994 7773
rect 2994 7744 3033 7773
rect 3033 7744 3045 7773
rect 3057 7744 3067 7773
rect 3067 7744 3106 7773
rect 3106 7744 3109 7773
rect 3121 7744 3140 7773
rect 3140 7744 3173 7773
rect 3185 7744 3213 7773
rect 3213 7744 3237 7773
rect 3249 7773 3301 7796
rect 3249 7744 3252 7773
rect 3252 7744 3286 7773
rect 3286 7744 3301 7773
rect 3313 7773 3365 7796
rect 3313 7744 3325 7773
rect 3325 7744 3359 7773
rect 3359 7744 3365 7773
rect 3377 7773 3429 7796
rect 3441 7773 3493 7796
rect 3505 7773 3557 7796
rect 3569 7773 3621 7796
rect 3377 7744 3398 7773
rect 3398 7744 3429 7773
rect 3441 7744 3471 7773
rect 3471 7744 3493 7773
rect 3505 7744 3544 7773
rect 3544 7744 3557 7773
rect 3569 7744 3578 7773
rect 3578 7744 3617 7773
rect 3617 7744 3621 7773
rect 631 7670 683 7722
rect 749 7680 801 7732
rect 631 7606 683 7658
rect 749 7616 801 7668
rect 631 7542 683 7594
rect 749 7552 801 7604
rect 631 7478 683 7530
rect 749 7488 801 7540
rect 631 7414 683 7466
rect 749 7424 801 7476
rect 631 7350 683 7402
rect 749 7360 801 7412
rect 631 7286 683 7338
rect 749 7296 801 7348
rect 631 7222 683 7274
rect 749 7231 801 7283
rect 631 7158 683 7210
rect 749 7166 801 7218
rect 631 7094 683 7146
rect 749 7101 801 7153
rect 631 7030 683 7082
rect 749 7036 801 7088
rect 631 6966 683 7018
rect 749 6971 801 7023
rect 631 6902 683 6954
rect 749 6906 801 6958
rect 631 6838 683 6890
rect 749 6841 801 6893
rect 631 6774 683 6826
rect 749 6776 801 6828
rect 631 6710 683 6762
rect 749 6711 801 6763
rect 631 6646 683 6698
rect 749 6646 801 6698
rect 631 6582 683 6634
rect 749 6581 801 6633
rect 631 6518 683 6570
rect 749 6516 801 6568
rect 631 6454 683 6506
rect 749 6451 801 6503
rect 631 6390 683 6442
rect 749 6386 801 6438
rect 631 6326 683 6378
rect 749 6321 801 6373
rect 631 6262 683 6314
rect 749 6256 801 6308
rect 631 6198 683 6250
rect 749 6191 801 6243
rect 631 6134 683 6186
rect 749 6126 801 6178
rect 631 6070 683 6122
rect 749 6083 801 6113
rect 749 6061 801 6083
rect 631 6011 683 6058
rect 749 6044 801 6048
rect 631 6006 683 6011
rect 749 6010 770 6044
rect 770 6010 801 6044
rect 749 5996 801 6010
rect 631 5972 683 5994
rect 631 5942 660 5972
rect 660 5942 683 5972
rect 749 5971 801 5983
rect 749 5937 770 5971
rect 770 5937 801 5971
rect 749 5931 801 5937
rect 631 5899 683 5929
rect 631 5877 660 5899
rect 660 5877 683 5899
rect 749 5898 801 5918
rect 749 5866 770 5898
rect 770 5866 801 5898
rect 631 5826 683 5864
rect 631 5812 660 5826
rect 660 5812 683 5826
rect 631 5792 660 5799
rect 660 5792 683 5799
rect 749 5825 801 5853
rect 8895 7428 8947 7434
rect 8895 7394 8899 7428
rect 8899 7394 8933 7428
rect 8933 7394 8947 7428
rect 8895 7382 8947 7394
rect 8959 7428 9011 7434
rect 8959 7394 8971 7428
rect 8971 7394 9005 7428
rect 9005 7394 9011 7428
rect 8959 7382 9011 7394
rect 3446 7243 3498 7295
rect 3511 7243 3563 7295
rect 3576 7243 3628 7295
rect 3641 7243 3693 7295
rect 3706 7264 3719 7295
rect 3719 7264 3753 7295
rect 3753 7264 3758 7295
rect 3706 7243 3758 7264
rect 3771 7243 3823 7295
rect 3836 7243 3888 7295
rect 3901 7243 3953 7295
rect 3966 7243 4018 7295
rect 4031 7264 4065 7295
rect 4065 7264 4083 7295
rect 4031 7243 4083 7264
rect 4096 7243 4148 7295
rect 4161 7243 4213 7295
rect 4226 7243 4278 7295
rect 4291 7243 4343 7295
rect 4356 7264 4377 7295
rect 4377 7264 4408 7295
rect 4356 7243 4408 7264
rect 4421 7243 4473 7295
rect 4486 7243 4538 7295
rect 4551 7243 4603 7295
rect 4616 7264 4655 7295
rect 4655 7264 4668 7295
rect 4681 7264 4689 7295
rect 4689 7264 4733 7295
rect 4616 7243 4668 7264
rect 4681 7243 4733 7264
rect 4746 7243 4798 7295
rect 4811 7243 4863 7295
rect 4876 7243 4928 7295
rect 4941 7264 4967 7295
rect 4967 7264 4993 7295
rect 4941 7243 4993 7264
rect 5006 7243 5058 7295
rect 5071 7243 5123 7295
rect 5136 7243 5188 7295
rect 5201 7243 5253 7295
rect 5266 7264 5279 7295
rect 5279 7264 5313 7295
rect 5313 7264 5318 7295
rect 5266 7243 5318 7264
rect 5331 7243 5383 7295
rect 5396 7243 5448 7295
rect 5461 7243 5513 7295
rect 5526 7243 5578 7295
rect 5591 7264 5625 7295
rect 5625 7264 5903 7295
rect 5903 7264 5937 7295
rect 5937 7264 6215 7295
rect 6215 7264 6249 7295
rect 6249 7264 6527 7295
rect 6527 7264 6561 7295
rect 6561 7264 6839 7295
rect 6839 7264 6873 7295
rect 6873 7264 7151 7295
rect 7151 7264 7185 7295
rect 7185 7264 7463 7295
rect 7463 7264 7497 7295
rect 7497 7264 7775 7295
rect 7775 7264 7809 7295
rect 7809 7264 8087 7295
rect 8087 7264 8121 7295
rect 8121 7264 8399 7295
rect 8399 7264 8433 7295
rect 8433 7264 8711 7295
rect 8711 7264 8745 7295
rect 8745 7264 9023 7295
rect 9023 7264 9057 7295
rect 9057 7264 9099 7295
rect 3446 7179 3498 7231
rect 3511 7179 3563 7231
rect 3576 7179 3628 7231
rect 3641 7179 3693 7231
rect 3706 7224 3758 7231
rect 3706 7190 3719 7224
rect 3719 7190 3753 7224
rect 3753 7190 3758 7224
rect 3706 7179 3758 7190
rect 3771 7179 3823 7231
rect 3836 7179 3888 7231
rect 3901 7179 3953 7231
rect 3966 7179 4018 7231
rect 4031 7224 4083 7231
rect 4031 7190 4065 7224
rect 4065 7190 4083 7224
rect 4031 7179 4083 7190
rect 4096 7179 4148 7231
rect 4161 7179 4213 7231
rect 4226 7179 4278 7231
rect 4291 7179 4343 7231
rect 4356 7224 4408 7231
rect 4356 7190 4377 7224
rect 4377 7190 4408 7224
rect 4356 7179 4408 7190
rect 4421 7179 4473 7231
rect 4486 7179 4538 7231
rect 4551 7179 4603 7231
rect 4616 7224 4668 7231
rect 4681 7224 4733 7231
rect 4616 7190 4655 7224
rect 4655 7190 4668 7224
rect 4681 7190 4689 7224
rect 4689 7190 4733 7224
rect 4616 7179 4668 7190
rect 4681 7179 4733 7190
rect 4746 7179 4798 7231
rect 4811 7179 4863 7231
rect 4876 7179 4928 7231
rect 4941 7224 4993 7231
rect 4941 7190 4967 7224
rect 4967 7190 4993 7224
rect 4941 7179 4993 7190
rect 5006 7179 5058 7231
rect 5071 7179 5123 7231
rect 5136 7179 5188 7231
rect 5201 7179 5253 7231
rect 5266 7224 5318 7231
rect 5266 7190 5279 7224
rect 5279 7190 5313 7224
rect 5313 7190 5318 7224
rect 5266 7179 5318 7190
rect 5331 7179 5383 7231
rect 5396 7179 5448 7231
rect 5461 7179 5513 7231
rect 5526 7179 5578 7231
rect 5591 7224 9099 7264
rect 5591 7190 5625 7224
rect 5625 7190 5903 7224
rect 5903 7190 5937 7224
rect 5937 7190 6215 7224
rect 6215 7190 6249 7224
rect 6249 7190 6527 7224
rect 6527 7190 6561 7224
rect 6561 7190 6839 7224
rect 6839 7190 6873 7224
rect 6873 7190 7151 7224
rect 7151 7190 7185 7224
rect 7185 7190 7463 7224
rect 7463 7190 7497 7224
rect 7497 7190 7775 7224
rect 7775 7190 7809 7224
rect 7809 7190 8087 7224
rect 8087 7190 8121 7224
rect 8121 7190 8399 7224
rect 8399 7190 8433 7224
rect 8433 7190 8711 7224
rect 8711 7190 8745 7224
rect 8745 7190 9023 7224
rect 9023 7190 9057 7224
rect 9057 7190 9099 7224
rect 3446 7115 3498 7167
rect 3511 7115 3563 7167
rect 3576 7115 3628 7167
rect 3641 7115 3693 7167
rect 3706 7150 3758 7167
rect 3706 7116 3719 7150
rect 3719 7116 3753 7150
rect 3753 7116 3758 7150
rect 3706 7115 3758 7116
rect 3771 7115 3823 7167
rect 3836 7115 3888 7167
rect 3901 7115 3953 7167
rect 3966 7115 4018 7167
rect 4031 7150 4083 7167
rect 4031 7116 4065 7150
rect 4065 7116 4083 7150
rect 4031 7115 4083 7116
rect 4096 7115 4148 7167
rect 4161 7115 4213 7167
rect 4226 7115 4278 7167
rect 4291 7115 4343 7167
rect 4356 7150 4408 7167
rect 4356 7116 4377 7150
rect 4377 7116 4408 7150
rect 4356 7115 4408 7116
rect 4421 7115 4473 7167
rect 4486 7115 4538 7167
rect 4551 7115 4603 7167
rect 4616 7150 4668 7167
rect 4681 7150 4733 7167
rect 4616 7116 4655 7150
rect 4655 7116 4668 7150
rect 4681 7116 4689 7150
rect 4689 7116 4733 7150
rect 4616 7115 4668 7116
rect 4681 7115 4733 7116
rect 4746 7115 4798 7167
rect 4811 7115 4863 7167
rect 4876 7115 4928 7167
rect 4941 7150 4993 7167
rect 4941 7116 4967 7150
rect 4967 7116 4993 7150
rect 4941 7115 4993 7116
rect 5006 7115 5058 7167
rect 5071 7115 5123 7167
rect 5136 7115 5188 7167
rect 5201 7115 5253 7167
rect 5266 7150 5318 7167
rect 5266 7116 5279 7150
rect 5279 7116 5313 7150
rect 5313 7116 5318 7150
rect 5266 7115 5318 7116
rect 5331 7115 5383 7167
rect 5396 7115 5448 7167
rect 5461 7115 5513 7167
rect 5526 7115 5578 7167
rect 5591 7150 9099 7190
rect 5591 7116 5625 7150
rect 5625 7116 5903 7150
rect 5903 7116 5937 7150
rect 5937 7116 6215 7150
rect 6215 7116 6249 7150
rect 6249 7116 6527 7150
rect 6527 7116 6561 7150
rect 6561 7116 6839 7150
rect 6839 7116 6873 7150
rect 6873 7116 7151 7150
rect 7151 7116 7185 7150
rect 7185 7116 7463 7150
rect 7463 7116 7497 7150
rect 7497 7116 7775 7150
rect 7775 7116 7809 7150
rect 7809 7116 8087 7150
rect 8087 7116 8121 7150
rect 8121 7116 8399 7150
rect 8399 7116 8433 7150
rect 8433 7116 8711 7150
rect 8711 7116 8745 7150
rect 8745 7116 9023 7150
rect 9023 7116 9057 7150
rect 9057 7116 9099 7150
rect 3446 7051 3498 7103
rect 3511 7051 3563 7103
rect 3576 7051 3628 7103
rect 3641 7051 3693 7103
rect 3706 7076 3758 7103
rect 3706 7051 3719 7076
rect 3719 7051 3753 7076
rect 3753 7051 3758 7076
rect 3771 7051 3823 7103
rect 3836 7051 3888 7103
rect 3901 7051 3953 7103
rect 3966 7051 4018 7103
rect 4031 7076 4083 7103
rect 4031 7051 4065 7076
rect 4065 7051 4083 7076
rect 4096 7051 4148 7103
rect 4161 7051 4213 7103
rect 4226 7051 4278 7103
rect 4291 7051 4343 7103
rect 4356 7076 4408 7103
rect 4356 7051 4377 7076
rect 4377 7051 4408 7076
rect 4421 7051 4473 7103
rect 4486 7051 4538 7103
rect 4551 7051 4603 7103
rect 4616 7076 4668 7103
rect 4681 7076 4733 7103
rect 4616 7051 4655 7076
rect 4655 7051 4668 7076
rect 4681 7051 4689 7076
rect 4689 7051 4733 7076
rect 4746 7051 4798 7103
rect 4811 7051 4863 7103
rect 4876 7051 4928 7103
rect 4941 7076 4993 7103
rect 4941 7051 4967 7076
rect 4967 7051 4993 7076
rect 5006 7051 5058 7103
rect 5071 7051 5123 7103
rect 5136 7051 5188 7103
rect 5201 7051 5253 7103
rect 5266 7076 5318 7103
rect 5266 7051 5279 7076
rect 5279 7051 5313 7076
rect 5313 7051 5318 7076
rect 5331 7051 5383 7103
rect 5396 7051 5448 7103
rect 5461 7051 5513 7103
rect 5526 7051 5578 7103
rect 5591 7076 9099 7116
rect 5591 7042 5625 7076
rect 5625 7042 5903 7076
rect 5903 7042 5937 7076
rect 5937 7042 6215 7076
rect 6215 7042 6249 7076
rect 6249 7042 6527 7076
rect 6527 7042 6561 7076
rect 6561 7042 6839 7076
rect 6839 7042 6873 7076
rect 6873 7042 7151 7076
rect 7151 7042 7185 7076
rect 7185 7042 7463 7076
rect 7463 7042 7497 7076
rect 7497 7042 7775 7076
rect 7775 7042 7809 7076
rect 7809 7042 8087 7076
rect 8087 7042 8121 7076
rect 8121 7042 8399 7076
rect 8399 7042 8433 7076
rect 8433 7042 8711 7076
rect 8711 7042 8745 7076
rect 8745 7042 9023 7076
rect 9023 7042 9057 7076
rect 9057 7042 9099 7076
rect 3446 6987 3498 7039
rect 3511 6987 3563 7039
rect 3576 6987 3628 7039
rect 3641 6987 3693 7039
rect 3706 7002 3758 7039
rect 3706 6987 3719 7002
rect 3719 6987 3753 7002
rect 3753 6987 3758 7002
rect 3771 6987 3823 7039
rect 3836 6987 3888 7039
rect 3901 6987 3953 7039
rect 3966 6987 4018 7039
rect 4031 7001 4083 7039
rect 4031 6987 4065 7001
rect 4065 6987 4083 7001
rect 4096 6987 4148 7039
rect 4161 6987 4213 7039
rect 4226 6987 4278 7039
rect 4291 6987 4343 7039
rect 4356 7002 4408 7039
rect 4356 6987 4377 7002
rect 4377 6987 4408 7002
rect 4421 6987 4473 7039
rect 4486 6987 4538 7039
rect 4551 6987 4603 7039
rect 4616 7001 4668 7039
rect 4681 7001 4733 7039
rect 4616 6987 4655 7001
rect 4655 6987 4668 7001
rect 4681 6987 4689 7001
rect 4689 6987 4733 7001
rect 4746 6987 4798 7039
rect 4811 6987 4863 7039
rect 4876 6987 4928 7039
rect 4941 7002 4993 7039
rect 4941 6987 4967 7002
rect 4967 6987 4993 7002
rect 5006 6987 5058 7039
rect 5071 6987 5123 7039
rect 5136 6987 5188 7039
rect 5201 6987 5253 7039
rect 5266 7001 5318 7039
rect 5266 6987 5279 7001
rect 5279 6987 5313 7001
rect 5313 6987 5318 7001
rect 5331 6987 5383 7039
rect 5396 6987 5448 7039
rect 5461 6987 5513 7039
rect 5526 6987 5578 7039
rect 5591 7002 9099 7042
rect 3446 6923 3498 6975
rect 3511 6923 3563 6975
rect 3576 6923 3628 6975
rect 3641 6923 3693 6975
rect 3706 6968 3719 6975
rect 3719 6968 3753 6975
rect 3753 6968 3758 6975
rect 3706 6927 3758 6968
rect 3706 6923 3719 6927
rect 3719 6923 3753 6927
rect 3753 6923 3758 6927
rect 3771 6923 3823 6975
rect 3836 6923 3888 6975
rect 3901 6923 3953 6975
rect 3966 6923 4018 6975
rect 4031 6967 4065 6975
rect 4065 6967 4083 6975
rect 4031 6926 4083 6967
rect 4031 6923 4065 6926
rect 4065 6923 4083 6926
rect 4096 6923 4148 6975
rect 4161 6923 4213 6975
rect 4226 6923 4278 6975
rect 4291 6923 4343 6975
rect 4356 6968 4377 6975
rect 4377 6968 4408 6975
rect 4356 6927 4408 6968
rect 4356 6923 4377 6927
rect 4377 6923 4408 6927
rect 4421 6923 4473 6975
rect 4486 6923 4538 6975
rect 4551 6923 4603 6975
rect 4616 6967 4655 6975
rect 4655 6967 4668 6975
rect 4681 6967 4689 6975
rect 4689 6967 4733 6975
rect 4616 6926 4668 6967
rect 4681 6926 4733 6967
rect 4616 6923 4655 6926
rect 4655 6923 4668 6926
rect 4681 6923 4689 6926
rect 4689 6923 4733 6926
rect 4746 6923 4798 6975
rect 4811 6923 4863 6975
rect 4876 6923 4928 6975
rect 4941 6968 4967 6975
rect 4967 6968 4993 6975
rect 4941 6927 4993 6968
rect 4941 6923 4967 6927
rect 4967 6923 4993 6927
rect 5006 6923 5058 6975
rect 5071 6923 5123 6975
rect 5136 6923 5188 6975
rect 5201 6923 5253 6975
rect 5266 6967 5279 6975
rect 5279 6967 5313 6975
rect 5313 6967 5318 6975
rect 5266 6926 5318 6967
rect 5266 6923 5279 6926
rect 5279 6923 5313 6926
rect 5313 6923 5318 6926
rect 5331 6923 5383 6975
rect 5396 6923 5448 6975
rect 5461 6923 5513 6975
rect 5526 6923 5578 6975
rect 5591 6968 5625 7002
rect 5625 7001 6215 7002
rect 5625 6968 5903 7001
rect 5591 6967 5903 6968
rect 5903 6967 5937 7001
rect 5937 6968 6215 7001
rect 6215 6968 6249 7002
rect 6249 7001 6839 7002
rect 6249 6968 6527 7001
rect 5937 6967 6527 6968
rect 6527 6967 6561 7001
rect 6561 6968 6839 7001
rect 6839 6968 6873 7002
rect 6873 7001 7463 7002
rect 6873 6968 7151 7001
rect 6561 6967 7151 6968
rect 7151 6967 7185 7001
rect 7185 6968 7463 7001
rect 7463 6968 7497 7002
rect 7497 7001 8399 7002
rect 7497 6968 7775 7001
rect 7185 6967 7775 6968
rect 7775 6967 7809 7001
rect 7809 6967 8087 7001
rect 8087 6967 8121 7001
rect 8121 6968 8399 7001
rect 8399 6968 8433 7002
rect 8433 7001 9023 7002
rect 8433 6968 8711 7001
rect 8121 6967 8711 6968
rect 8711 6967 8745 7001
rect 8745 6968 9023 7001
rect 9023 6968 9057 7002
rect 9057 6968 9099 7002
rect 8745 6967 9099 6968
rect 5591 6927 9099 6967
rect 3446 6859 3498 6911
rect 3511 6859 3563 6911
rect 3576 6859 3628 6911
rect 3641 6859 3693 6911
rect 3706 6893 3719 6911
rect 3719 6893 3753 6911
rect 3753 6893 3758 6911
rect 3706 6859 3758 6893
rect 3771 6859 3823 6911
rect 3836 6859 3888 6911
rect 3901 6859 3953 6911
rect 3966 6859 4018 6911
rect 4031 6892 4065 6911
rect 4065 6892 4083 6911
rect 4031 6859 4083 6892
rect 4096 6859 4148 6911
rect 4161 6859 4213 6911
rect 4226 6859 4278 6911
rect 4291 6859 4343 6911
rect 4356 6893 4377 6911
rect 4377 6893 4408 6911
rect 4356 6859 4408 6893
rect 4421 6859 4473 6911
rect 4486 6859 4538 6911
rect 4551 6859 4603 6911
rect 4616 6892 4655 6911
rect 4655 6892 4668 6911
rect 4681 6892 4689 6911
rect 4689 6892 4733 6911
rect 4616 6859 4668 6892
rect 4681 6859 4733 6892
rect 4746 6859 4798 6911
rect 4811 6859 4863 6911
rect 4876 6859 4928 6911
rect 4941 6893 4967 6911
rect 4967 6893 4993 6911
rect 4941 6859 4993 6893
rect 5006 6859 5058 6911
rect 5071 6859 5123 6911
rect 5136 6859 5188 6911
rect 5201 6859 5253 6911
rect 5266 6892 5279 6911
rect 5279 6892 5313 6911
rect 5313 6892 5318 6911
rect 5266 6859 5318 6892
rect 5331 6859 5383 6911
rect 5396 6859 5448 6911
rect 5461 6859 5513 6911
rect 5526 6859 5578 6911
rect 5591 6893 5625 6927
rect 5625 6926 6215 6927
rect 5625 6893 5903 6926
rect 5591 6892 5903 6893
rect 5903 6892 5937 6926
rect 5937 6893 6215 6926
rect 6215 6893 6249 6927
rect 6249 6926 6839 6927
rect 6249 6893 6527 6926
rect 5937 6892 6527 6893
rect 6527 6892 6561 6926
rect 6561 6893 6839 6926
rect 6839 6893 6873 6927
rect 6873 6926 7463 6927
rect 6873 6893 7151 6926
rect 6561 6892 7151 6893
rect 7151 6892 7185 6926
rect 7185 6893 7463 6926
rect 7463 6893 7497 6927
rect 7497 6926 8399 6927
rect 7497 6893 7775 6926
rect 7185 6892 7775 6893
rect 7775 6892 7809 6926
rect 7809 6892 8087 6926
rect 8087 6892 8121 6926
rect 8121 6893 8399 6926
rect 8399 6893 8433 6927
rect 8433 6926 9023 6927
rect 8433 6893 8711 6926
rect 8121 6892 8711 6893
rect 8711 6892 8745 6926
rect 8745 6893 9023 6926
rect 9023 6893 9057 6927
rect 9057 6893 9099 6927
rect 8745 6892 9099 6893
rect 5591 6852 9099 6892
rect 3446 6795 3498 6847
rect 3511 6795 3563 6847
rect 3576 6795 3628 6847
rect 3641 6795 3693 6847
rect 3706 6818 3719 6847
rect 3719 6818 3753 6847
rect 3753 6818 3758 6847
rect 3706 6795 3758 6818
rect 3771 6795 3823 6847
rect 3836 6795 3888 6847
rect 3901 6795 3953 6847
rect 3966 6795 4018 6847
rect 4031 6817 4065 6847
rect 4065 6817 4083 6847
rect 4031 6795 4083 6817
rect 4096 6795 4148 6847
rect 4161 6795 4213 6847
rect 4226 6795 4278 6847
rect 4291 6795 4343 6847
rect 4356 6818 4377 6847
rect 4377 6818 4408 6847
rect 4356 6795 4408 6818
rect 4421 6795 4473 6847
rect 4486 6795 4538 6847
rect 4551 6795 4603 6847
rect 4616 6817 4655 6847
rect 4655 6817 4668 6847
rect 4681 6817 4689 6847
rect 4689 6817 4733 6847
rect 4616 6795 4668 6817
rect 4681 6795 4733 6817
rect 4746 6795 4798 6847
rect 4811 6795 4863 6847
rect 4876 6795 4928 6847
rect 4941 6818 4967 6847
rect 4967 6818 4993 6847
rect 4941 6795 4993 6818
rect 5006 6795 5058 6847
rect 5071 6795 5123 6847
rect 5136 6795 5188 6847
rect 5201 6795 5253 6847
rect 5266 6817 5279 6847
rect 5279 6817 5313 6847
rect 5313 6817 5318 6847
rect 5266 6795 5318 6817
rect 5331 6795 5383 6847
rect 5396 6795 5448 6847
rect 5461 6795 5513 6847
rect 5526 6795 5578 6847
rect 5591 6818 5625 6852
rect 5625 6851 6215 6852
rect 5625 6818 5903 6851
rect 5591 6817 5903 6818
rect 5903 6817 5937 6851
rect 5937 6818 6215 6851
rect 6215 6818 6249 6852
rect 6249 6851 6839 6852
rect 6249 6818 6527 6851
rect 5937 6817 6527 6818
rect 6527 6817 6561 6851
rect 6561 6818 6839 6851
rect 6839 6818 6873 6852
rect 6873 6851 7463 6852
rect 6873 6818 7151 6851
rect 6561 6817 7151 6818
rect 7151 6817 7185 6851
rect 7185 6818 7463 6851
rect 7463 6818 7497 6852
rect 7497 6851 8399 6852
rect 7497 6818 7775 6851
rect 7185 6817 7775 6818
rect 7775 6817 7809 6851
rect 7809 6817 8087 6851
rect 8087 6817 8121 6851
rect 8121 6818 8399 6851
rect 8399 6818 8433 6852
rect 8433 6851 9023 6852
rect 8433 6818 8711 6851
rect 8121 6817 8711 6818
rect 8711 6817 8745 6851
rect 8745 6818 9023 6851
rect 9023 6818 9057 6852
rect 9057 6818 9099 6852
rect 8745 6817 9099 6818
rect 3446 6731 3498 6783
rect 3511 6731 3563 6783
rect 3576 6731 3628 6783
rect 3641 6731 3693 6783
rect 3706 6777 3758 6783
rect 3706 6743 3719 6777
rect 3719 6743 3753 6777
rect 3753 6743 3758 6777
rect 3706 6731 3758 6743
rect 3771 6731 3823 6783
rect 3836 6731 3888 6783
rect 3901 6731 3953 6783
rect 3966 6731 4018 6783
rect 4031 6776 4083 6783
rect 4031 6742 4065 6776
rect 4065 6742 4083 6776
rect 4031 6731 4083 6742
rect 4096 6731 4148 6783
rect 4161 6731 4213 6783
rect 4226 6731 4278 6783
rect 4291 6731 4343 6783
rect 4356 6777 4408 6783
rect 4356 6743 4377 6777
rect 4377 6743 4408 6777
rect 4356 6731 4408 6743
rect 4421 6731 4473 6783
rect 4486 6731 4538 6783
rect 4551 6731 4603 6783
rect 4616 6776 4668 6783
rect 4681 6776 4733 6783
rect 4616 6742 4655 6776
rect 4655 6742 4668 6776
rect 4681 6742 4689 6776
rect 4689 6742 4733 6776
rect 4616 6731 4668 6742
rect 4681 6731 4733 6742
rect 4746 6731 4798 6783
rect 4811 6731 4863 6783
rect 4876 6731 4928 6783
rect 4941 6777 4993 6783
rect 4941 6743 4967 6777
rect 4967 6743 4993 6777
rect 4941 6731 4993 6743
rect 5006 6731 5058 6783
rect 5071 6731 5123 6783
rect 5136 6731 5188 6783
rect 5201 6731 5253 6783
rect 5266 6776 5318 6783
rect 5266 6742 5279 6776
rect 5279 6742 5313 6776
rect 5313 6742 5318 6776
rect 5266 6731 5318 6742
rect 5331 6731 5383 6783
rect 5396 6731 5448 6783
rect 5461 6731 5513 6783
rect 5526 6731 5578 6783
rect 5591 6777 9099 6817
rect 5591 6743 5625 6777
rect 5625 6776 6215 6777
rect 5625 6743 5903 6776
rect 5591 6742 5903 6743
rect 5903 6742 5937 6776
rect 5937 6743 6215 6776
rect 6215 6743 6249 6777
rect 6249 6776 6839 6777
rect 6249 6743 6527 6776
rect 5937 6742 6527 6743
rect 6527 6742 6561 6776
rect 6561 6743 6839 6776
rect 6839 6743 6873 6777
rect 6873 6776 7463 6777
rect 6873 6743 7151 6776
rect 6561 6742 7151 6743
rect 7151 6742 7185 6776
rect 7185 6743 7463 6776
rect 7463 6743 7497 6777
rect 7497 6776 8399 6777
rect 7497 6743 7775 6776
rect 7185 6742 7775 6743
rect 7775 6742 7809 6776
rect 7809 6742 8087 6776
rect 8087 6742 8121 6776
rect 8121 6743 8399 6776
rect 8399 6743 8433 6777
rect 8433 6776 9023 6777
rect 8433 6743 8711 6776
rect 8121 6742 8711 6743
rect 8711 6742 8745 6776
rect 8745 6743 9023 6776
rect 9023 6743 9057 6777
rect 9057 6743 9099 6777
rect 8745 6742 9099 6743
rect 3446 6667 3498 6719
rect 3511 6667 3563 6719
rect 3576 6667 3628 6719
rect 3641 6667 3693 6719
rect 3706 6702 3758 6719
rect 3706 6668 3719 6702
rect 3719 6668 3753 6702
rect 3753 6668 3758 6702
rect 3706 6667 3758 6668
rect 3771 6667 3823 6719
rect 3836 6667 3888 6719
rect 3901 6667 3953 6719
rect 3966 6667 4018 6719
rect 4031 6701 4083 6719
rect 4031 6667 4065 6701
rect 4065 6667 4083 6701
rect 4096 6667 4148 6719
rect 4161 6667 4213 6719
rect 4226 6667 4278 6719
rect 4291 6667 4343 6719
rect 4356 6702 4408 6719
rect 4356 6668 4377 6702
rect 4377 6668 4408 6702
rect 4356 6667 4408 6668
rect 4421 6667 4473 6719
rect 4486 6667 4538 6719
rect 4551 6667 4603 6719
rect 4616 6701 4668 6719
rect 4681 6701 4733 6719
rect 4616 6667 4655 6701
rect 4655 6667 4668 6701
rect 4681 6667 4689 6701
rect 4689 6667 4733 6701
rect 4746 6667 4798 6719
rect 4811 6667 4863 6719
rect 4876 6667 4928 6719
rect 4941 6702 4993 6719
rect 4941 6668 4967 6702
rect 4967 6668 4993 6702
rect 4941 6667 4993 6668
rect 5006 6667 5058 6719
rect 5071 6667 5123 6719
rect 5136 6667 5188 6719
rect 5201 6667 5253 6719
rect 5266 6701 5318 6719
rect 5266 6667 5279 6701
rect 5279 6667 5313 6701
rect 5313 6667 5318 6701
rect 5331 6667 5383 6719
rect 5396 6667 5448 6719
rect 5461 6667 5513 6719
rect 5526 6667 5578 6719
rect 5591 6702 9099 6742
rect 5591 6668 5625 6702
rect 5625 6701 6215 6702
rect 5625 6668 5903 6701
rect 5591 6667 5903 6668
rect 5903 6667 5937 6701
rect 5937 6668 6215 6701
rect 6215 6668 6249 6702
rect 6249 6701 6839 6702
rect 6249 6668 6527 6701
rect 5937 6667 6527 6668
rect 6527 6667 6561 6701
rect 6561 6668 6839 6701
rect 6839 6668 6873 6702
rect 6873 6701 7463 6702
rect 6873 6668 7151 6701
rect 6561 6667 7151 6668
rect 7151 6667 7185 6701
rect 7185 6668 7463 6701
rect 7463 6668 7497 6702
rect 7497 6701 8399 6702
rect 7497 6668 7775 6701
rect 7185 6667 7775 6668
rect 7775 6667 7809 6701
rect 7809 6667 8087 6701
rect 8087 6667 8121 6701
rect 8121 6668 8399 6701
rect 8399 6668 8433 6702
rect 8433 6701 9023 6702
rect 8433 6668 8711 6701
rect 8121 6667 8711 6668
rect 8711 6667 8745 6701
rect 8745 6668 9023 6701
rect 9023 6668 9057 6702
rect 9057 6668 9099 6702
rect 8745 6667 9099 6668
rect 3857 6538 3875 6570
rect 3875 6538 3909 6570
rect 3857 6518 3909 6538
rect 3981 6518 4033 6570
rect 8941 6526 8993 6578
rect 9011 6526 9063 6578
rect 3857 6466 3875 6500
rect 3875 6466 3909 6500
rect 3857 6448 3909 6466
rect 3981 6448 4033 6500
rect 8941 6462 8993 6514
rect 9011 6462 9063 6514
rect 3857 6427 3909 6430
rect 3857 6393 3875 6427
rect 3875 6393 3909 6427
rect 3857 6378 3909 6393
rect 3981 6378 4033 6430
rect 8941 6398 8993 6450
rect 9011 6398 9063 6450
rect 3857 6354 3909 6359
rect 3857 6320 3875 6354
rect 3875 6320 3909 6354
rect 3857 6307 3909 6320
rect 3981 6307 4033 6359
rect 8941 6334 8993 6386
rect 9011 6334 9063 6386
rect 3857 6281 3909 6288
rect 3857 6247 3875 6281
rect 3875 6247 3909 6281
rect 3857 6236 3909 6247
rect 3981 6236 4033 6288
rect 8941 6270 8993 6322
rect 9011 6270 9063 6322
rect 3857 6208 3909 6217
rect 3857 6174 3875 6208
rect 3875 6174 3909 6208
rect 3857 6165 3909 6174
rect 3981 6165 4033 6217
rect 8941 6206 8993 6258
rect 9011 6206 9063 6258
rect 3857 6135 3909 6146
rect 3857 6101 3875 6135
rect 3875 6101 3909 6135
rect 3857 6094 3909 6101
rect 3981 6094 4033 6146
rect 8941 6142 8993 6194
rect 9011 6142 9063 6194
rect 8941 6078 8993 6130
rect 9011 6078 9063 6130
rect 3857 6062 3909 6075
rect 3857 6028 3875 6062
rect 3875 6028 3909 6062
rect 3857 6023 3909 6028
rect 3981 6023 4033 6075
rect 8941 6013 8993 6065
rect 9011 6013 9063 6065
rect 3857 5989 3909 6004
rect 3857 5955 3875 5989
rect 3875 5955 3909 5989
rect 3857 5952 3909 5955
rect 3981 5952 4033 6004
rect 8941 5948 8993 6000
rect 9011 5948 9063 6000
rect 749 5801 770 5825
rect 770 5801 801 5825
rect 631 5753 683 5792
rect 631 5747 660 5753
rect 660 5747 683 5753
rect 631 5719 660 5734
rect 660 5719 683 5734
rect 749 5752 801 5788
rect 749 5736 770 5752
rect 770 5736 801 5752
rect 631 5682 683 5719
rect 749 5718 770 5723
rect 770 5718 801 5723
rect 631 5646 660 5669
rect 660 5646 683 5669
rect 749 5679 801 5718
rect 749 5671 770 5679
rect 770 5671 801 5679
rect 631 5617 683 5646
rect 749 5645 770 5658
rect 770 5645 801 5658
rect 10677 7698 10729 7750
rect 10677 7634 10729 7686
rect 10934 7858 10986 7864
rect 10934 7824 10939 7858
rect 10939 7824 10973 7858
rect 10973 7824 10986 7858
rect 10934 7812 10986 7824
rect 11000 7812 11052 7864
rect 11066 7812 11118 7864
rect 11132 7812 11184 7864
rect 11198 7812 11250 7864
rect 11264 7858 11316 7864
rect 11264 7824 11285 7858
rect 11285 7824 11316 7858
rect 11264 7812 11316 7824
rect 11330 7812 11382 7864
rect 10934 7785 10986 7793
rect 10934 7751 10939 7785
rect 10939 7751 10973 7785
rect 10973 7751 10986 7785
rect 10934 7741 10986 7751
rect 11000 7741 11052 7793
rect 11066 7741 11118 7793
rect 11132 7741 11184 7793
rect 11198 7741 11250 7793
rect 11264 7785 11316 7793
rect 11264 7751 11285 7785
rect 11285 7751 11316 7785
rect 11264 7741 11316 7751
rect 11330 7741 11382 7793
rect 10934 7712 10986 7722
rect 10934 7678 10939 7712
rect 10939 7678 10973 7712
rect 10973 7678 10986 7712
rect 10934 7670 10986 7678
rect 11000 7670 11052 7722
rect 11066 7670 11118 7722
rect 11132 7670 11184 7722
rect 11198 7670 11250 7722
rect 11264 7712 11316 7722
rect 11264 7678 11285 7712
rect 11285 7678 11316 7712
rect 11264 7670 11316 7678
rect 11330 7670 11382 7722
rect 10934 7639 10986 7651
rect 10934 7605 10939 7639
rect 10939 7605 10973 7639
rect 10973 7605 10986 7639
rect 10934 7599 10986 7605
rect 11000 7599 11052 7651
rect 11066 7599 11118 7651
rect 11132 7599 11184 7651
rect 11198 7599 11250 7651
rect 11264 7639 11316 7651
rect 11264 7605 11285 7639
rect 11285 7605 11316 7639
rect 11264 7599 11316 7605
rect 11330 7599 11382 7651
rect 10934 7566 10986 7579
rect 10934 7532 10939 7566
rect 10939 7532 10973 7566
rect 10973 7532 10986 7566
rect 10934 7527 10986 7532
rect 11000 7527 11052 7579
rect 11066 7527 11118 7579
rect 11132 7527 11184 7579
rect 11198 7527 11250 7579
rect 11264 7566 11316 7579
rect 11264 7532 11285 7566
rect 11285 7532 11316 7566
rect 11264 7527 11316 7532
rect 11330 7527 11382 7579
rect 10934 7493 10986 7507
rect 10934 7459 10939 7493
rect 10939 7459 10973 7493
rect 10973 7459 10986 7493
rect 10934 7455 10986 7459
rect 11000 7455 11052 7507
rect 11066 7455 11118 7507
rect 11132 7455 11184 7507
rect 11198 7455 11250 7507
rect 11264 7493 11316 7507
rect 11264 7459 11285 7493
rect 11285 7459 11316 7493
rect 11264 7455 11316 7459
rect 11330 7455 11382 7507
rect 10934 7420 10986 7435
rect 10934 7386 10939 7420
rect 10939 7386 10973 7420
rect 10973 7386 10986 7420
rect 10934 7383 10986 7386
rect 11000 7383 11052 7435
rect 11066 7383 11118 7435
rect 11132 7383 11184 7435
rect 11198 7383 11250 7435
rect 11264 7420 11316 7435
rect 11264 7386 11285 7420
rect 11285 7386 11316 7420
rect 11264 7383 11316 7386
rect 11330 7383 11382 7435
rect 10934 7346 10986 7363
rect 10934 7312 10939 7346
rect 10939 7312 10973 7346
rect 10973 7312 10986 7346
rect 10934 7311 10986 7312
rect 11000 7311 11052 7363
rect 11066 7311 11118 7363
rect 11132 7311 11184 7363
rect 11198 7311 11250 7363
rect 11264 7346 11316 7363
rect 11264 7312 11285 7346
rect 11285 7312 11316 7346
rect 11264 7311 11316 7312
rect 11330 7311 11382 7363
rect 10934 7272 10986 7291
rect 10934 7239 10939 7272
rect 10939 7239 10973 7272
rect 10973 7239 10986 7272
rect 11000 7239 11052 7291
rect 11066 7239 11118 7291
rect 11132 7239 11184 7291
rect 11198 7239 11250 7291
rect 11264 7272 11316 7291
rect 11264 7239 11285 7272
rect 11285 7239 11316 7272
rect 11330 7239 11382 7291
rect 10985 7108 11037 7160
rect 11111 7154 11163 7160
rect 11111 7120 11127 7154
rect 11127 7120 11163 7154
rect 11111 7108 11163 7120
rect 10985 7043 11037 7095
rect 11111 7080 11163 7095
rect 11111 7046 11127 7080
rect 11127 7046 11163 7080
rect 11111 7043 11163 7046
rect 10985 6978 11037 7030
rect 11111 7006 11163 7030
rect 11111 6978 11127 7006
rect 11127 6978 11163 7006
rect 10985 6913 11037 6965
rect 11111 6932 11163 6965
rect 11111 6913 11127 6932
rect 11127 6913 11163 6932
rect 10985 6847 11037 6899
rect 11111 6898 11127 6899
rect 11127 6898 11163 6899
rect 11111 6858 11163 6898
rect 11111 6847 11127 6858
rect 11127 6847 11163 6858
rect 10985 6781 11037 6833
rect 11111 6824 11127 6833
rect 11127 6824 11163 6833
rect 11111 6783 11163 6824
rect 11111 6781 11127 6783
rect 11127 6781 11163 6783
rect 10985 6715 11037 6767
rect 11111 6749 11127 6767
rect 11127 6749 11163 6767
rect 11111 6715 11163 6749
rect 10985 6649 11037 6701
rect 11111 6674 11127 6701
rect 11127 6674 11163 6701
rect 11111 6649 11163 6674
rect 10985 6583 11037 6635
rect 11111 6633 11163 6635
rect 11111 6599 11127 6633
rect 11127 6599 11163 6633
rect 11111 6583 11163 6599
rect 10985 6517 11037 6569
rect 11111 6558 11163 6569
rect 11111 6524 11127 6558
rect 11127 6524 11163 6558
rect 11111 6517 11163 6524
rect 631 5573 660 5604
rect 660 5573 683 5604
rect 749 5606 801 5645
rect 631 5552 683 5573
rect 749 5541 770 5593
rect 770 5541 801 5593
rect 813 5541 865 5593
rect 877 5541 929 5593
rect 941 5541 993 5593
rect 1005 5541 1057 5593
rect 1069 5541 1121 5593
rect 1133 5541 1185 5593
rect 1197 5541 1249 5593
rect 1261 5541 1313 5593
rect 1325 5541 1377 5593
rect 1389 5541 1441 5593
rect 1453 5541 1505 5593
rect 1517 5541 1569 5593
rect 1581 5541 1633 5593
rect 1646 5541 1698 5593
rect 1711 5541 1763 5593
rect 1776 5541 1828 5593
rect 1841 5541 1893 5593
rect 1906 5541 1958 5593
rect 1971 5541 2023 5593
rect 2036 5541 2088 5593
rect 2101 5541 2153 5593
rect 2166 5541 2218 5593
rect 631 5534 683 5539
rect 631 5500 660 5534
rect 660 5500 683 5534
rect 631 5487 683 5500
rect 697 5428 698 5475
rect 698 5428 749 5475
rect 763 5428 815 5475
rect 829 5428 881 5475
rect 895 5428 947 5475
rect 961 5428 1013 5475
rect 1027 5428 1079 5475
rect 1094 5428 1146 5475
rect 1161 5428 1213 5475
rect 1228 5428 1280 5475
rect 1295 5428 1347 5475
rect 1362 5428 1414 5475
rect 1429 5428 1481 5475
rect 1496 5428 1548 5475
rect 1563 5428 1615 5475
rect 1630 5428 1682 5475
rect 1697 5428 1749 5475
rect 1764 5428 1816 5475
rect 1831 5428 1883 5475
rect 1898 5428 1950 5475
rect 1965 5428 2017 5475
rect 2032 5428 2084 5475
rect 2099 5428 2151 5475
rect 2166 5428 2218 5475
rect 697 5423 749 5428
rect 763 5423 815 5428
rect 829 5423 881 5428
rect 895 5423 947 5428
rect 961 5423 1013 5428
rect 1027 5423 1079 5428
rect 1094 5423 1146 5428
rect 1161 5423 1213 5428
rect 1228 5423 1280 5428
rect 1295 5423 1347 5428
rect 1362 5423 1414 5428
rect 1429 5423 1481 5428
rect 1496 5423 1548 5428
rect 1563 5423 1615 5428
rect 1630 5423 1682 5428
rect 1697 5423 1749 5428
rect 1764 5423 1816 5428
rect 1831 5423 1883 5428
rect 1898 5423 1950 5428
rect 1965 5423 2017 5428
rect 2032 5423 2084 5428
rect 2099 5423 2151 5428
rect 2166 5423 2218 5428
rect 3854 5313 3906 5365
rect 3918 5313 3970 5365
rect 3982 5313 4034 5365
rect 2771 3952 2823 4004
rect 2838 3952 2890 4004
rect 2905 3952 2957 4004
rect 2972 3952 3024 4004
rect 3039 3952 3091 4004
rect 3106 3952 3158 4004
rect 3173 3952 3225 4004
rect 3240 3952 3292 4004
rect 3307 3952 3359 4004
rect 3374 3952 3426 4004
rect 3441 3952 3493 4004
rect 3508 3952 3560 4004
rect 3575 3952 3627 4004
rect 3642 3952 3694 4004
rect 3708 3952 3760 4004
rect 3774 3952 3826 4004
rect 2771 3884 2823 3936
rect 2838 3884 2890 3936
rect 2905 3884 2957 3936
rect 2972 3884 3024 3936
rect 3039 3884 3091 3936
rect 3106 3884 3158 3936
rect 3173 3884 3225 3936
rect 3240 3884 3292 3936
rect 3307 3884 3359 3936
rect 3374 3884 3426 3936
rect 3441 3884 3493 3936
rect 3508 3884 3560 3936
rect 3575 3884 3627 3936
rect 3642 3884 3694 3936
rect 3708 3884 3760 3936
rect 3774 3884 3826 3936
rect 2771 3816 2823 3868
rect 2838 3816 2890 3868
rect 2905 3816 2957 3868
rect 2972 3816 3024 3868
rect 3039 3816 3091 3868
rect 3106 3816 3158 3868
rect 3173 3816 3225 3868
rect 3240 3816 3292 3868
rect 3307 3816 3359 3868
rect 3374 3816 3426 3868
rect 3441 3816 3493 3868
rect 3508 3816 3560 3868
rect 3575 3816 3627 3868
rect 3642 3816 3694 3868
rect 3708 3816 3760 3868
rect 3774 3816 3826 3868
rect 2771 3748 2823 3800
rect 2838 3748 2890 3800
rect 2905 3748 2957 3800
rect 2972 3748 3024 3800
rect 3039 3748 3091 3800
rect 3106 3748 3158 3800
rect 3173 3748 3225 3800
rect 3240 3748 3292 3800
rect 3307 3748 3359 3800
rect 3374 3748 3426 3800
rect 3441 3748 3493 3800
rect 3508 3748 3560 3800
rect 3575 3748 3627 3800
rect 3642 3748 3694 3800
rect 3708 3748 3760 3800
rect 3774 3748 3826 3800
rect 2771 3680 2823 3732
rect 2838 3680 2890 3732
rect 2905 3680 2957 3732
rect 2972 3680 3024 3732
rect 3039 3680 3091 3732
rect 3106 3680 3158 3732
rect 3173 3680 3225 3732
rect 3240 3680 3292 3732
rect 3307 3680 3359 3732
rect 3374 3680 3426 3732
rect 3441 3680 3493 3732
rect 3508 3680 3560 3732
rect 3575 3680 3627 3732
rect 3642 3680 3694 3732
rect 3708 3680 3760 3732
rect 3774 3680 3826 3732
rect 2771 3612 2823 3664
rect 2838 3612 2890 3664
rect 2905 3612 2957 3664
rect 2972 3612 3024 3664
rect 3039 3612 3091 3664
rect 3106 3612 3158 3664
rect 3173 3612 3225 3664
rect 3240 3612 3292 3664
rect 3307 3612 3359 3664
rect 3374 3612 3426 3664
rect 3441 3612 3493 3664
rect 3508 3612 3560 3664
rect 3575 3612 3627 3664
rect 3642 3612 3694 3664
rect 3708 3612 3760 3664
rect 3774 3612 3826 3664
rect 2771 3544 2823 3596
rect 2838 3544 2890 3596
rect 2905 3544 2957 3596
rect 2972 3544 3024 3596
rect 3039 3544 3091 3596
rect 3106 3544 3158 3596
rect 3173 3544 3225 3596
rect 3240 3544 3292 3596
rect 3307 3544 3359 3596
rect 3374 3544 3426 3596
rect 3441 3544 3493 3596
rect 3508 3544 3560 3596
rect 3575 3544 3627 3596
rect 3642 3544 3694 3596
rect 3708 3544 3760 3596
rect 3774 3544 3826 3596
rect 2771 3476 2823 3528
rect 2838 3476 2890 3528
rect 2905 3476 2957 3528
rect 2972 3476 3024 3528
rect 3039 3476 3091 3528
rect 3106 3476 3158 3528
rect 3173 3476 3225 3528
rect 3240 3476 3292 3528
rect 3307 3476 3359 3528
rect 3374 3476 3426 3528
rect 3441 3476 3493 3528
rect 3508 3476 3560 3528
rect 3575 3476 3627 3528
rect 3642 3476 3694 3528
rect 3708 3476 3760 3528
rect 3774 3476 3826 3528
rect 2766 2740 2818 2792
rect 2831 2740 2883 2792
rect 2896 2740 2948 2792
rect 2961 2740 3013 2792
rect 3026 2740 3078 2792
rect 3091 2740 3143 2792
rect 3156 2740 3208 2792
rect 3221 2740 3273 2792
rect 3285 2740 3337 2792
rect 3349 2740 3401 2792
rect 3413 2740 3465 2792
rect 3477 2740 3529 2792
rect 3541 2740 3593 2792
rect 3605 2740 3657 2792
rect 3669 2740 3721 2792
rect 3733 2740 3785 2792
rect 3797 2740 3849 2792
rect 3861 2740 3913 2792
rect 3925 2740 3977 2792
rect 3989 2740 4041 2792
rect 4053 2740 4105 2792
rect 4117 2740 4169 2792
rect 4181 2740 4233 2792
rect 4245 2740 4297 2792
rect 4309 2740 4361 2792
rect 4373 2740 4425 2792
rect 4437 2740 4489 2792
rect 4501 2740 4553 2792
rect 4565 2740 4617 2792
rect 4629 2740 4681 2792
rect 4693 2740 4745 2792
rect 4757 2740 4809 2792
rect 4821 2740 4873 2792
rect 2766 2674 2818 2726
rect 2831 2674 2883 2726
rect 2896 2674 2948 2726
rect 2961 2674 3013 2726
rect 3026 2674 3078 2726
rect 3091 2674 3143 2726
rect 3156 2674 3208 2726
rect 3221 2674 3273 2726
rect 3285 2674 3337 2726
rect 3349 2674 3401 2726
rect 3413 2674 3465 2726
rect 3477 2674 3529 2726
rect 3541 2674 3593 2726
rect 3605 2674 3657 2726
rect 3669 2674 3721 2726
rect 3733 2674 3785 2726
rect 3797 2674 3849 2726
rect 3861 2674 3913 2726
rect 3925 2674 3977 2726
rect 3989 2674 4041 2726
rect 4053 2674 4105 2726
rect 4117 2674 4169 2726
rect 4181 2674 4233 2726
rect 4245 2674 4297 2726
rect 4309 2674 4361 2726
rect 4373 2674 4425 2726
rect 4437 2674 4489 2726
rect 4501 2674 4553 2726
rect 4565 2674 4617 2726
rect 4629 2674 4681 2726
rect 4693 2674 4745 2726
rect 4757 2674 4809 2726
rect 4821 2674 4873 2726
rect 2766 2608 2818 2660
rect 2831 2608 2883 2660
rect 2896 2608 2948 2660
rect 2961 2608 3013 2660
rect 3026 2608 3078 2660
rect 3091 2608 3143 2660
rect 3156 2608 3208 2660
rect 3221 2608 3273 2660
rect 3285 2608 3337 2660
rect 3349 2608 3401 2660
rect 3413 2608 3465 2660
rect 3477 2608 3529 2660
rect 3541 2608 3593 2660
rect 3605 2608 3657 2660
rect 3669 2608 3721 2660
rect 3733 2608 3785 2660
rect 3797 2608 3849 2660
rect 3861 2608 3913 2660
rect 3925 2608 3977 2660
rect 3989 2608 4041 2660
rect 4053 2608 4105 2660
rect 4117 2608 4169 2660
rect 4181 2608 4233 2660
rect 4245 2608 4297 2660
rect 4309 2608 4361 2660
rect 4373 2608 4425 2660
rect 4437 2608 4489 2660
rect 4501 2608 4553 2660
rect 4565 2608 4617 2660
rect 4629 2608 4681 2660
rect 4693 2608 4745 2660
rect 4757 2608 4809 2660
rect 4821 2608 4873 2660
rect 2766 2542 2818 2594
rect 2831 2542 2883 2594
rect 2896 2542 2948 2594
rect 2961 2542 3013 2594
rect 3026 2542 3078 2594
rect 3091 2542 3143 2594
rect 3156 2542 3208 2594
rect 3221 2542 3273 2594
rect 3285 2542 3337 2594
rect 3349 2542 3401 2594
rect 3413 2542 3465 2594
rect 3477 2542 3529 2594
rect 3541 2542 3593 2594
rect 3605 2542 3657 2594
rect 3669 2542 3721 2594
rect 3733 2542 3785 2594
rect 3797 2542 3849 2594
rect 3861 2542 3913 2594
rect 3925 2542 3977 2594
rect 3989 2542 4041 2594
rect 4053 2542 4105 2594
rect 4117 2542 4169 2594
rect 4181 2542 4233 2594
rect 4245 2542 4297 2594
rect 4309 2542 4361 2594
rect 4373 2542 4425 2594
rect 4437 2542 4489 2594
rect 4501 2542 4553 2594
rect 4565 2542 4617 2594
rect 4629 2542 4681 2594
rect 4693 2542 4745 2594
rect 4757 2542 4809 2594
rect 4821 2542 4873 2594
rect 2766 2476 2818 2528
rect 2831 2476 2883 2528
rect 2896 2476 2948 2528
rect 2961 2476 3013 2528
rect 3026 2476 3078 2528
rect 3091 2476 3143 2528
rect 3156 2476 3208 2528
rect 3221 2476 3273 2528
rect 3285 2476 3337 2528
rect 3349 2476 3401 2528
rect 3413 2476 3465 2528
rect 3477 2476 3529 2528
rect 3541 2476 3593 2528
rect 3605 2476 3657 2528
rect 3669 2476 3721 2528
rect 3733 2476 3785 2528
rect 3797 2476 3849 2528
rect 3861 2476 3913 2528
rect 3925 2476 3977 2528
rect 3989 2476 4041 2528
rect 4053 2476 4105 2528
rect 4117 2476 4169 2528
rect 4181 2476 4233 2528
rect 4245 2476 4297 2528
rect 4309 2476 4361 2528
rect 4373 2476 4425 2528
rect 4437 2476 4489 2528
rect 4501 2476 4553 2528
rect 4565 2476 4617 2528
rect 4629 2476 4681 2528
rect 4693 2476 4745 2528
rect 4757 2476 4809 2528
rect 4821 2476 4873 2528
rect 2766 2410 2818 2462
rect 2831 2410 2883 2462
rect 2896 2410 2948 2462
rect 2961 2410 3013 2462
rect 3026 2410 3078 2462
rect 3091 2410 3143 2462
rect 3156 2410 3208 2462
rect 3221 2410 3273 2462
rect 3285 2410 3337 2462
rect 3349 2410 3401 2462
rect 3413 2410 3465 2462
rect 3477 2410 3529 2462
rect 3541 2410 3593 2462
rect 3605 2410 3657 2462
rect 3669 2410 3721 2462
rect 3733 2410 3785 2462
rect 3797 2410 3849 2462
rect 3861 2410 3913 2462
rect 3925 2410 3977 2462
rect 3989 2410 4041 2462
rect 4053 2410 4105 2462
rect 4117 2410 4169 2462
rect 4181 2410 4233 2462
rect 4245 2410 4297 2462
rect 4309 2410 4361 2462
rect 4373 2410 4425 2462
rect 4437 2410 4489 2462
rect 4501 2410 4553 2462
rect 4565 2410 4617 2462
rect 4629 2410 4681 2462
rect 4693 2410 4745 2462
rect 4757 2410 4809 2462
rect 4821 2410 4873 2462
rect 2766 2344 2818 2396
rect 2831 2344 2883 2396
rect 2896 2344 2948 2396
rect 2961 2344 3013 2396
rect 3026 2344 3078 2396
rect 3091 2344 3143 2396
rect 3156 2344 3208 2396
rect 3221 2344 3273 2396
rect 3285 2344 3337 2396
rect 3349 2344 3401 2396
rect 3413 2344 3465 2396
rect 3477 2344 3529 2396
rect 3541 2344 3593 2396
rect 3605 2344 3657 2396
rect 3669 2344 3721 2396
rect 3733 2344 3785 2396
rect 3797 2344 3849 2396
rect 3861 2344 3913 2396
rect 3925 2344 3977 2396
rect 3989 2344 4041 2396
rect 4053 2344 4105 2396
rect 4117 2344 4169 2396
rect 4181 2344 4233 2396
rect 4245 2344 4297 2396
rect 4309 2344 4361 2396
rect 4373 2344 4425 2396
rect 4437 2344 4489 2396
rect 4501 2344 4553 2396
rect 4565 2344 4617 2396
rect 4629 2344 4681 2396
rect 4693 2344 4745 2396
rect 4757 2344 4809 2396
rect 4821 2344 4873 2396
rect 2766 2278 2818 2330
rect 2831 2278 2883 2330
rect 2896 2278 2948 2330
rect 2961 2278 3013 2330
rect 3026 2278 3078 2330
rect 3091 2278 3143 2330
rect 3156 2278 3208 2330
rect 3221 2278 3273 2330
rect 3285 2278 3337 2330
rect 3349 2278 3401 2330
rect 3413 2278 3465 2330
rect 3477 2278 3529 2330
rect 3541 2278 3593 2330
rect 3605 2278 3657 2330
rect 3669 2278 3721 2330
rect 3733 2278 3785 2330
rect 3797 2278 3849 2330
rect 3861 2278 3913 2330
rect 3925 2278 3977 2330
rect 3989 2278 4041 2330
rect 4053 2278 4105 2330
rect 4117 2278 4169 2330
rect 4181 2278 4233 2330
rect 4245 2278 4297 2330
rect 4309 2278 4361 2330
rect 4373 2278 4425 2330
rect 4437 2278 4489 2330
rect 4501 2278 4553 2330
rect 4565 2278 4617 2330
rect 4629 2278 4681 2330
rect 4693 2278 4745 2330
rect 4757 2278 4809 2330
rect 4821 2278 4873 2330
rect 2766 2212 2818 2264
rect 2831 2212 2883 2264
rect 2896 2212 2948 2264
rect 2961 2212 3013 2264
rect 3026 2212 3078 2264
rect 3091 2212 3143 2264
rect 3156 2212 3208 2264
rect 3221 2212 3273 2264
rect 3285 2212 3337 2264
rect 3349 2212 3401 2264
rect 3413 2212 3465 2264
rect 3477 2212 3529 2264
rect 3541 2212 3593 2264
rect 3605 2212 3657 2264
rect 3669 2212 3721 2264
rect 3733 2212 3785 2264
rect 3797 2212 3849 2264
rect 3861 2212 3913 2264
rect 3925 2212 3977 2264
rect 3989 2212 4041 2264
rect 4053 2212 4105 2264
rect 4117 2212 4169 2264
rect 4181 2212 4233 2264
rect 4245 2212 4297 2264
rect 4309 2212 4361 2264
rect 4373 2212 4425 2264
rect 4437 2212 4489 2264
rect 4501 2212 4553 2264
rect 4565 2212 4617 2264
rect 4629 2212 4681 2264
rect 4693 2212 4745 2264
rect 4757 2212 4809 2264
rect 4821 2212 4873 2264
rect 2776 1461 2828 1513
rect 2842 1461 2894 1513
rect 2908 1461 2960 1513
rect 2974 1461 3026 1513
rect 3040 1461 3092 1513
rect 3106 1461 3158 1513
rect 3172 1461 3224 1513
rect 3238 1461 3290 1513
rect 3304 1461 3356 1513
rect 3370 1461 3422 1513
rect 3436 1461 3488 1513
rect 3502 1461 3554 1513
rect 3568 1461 3620 1513
rect 3634 1461 3686 1513
rect 3700 1461 3752 1513
rect 3766 1461 3818 1513
rect 3832 1461 3884 1513
rect 3898 1461 3950 1513
rect 3964 1461 4016 1513
rect 4030 1461 4082 1513
rect 4096 1461 4148 1513
rect 4162 1461 4214 1513
rect 4228 1461 4280 1513
rect 4294 1461 4346 1513
rect 4360 1461 4412 1513
rect 4426 1461 4478 1513
rect 4492 1461 4544 1513
rect 4558 1461 4610 1513
rect 4624 1461 4676 1513
rect 4690 1461 4742 1513
rect 4756 1461 4808 1513
rect 4821 1461 4873 1513
rect 2776 1393 2828 1445
rect 2842 1393 2894 1445
rect 2908 1393 2960 1445
rect 2974 1393 3026 1445
rect 3040 1393 3092 1445
rect 3106 1393 3158 1445
rect 3172 1393 3224 1445
rect 3238 1393 3290 1445
rect 3304 1393 3356 1445
rect 3370 1393 3422 1445
rect 3436 1393 3488 1445
rect 3502 1393 3554 1445
rect 3568 1393 3620 1445
rect 3634 1393 3686 1445
rect 3700 1393 3752 1445
rect 3766 1393 3818 1445
rect 3832 1393 3884 1445
rect 3898 1393 3950 1445
rect 3964 1393 4016 1445
rect 4030 1393 4082 1445
rect 4096 1393 4148 1445
rect 4162 1393 4214 1445
rect 4228 1393 4280 1445
rect 4294 1393 4346 1445
rect 4360 1393 4412 1445
rect 4426 1393 4478 1445
rect 4492 1393 4544 1445
rect 4558 1393 4610 1445
rect 4624 1393 4676 1445
rect 4690 1393 4742 1445
rect 4756 1393 4808 1445
rect 4821 1393 4873 1445
rect 2776 1325 2828 1377
rect 2842 1325 2894 1377
rect 2908 1325 2960 1377
rect 2974 1325 3026 1377
rect 3040 1325 3092 1377
rect 3106 1325 3158 1377
rect 3172 1325 3224 1377
rect 3238 1325 3290 1377
rect 3304 1325 3356 1377
rect 3370 1325 3422 1377
rect 3436 1325 3488 1377
rect 3502 1325 3554 1377
rect 3568 1325 3620 1377
rect 3634 1325 3686 1377
rect 3700 1325 3752 1377
rect 3766 1325 3818 1377
rect 3832 1325 3884 1377
rect 3898 1325 3950 1377
rect 3964 1325 4016 1377
rect 4030 1325 4082 1377
rect 4096 1325 4148 1377
rect 4162 1325 4214 1377
rect 4228 1325 4280 1377
rect 4294 1325 4346 1377
rect 4360 1325 4412 1377
rect 4426 1325 4478 1377
rect 4492 1325 4544 1377
rect 4558 1325 4610 1377
rect 4624 1325 4676 1377
rect 4690 1325 4742 1377
rect 4756 1325 4808 1377
rect 4821 1325 4873 1377
rect 2776 1257 2828 1309
rect 2842 1257 2894 1309
rect 2908 1257 2960 1309
rect 2974 1257 3026 1309
rect 3040 1257 3092 1309
rect 3106 1257 3158 1309
rect 3172 1257 3224 1309
rect 3238 1257 3290 1309
rect 3304 1257 3356 1309
rect 3370 1257 3422 1309
rect 3436 1257 3488 1309
rect 3502 1257 3554 1309
rect 3568 1257 3620 1309
rect 3634 1257 3686 1309
rect 3700 1257 3752 1309
rect 3766 1257 3818 1309
rect 3832 1257 3884 1309
rect 3898 1257 3950 1309
rect 3964 1257 4016 1309
rect 4030 1257 4082 1309
rect 4096 1257 4148 1309
rect 4162 1257 4214 1309
rect 4228 1257 4280 1309
rect 4294 1257 4346 1309
rect 4360 1257 4412 1309
rect 4426 1257 4478 1309
rect 4492 1257 4544 1309
rect 4558 1257 4610 1309
rect 4624 1257 4676 1309
rect 4690 1257 4742 1309
rect 4756 1257 4808 1309
rect 4821 1257 4873 1309
rect 2776 1189 2828 1241
rect 2842 1189 2894 1241
rect 2908 1189 2960 1241
rect 2974 1189 3026 1241
rect 3040 1189 3092 1241
rect 3106 1189 3158 1241
rect 3172 1189 3224 1241
rect 3238 1189 3290 1241
rect 3304 1189 3356 1241
rect 3370 1189 3422 1241
rect 3436 1189 3488 1241
rect 3502 1189 3554 1241
rect 3568 1189 3620 1241
rect 3634 1189 3686 1241
rect 3700 1189 3752 1241
rect 3766 1189 3818 1241
rect 3832 1189 3884 1241
rect 3898 1189 3950 1241
rect 3964 1189 4016 1241
rect 4030 1189 4082 1241
rect 4096 1189 4148 1241
rect 4162 1189 4214 1241
rect 4228 1189 4280 1241
rect 4294 1189 4346 1241
rect 4360 1189 4412 1241
rect 4426 1189 4478 1241
rect 4492 1189 4544 1241
rect 4558 1189 4610 1241
rect 4624 1189 4676 1241
rect 4690 1189 4742 1241
rect 4756 1189 4808 1241
rect 4821 1189 4873 1241
rect 2776 1121 2828 1173
rect 2842 1121 2894 1173
rect 2908 1121 2960 1173
rect 2974 1121 3026 1173
rect 3040 1121 3092 1173
rect 3106 1121 3158 1173
rect 3172 1121 3224 1173
rect 3238 1121 3290 1173
rect 3304 1121 3356 1173
rect 3370 1121 3422 1173
rect 3436 1121 3488 1173
rect 3502 1121 3554 1173
rect 3568 1121 3620 1173
rect 3634 1121 3686 1173
rect 3700 1121 3752 1173
rect 3766 1121 3818 1173
rect 3832 1121 3884 1173
rect 3898 1121 3950 1173
rect 3964 1121 4016 1173
rect 4030 1121 4082 1173
rect 4096 1121 4148 1173
rect 4162 1121 4214 1173
rect 4228 1121 4280 1173
rect 4294 1121 4346 1173
rect 4360 1121 4412 1173
rect 4426 1121 4478 1173
rect 4492 1121 4544 1173
rect 4558 1121 4610 1173
rect 4624 1121 4676 1173
rect 4690 1121 4742 1173
rect 4756 1121 4808 1173
rect 4821 1121 4873 1173
rect 2776 1053 2828 1105
rect 2842 1053 2894 1105
rect 2908 1053 2960 1105
rect 2974 1053 3026 1105
rect 3040 1053 3092 1105
rect 3106 1053 3158 1105
rect 3172 1053 3224 1105
rect 3238 1053 3290 1105
rect 3304 1053 3356 1105
rect 3370 1053 3422 1105
rect 3436 1053 3488 1105
rect 3502 1053 3554 1105
rect 3568 1053 3620 1105
rect 3634 1053 3686 1105
rect 3700 1053 3752 1105
rect 3766 1053 3818 1105
rect 3832 1053 3884 1105
rect 3898 1053 3950 1105
rect 3964 1053 4016 1105
rect 4030 1053 4082 1105
rect 4096 1053 4148 1105
rect 4162 1053 4214 1105
rect 4228 1053 4280 1105
rect 4294 1053 4346 1105
rect 4360 1053 4412 1105
rect 4426 1053 4478 1105
rect 4492 1053 4544 1105
rect 4558 1053 4610 1105
rect 4624 1053 4676 1105
rect 4690 1053 4742 1105
rect 4756 1053 4808 1105
rect 4821 1053 4873 1105
rect 2776 985 2828 1037
rect 2842 985 2894 1037
rect 2908 985 2960 1037
rect 2974 985 3026 1037
rect 3040 985 3092 1037
rect 3106 985 3158 1037
rect 3172 985 3224 1037
rect 3238 985 3290 1037
rect 3304 985 3356 1037
rect 3370 985 3422 1037
rect 3436 985 3488 1037
rect 3502 985 3554 1037
rect 3568 985 3620 1037
rect 3634 985 3686 1037
rect 3700 985 3752 1037
rect 3766 985 3818 1037
rect 3832 985 3884 1037
rect 3898 985 3950 1037
rect 3964 985 4016 1037
rect 4030 985 4082 1037
rect 4096 985 4148 1037
rect 4162 985 4214 1037
rect 4228 985 4280 1037
rect 4294 985 4346 1037
rect 4360 985 4412 1037
rect 4426 985 4478 1037
rect 4492 985 4544 1037
rect 4558 985 4610 1037
rect 4624 985 4676 1037
rect 4690 985 4742 1037
rect 4756 985 4808 1037
rect 4821 985 4873 1037
rect 6749 1054 6801 1106
rect 6749 970 6801 1022
rect 8703 1054 8755 1106
rect 8703 970 8755 1022
rect 6707 515 6759 567
rect 6791 515 6843 567
rect 8661 515 8713 567
rect 8745 515 8797 567
rect 5190 325 5242 377
rect 5256 325 5308 377
rect 5322 325 5374 377
rect 5388 325 5440 377
rect 5453 325 5505 377
rect 5518 325 5570 377
rect 5190 261 5242 313
rect 5256 261 5308 313
rect 5322 261 5374 313
rect 5388 261 5440 313
rect 5453 261 5505 313
rect 5518 261 5570 313
rect 5190 200 5242 249
rect 5256 200 5308 249
rect 5322 200 5374 249
rect 5388 200 5440 249
rect 5453 200 5505 249
rect 5518 200 5570 249
rect 5190 197 5242 200
rect 5256 197 5308 200
rect 5322 197 5374 200
rect 5388 197 5440 200
rect 5453 197 5505 200
rect 5518 197 5570 200
<< metal2 >>
rect 187 39009 13440 39015
rect 187 38953 2534 39009
rect 2590 38953 2617 39009
rect 2673 38953 2700 39009
rect 2756 38953 2783 39009
rect 2839 38953 2866 39009
rect 2924 38957 2940 39009
rect 3005 38957 3008 39009
rect 2922 38953 2949 38957
rect 3005 38953 3032 38957
rect 3088 38953 3115 39009
rect 3171 38953 3198 39009
rect 3254 38953 3281 39009
rect 3337 38953 3364 39009
rect 3420 38953 3447 39009
rect 3503 38953 3530 39009
rect 3586 38953 3613 39009
rect 3669 38953 3696 39009
rect 3752 38953 3779 39009
rect 3844 38957 3860 39009
rect 3918 38957 3928 39009
rect 3835 38953 3862 38957
rect 3918 38953 3945 38957
rect 4001 38953 4028 39009
rect 4084 38953 4111 39009
rect 4167 38953 4194 39009
rect 4250 38953 4276 39009
rect 4332 38953 4358 39009
rect 4414 38953 4440 39009
rect 4496 38953 4522 39009
rect 4578 38953 4604 39009
rect 4660 38953 4686 39009
rect 4764 38957 4768 39009
rect 4832 38957 4848 39009
rect 4742 38953 4768 38957
rect 4824 38953 4850 38957
rect 4906 38953 4932 39009
rect 4988 38953 5195 39009
rect 5251 38953 5276 39009
rect 5332 38953 5357 39009
rect 5413 38953 5438 39009
rect 5494 38953 5519 39009
rect 5575 38953 5600 39009
rect 5752 38957 5762 39009
rect 5820 38957 5843 39009
rect 5656 38953 5681 38957
rect 5737 38953 5762 38957
rect 5818 38953 5843 38957
rect 5899 38953 5924 39009
rect 5980 38953 6005 39009
rect 6061 38953 6086 39009
rect 6142 38953 6167 39009
rect 6223 38953 6248 39009
rect 6304 38953 6329 39009
rect 6385 38953 6410 39009
rect 6466 38953 6491 39009
rect 6547 38957 6552 39009
rect 6547 38953 6572 38957
rect 6628 38953 6653 38957
rect 6709 38953 6734 38957
rect 6790 38953 6815 39009
rect 6871 38953 6896 39009
rect 6952 38953 6977 39009
rect 7033 38953 7058 39009
rect 7114 38953 7139 39009
rect 7195 38953 7221 39009
rect 7277 38953 7303 39009
rect 7359 38957 7472 39009
rect 7524 38957 7540 39009
rect 7592 38957 7608 39009
rect 7660 38957 8392 39009
rect 8444 38957 8460 39009
rect 8512 38957 8528 39009
rect 8580 38957 9312 39009
rect 9364 38957 9380 39009
rect 9432 38957 9448 39009
rect 9500 38957 10232 39009
rect 10284 38957 10300 39009
rect 10352 38957 10368 39009
rect 10420 38957 11152 39009
rect 11204 38957 11220 39009
rect 11272 38957 11288 39009
rect 11340 38957 12072 39009
rect 12124 38957 12140 39009
rect 12192 38957 12208 39009
rect 12260 38957 12992 39009
rect 13044 38957 13060 39009
rect 13112 38957 13128 39009
rect 13180 38957 13440 39009
rect 7359 38953 13440 38957
rect 187 38945 13440 38953
rect 187 38944 12992 38945
rect 187 38925 2872 38944
rect 187 38869 2534 38925
rect 2590 38869 2617 38925
rect 2673 38869 2700 38925
rect 2756 38869 2783 38925
rect 2839 38869 2866 38925
rect 2924 38892 2940 38944
rect 2992 38925 3008 38944
rect 3060 38925 3792 38944
rect 3005 38892 3008 38925
rect 2922 38879 2949 38892
rect 3005 38879 3032 38892
rect 187 38841 2872 38869
rect 187 38785 2534 38841
rect 2590 38785 2617 38841
rect 2673 38785 2700 38841
rect 2756 38785 2783 38841
rect 2839 38785 2866 38841
rect 2924 38827 2940 38879
rect 3005 38869 3008 38879
rect 3088 38869 3115 38925
rect 3171 38869 3198 38925
rect 3254 38869 3281 38925
rect 3337 38869 3364 38925
rect 3420 38869 3447 38925
rect 3503 38869 3530 38925
rect 3586 38869 3613 38925
rect 3669 38869 3696 38925
rect 3752 38869 3779 38925
rect 3844 38892 3860 38944
rect 3912 38925 3928 38944
rect 3980 38925 4712 38944
rect 4764 38925 4780 38944
rect 3918 38892 3928 38925
rect 3835 38879 3862 38892
rect 3918 38879 3945 38892
rect 2992 38841 3008 38869
rect 3060 38841 3792 38869
rect 3005 38827 3008 38841
rect 2922 38814 2949 38827
rect 3005 38814 3032 38827
rect 187 38762 2872 38785
rect 2924 38762 2940 38814
rect 3005 38785 3008 38814
rect 3088 38785 3115 38841
rect 3171 38785 3198 38841
rect 3254 38785 3281 38841
rect 3337 38785 3364 38841
rect 3420 38785 3447 38841
rect 3503 38785 3530 38841
rect 3586 38785 3613 38841
rect 3669 38785 3696 38841
rect 3752 38785 3779 38841
rect 3844 38827 3860 38879
rect 3918 38869 3928 38879
rect 4001 38869 4028 38925
rect 4084 38869 4111 38925
rect 4167 38869 4194 38925
rect 4250 38869 4276 38925
rect 4332 38869 4358 38925
rect 4414 38869 4440 38925
rect 4496 38869 4522 38925
rect 4578 38869 4604 38925
rect 4660 38869 4686 38925
rect 4764 38892 4768 38925
rect 4832 38892 4848 38944
rect 4900 38925 5632 38944
rect 5684 38925 5700 38944
rect 5752 38925 5768 38944
rect 5820 38925 6552 38944
rect 6604 38925 6620 38944
rect 6672 38925 6688 38944
rect 6740 38925 7472 38944
rect 4742 38879 4768 38892
rect 4824 38879 4850 38892
rect 4764 38869 4768 38879
rect 3912 38841 3928 38869
rect 3980 38841 4712 38869
rect 4764 38841 4780 38869
rect 3918 38827 3928 38841
rect 3835 38814 3862 38827
rect 3918 38814 3945 38827
rect 2992 38762 3008 38785
rect 3060 38762 3792 38785
rect 3844 38762 3860 38814
rect 3918 38785 3928 38814
rect 4001 38785 4028 38841
rect 4084 38785 4111 38841
rect 4167 38785 4194 38841
rect 4250 38785 4276 38841
rect 4332 38785 4358 38841
rect 4414 38785 4440 38841
rect 4496 38785 4522 38841
rect 4578 38785 4604 38841
rect 4660 38785 4686 38841
rect 4764 38827 4768 38841
rect 4832 38827 4848 38879
rect 4906 38869 4932 38925
rect 4988 38869 5195 38925
rect 5251 38869 5276 38925
rect 5332 38869 5357 38925
rect 5413 38869 5438 38925
rect 5494 38869 5519 38925
rect 5575 38869 5600 38925
rect 5752 38892 5762 38925
rect 5820 38892 5843 38925
rect 5656 38879 5681 38892
rect 5737 38879 5762 38892
rect 5818 38879 5843 38892
rect 5752 38869 5762 38879
rect 5820 38869 5843 38879
rect 5899 38869 5924 38925
rect 5980 38869 6005 38925
rect 6061 38869 6086 38925
rect 6142 38869 6167 38925
rect 6223 38869 6248 38925
rect 6304 38869 6329 38925
rect 6385 38869 6410 38925
rect 6466 38869 6491 38925
rect 6547 38892 6552 38925
rect 6547 38879 6572 38892
rect 6628 38879 6653 38892
rect 6709 38879 6734 38892
rect 6547 38869 6552 38879
rect 6790 38869 6815 38925
rect 6871 38869 6896 38925
rect 6952 38869 6977 38925
rect 7033 38869 7058 38925
rect 7114 38869 7139 38925
rect 7195 38869 7221 38925
rect 7277 38869 7303 38925
rect 7359 38892 7472 38925
rect 7524 38892 7540 38944
rect 7592 38892 7608 38944
rect 7660 38892 8392 38944
rect 8444 38892 8460 38944
rect 8512 38892 8528 38944
rect 8580 38892 9312 38944
rect 9364 38892 9380 38944
rect 9432 38892 9448 38944
rect 9500 38892 10232 38944
rect 10284 38892 10300 38944
rect 10352 38892 10368 38944
rect 10420 38892 11152 38944
rect 11204 38892 11220 38944
rect 11272 38892 11288 38944
rect 11340 38892 12072 38944
rect 12124 38892 12140 38944
rect 12192 38892 12208 38944
rect 12260 38893 12992 38944
rect 13044 38893 13060 38945
rect 13112 38893 13128 38945
rect 13180 38893 13440 38945
rect 12260 38892 13440 38893
rect 7359 38881 13440 38892
rect 7359 38879 12992 38881
rect 7359 38869 7472 38879
rect 4900 38841 5632 38869
rect 5684 38841 5700 38869
rect 5752 38841 5768 38869
rect 5820 38841 6552 38869
rect 6604 38841 6620 38869
rect 6672 38841 6688 38869
rect 6740 38841 7472 38869
rect 4742 38814 4768 38827
rect 4824 38814 4850 38827
rect 4764 38785 4768 38814
rect 3912 38762 3928 38785
rect 3980 38762 4712 38785
rect 4764 38762 4780 38785
rect 4832 38762 4848 38814
rect 4906 38785 4932 38841
rect 4988 38785 5195 38841
rect 5251 38785 5276 38841
rect 5332 38785 5357 38841
rect 5413 38785 5438 38841
rect 5494 38785 5519 38841
rect 5575 38785 5600 38841
rect 5752 38827 5762 38841
rect 5820 38827 5843 38841
rect 5656 38814 5681 38827
rect 5737 38814 5762 38827
rect 5818 38814 5843 38827
rect 5752 38785 5762 38814
rect 5820 38785 5843 38814
rect 5899 38785 5924 38841
rect 5980 38785 6005 38841
rect 6061 38785 6086 38841
rect 6142 38785 6167 38841
rect 6223 38785 6248 38841
rect 6304 38785 6329 38841
rect 6385 38785 6410 38841
rect 6466 38785 6491 38841
rect 6547 38827 6552 38841
rect 6547 38814 6572 38827
rect 6628 38814 6653 38827
rect 6709 38814 6734 38827
rect 6547 38785 6552 38814
rect 6790 38785 6815 38841
rect 6871 38785 6896 38841
rect 6952 38785 6977 38841
rect 7033 38785 7058 38841
rect 7114 38785 7139 38841
rect 7195 38785 7221 38841
rect 7277 38785 7303 38841
rect 7359 38827 7472 38841
rect 7524 38827 7540 38879
rect 7592 38827 7608 38879
rect 7660 38827 8392 38879
rect 8444 38827 8460 38879
rect 8512 38827 8528 38879
rect 8580 38827 9312 38879
rect 9364 38827 9380 38879
rect 9432 38827 9448 38879
rect 9500 38827 10232 38879
rect 10284 38827 10300 38879
rect 10352 38827 10368 38879
rect 10420 38827 11152 38879
rect 11204 38827 11220 38879
rect 11272 38827 11288 38879
rect 11340 38827 12072 38879
rect 12124 38827 12140 38879
rect 12192 38827 12208 38879
rect 12260 38829 12992 38879
rect 13044 38829 13060 38881
rect 13112 38829 13128 38881
rect 13180 38829 13440 38881
rect 12260 38827 13440 38829
rect 7359 38817 13440 38827
rect 7359 38814 12992 38817
rect 7359 38785 7472 38814
rect 4900 38762 5632 38785
rect 5684 38762 5700 38785
rect 5752 38762 5768 38785
rect 5820 38762 6552 38785
rect 6604 38762 6620 38785
rect 6672 38762 6688 38785
rect 6740 38762 7472 38785
rect 7524 38762 7540 38814
rect 7592 38762 7608 38814
rect 7660 38762 8392 38814
rect 8444 38762 8460 38814
rect 8512 38762 8528 38814
rect 8580 38762 9312 38814
rect 9364 38762 9380 38814
rect 9432 38762 9448 38814
rect 9500 38762 10232 38814
rect 10284 38762 10300 38814
rect 10352 38762 10368 38814
rect 10420 38762 11152 38814
rect 11204 38762 11220 38814
rect 11272 38762 11288 38814
rect 11340 38762 12072 38814
rect 12124 38762 12140 38814
rect 12192 38762 12208 38814
rect 12260 38765 12992 38814
rect 13044 38765 13060 38817
rect 13112 38765 13128 38817
rect 13180 38765 13440 38817
rect 12260 38762 13440 38765
rect 187 38757 13440 38762
rect 187 38701 2534 38757
rect 2590 38701 2617 38757
rect 2673 38701 2700 38757
rect 2756 38701 2783 38757
rect 2839 38701 2866 38757
rect 2922 38749 2949 38757
rect 3005 38749 3032 38757
rect 187 38697 2872 38701
rect 2924 38697 2940 38749
rect 3005 38701 3008 38749
rect 3088 38701 3115 38757
rect 3171 38701 3198 38757
rect 3254 38701 3281 38757
rect 3337 38701 3364 38757
rect 3420 38701 3447 38757
rect 3503 38701 3530 38757
rect 3586 38701 3613 38757
rect 3669 38701 3696 38757
rect 3752 38701 3779 38757
rect 3835 38749 3862 38757
rect 3918 38749 3945 38757
rect 2992 38697 3008 38701
rect 3060 38697 3792 38701
rect 3844 38697 3860 38749
rect 3918 38701 3928 38749
rect 4001 38701 4028 38757
rect 4084 38701 4111 38757
rect 4167 38701 4194 38757
rect 4250 38701 4276 38757
rect 4332 38701 4358 38757
rect 4414 38701 4440 38757
rect 4496 38701 4522 38757
rect 4578 38701 4604 38757
rect 4660 38701 4686 38757
rect 4742 38749 4768 38757
rect 4824 38749 4850 38757
rect 4764 38701 4768 38749
rect 3912 38697 3928 38701
rect 3980 38697 4712 38701
rect 4764 38697 4780 38701
rect 4832 38697 4848 38749
rect 4906 38701 4932 38757
rect 4988 38701 5195 38757
rect 5251 38701 5276 38757
rect 5332 38701 5357 38757
rect 5413 38701 5438 38757
rect 5494 38701 5519 38757
rect 5575 38701 5600 38757
rect 5656 38749 5681 38757
rect 5737 38749 5762 38757
rect 5818 38749 5843 38757
rect 5752 38701 5762 38749
rect 5820 38701 5843 38749
rect 5899 38701 5924 38757
rect 5980 38701 6005 38757
rect 6061 38701 6086 38757
rect 6142 38701 6167 38757
rect 6223 38701 6248 38757
rect 6304 38701 6329 38757
rect 6385 38701 6410 38757
rect 6466 38701 6491 38757
rect 6547 38749 6572 38757
rect 6628 38749 6653 38757
rect 6709 38749 6734 38757
rect 6547 38701 6552 38749
rect 6790 38701 6815 38757
rect 6871 38701 6896 38757
rect 6952 38701 6977 38757
rect 7033 38701 7058 38757
rect 7114 38701 7139 38757
rect 7195 38701 7221 38757
rect 7277 38701 7303 38757
rect 7359 38753 13440 38757
rect 7359 38749 12992 38753
rect 7359 38701 7472 38749
rect 4900 38697 5632 38701
rect 5684 38697 5700 38701
rect 5752 38697 5768 38701
rect 5820 38697 6552 38701
rect 6604 38697 6620 38701
rect 6672 38697 6688 38701
rect 6740 38697 7472 38701
rect 7524 38697 7540 38749
rect 7592 38697 7608 38749
rect 7660 38697 8392 38749
rect 8444 38697 8460 38749
rect 8512 38697 8528 38749
rect 8580 38697 9312 38749
rect 9364 38697 9380 38749
rect 9432 38697 9448 38749
rect 9500 38697 10232 38749
rect 10284 38697 10300 38749
rect 10352 38697 10368 38749
rect 10420 38697 11152 38749
rect 11204 38697 11220 38749
rect 11272 38697 11288 38749
rect 11340 38697 12072 38749
rect 12124 38697 12140 38749
rect 12192 38697 12208 38749
rect 12260 38701 12992 38749
rect 13044 38701 13060 38753
rect 13112 38701 13128 38753
rect 13180 38701 13440 38753
rect 12260 38697 13440 38701
rect 187 38689 13440 38697
rect 187 38684 12992 38689
rect 187 38673 2872 38684
rect 187 38617 2534 38673
rect 2590 38617 2617 38673
rect 2673 38617 2700 38673
rect 2756 38617 2783 38673
rect 2839 38617 2866 38673
rect 2924 38632 2940 38684
rect 2992 38673 3008 38684
rect 3060 38673 3792 38684
rect 3005 38632 3008 38673
rect 2922 38619 2949 38632
rect 3005 38619 3032 38632
rect 187 38589 2872 38617
rect 187 38533 2534 38589
rect 2590 38533 2617 38589
rect 2673 38533 2700 38589
rect 2756 38533 2783 38589
rect 2839 38533 2866 38589
rect 2924 38567 2940 38619
rect 3005 38617 3008 38619
rect 3088 38617 3115 38673
rect 3171 38617 3198 38673
rect 3254 38617 3281 38673
rect 3337 38617 3364 38673
rect 3420 38617 3447 38673
rect 3503 38617 3530 38673
rect 3586 38617 3613 38673
rect 3669 38617 3696 38673
rect 3752 38617 3779 38673
rect 3844 38632 3860 38684
rect 3912 38673 3928 38684
rect 3980 38673 4712 38684
rect 4764 38673 4780 38684
rect 3918 38632 3928 38673
rect 3835 38619 3862 38632
rect 3918 38619 3945 38632
rect 2992 38589 3008 38617
rect 3060 38589 3792 38617
rect 3005 38567 3008 38589
rect 2922 38554 2949 38567
rect 3005 38554 3032 38567
rect 187 38505 2872 38533
rect 187 38449 2534 38505
rect 2590 38449 2617 38505
rect 2673 38449 2700 38505
rect 2756 38449 2783 38505
rect 2839 38449 2866 38505
rect 2924 38502 2940 38554
rect 3005 38533 3008 38554
rect 3088 38533 3115 38589
rect 3171 38533 3198 38589
rect 3254 38533 3281 38589
rect 3337 38533 3364 38589
rect 3420 38533 3447 38589
rect 3503 38533 3530 38589
rect 3586 38533 3613 38589
rect 3669 38533 3696 38589
rect 3752 38533 3779 38589
rect 3844 38567 3860 38619
rect 3918 38617 3928 38619
rect 4001 38617 4028 38673
rect 4084 38617 4111 38673
rect 4167 38617 4194 38673
rect 4250 38617 4276 38673
rect 4332 38617 4358 38673
rect 4414 38617 4440 38673
rect 4496 38617 4522 38673
rect 4578 38617 4604 38673
rect 4660 38617 4686 38673
rect 4764 38632 4768 38673
rect 4832 38632 4848 38684
rect 4900 38673 5632 38684
rect 5684 38673 5700 38684
rect 5752 38673 5768 38684
rect 5820 38673 6552 38684
rect 6604 38673 6620 38684
rect 6672 38673 6688 38684
rect 6740 38673 7472 38684
rect 4742 38619 4768 38632
rect 4824 38619 4850 38632
rect 4764 38617 4768 38619
rect 3912 38589 3928 38617
rect 3980 38589 4712 38617
rect 4764 38589 4780 38617
rect 3918 38567 3928 38589
rect 3835 38554 3862 38567
rect 3918 38554 3945 38567
rect 2992 38505 3008 38533
rect 3060 38505 3792 38533
rect 3005 38502 3008 38505
rect 2922 38490 2949 38502
rect 3005 38490 3032 38502
rect 187 38438 2872 38449
rect 2924 38438 2940 38490
rect 3005 38449 3008 38490
rect 3088 38449 3115 38505
rect 3171 38449 3198 38505
rect 3254 38449 3281 38505
rect 3337 38449 3364 38505
rect 3420 38449 3447 38505
rect 3503 38449 3530 38505
rect 3586 38449 3613 38505
rect 3669 38449 3696 38505
rect 3752 38449 3779 38505
rect 3844 38502 3860 38554
rect 3918 38533 3928 38554
rect 4001 38533 4028 38589
rect 4084 38533 4111 38589
rect 4167 38533 4194 38589
rect 4250 38533 4276 38589
rect 4332 38533 4358 38589
rect 4414 38533 4440 38589
rect 4496 38533 4522 38589
rect 4578 38533 4604 38589
rect 4660 38533 4686 38589
rect 4764 38567 4768 38589
rect 4832 38567 4848 38619
rect 4906 38617 4932 38673
rect 4988 38617 5195 38673
rect 5251 38617 5276 38673
rect 5332 38617 5357 38673
rect 5413 38617 5438 38673
rect 5494 38617 5519 38673
rect 5575 38617 5600 38673
rect 5752 38632 5762 38673
rect 5820 38632 5843 38673
rect 5656 38619 5681 38632
rect 5737 38619 5762 38632
rect 5818 38619 5843 38632
rect 5752 38617 5762 38619
rect 5820 38617 5843 38619
rect 5899 38617 5924 38673
rect 5980 38617 6005 38673
rect 6061 38617 6086 38673
rect 6142 38617 6167 38673
rect 6223 38617 6248 38673
rect 6304 38617 6329 38673
rect 6385 38617 6410 38673
rect 6466 38617 6491 38673
rect 6547 38632 6552 38673
rect 6547 38619 6572 38632
rect 6628 38619 6653 38632
rect 6709 38619 6734 38632
rect 6547 38617 6552 38619
rect 6790 38617 6815 38673
rect 6871 38617 6896 38673
rect 6952 38617 6977 38673
rect 7033 38617 7058 38673
rect 7114 38617 7139 38673
rect 7195 38617 7221 38673
rect 7277 38617 7303 38673
rect 7359 38632 7472 38673
rect 7524 38632 7540 38684
rect 7592 38632 7608 38684
rect 7660 38632 8392 38684
rect 8444 38632 8460 38684
rect 8512 38632 8528 38684
rect 8580 38632 9312 38684
rect 9364 38632 9380 38684
rect 9432 38632 9448 38684
rect 9500 38632 10232 38684
rect 10284 38632 10300 38684
rect 10352 38632 10368 38684
rect 10420 38632 11152 38684
rect 11204 38632 11220 38684
rect 11272 38632 11288 38684
rect 11340 38632 12072 38684
rect 12124 38632 12140 38684
rect 12192 38632 12208 38684
rect 12260 38637 12992 38684
rect 13044 38637 13060 38689
rect 13112 38637 13128 38689
rect 13180 38637 13440 38689
rect 12260 38632 13440 38637
rect 7359 38625 13440 38632
rect 7359 38619 12992 38625
rect 7359 38617 7472 38619
rect 4900 38589 5632 38617
rect 5684 38589 5700 38617
rect 5752 38589 5768 38617
rect 5820 38589 6552 38617
rect 6604 38589 6620 38617
rect 6672 38589 6688 38617
rect 6740 38589 7472 38617
rect 4742 38554 4768 38567
rect 4824 38554 4850 38567
rect 4764 38533 4768 38554
rect 3912 38505 3928 38533
rect 3980 38505 4712 38533
rect 4764 38505 4780 38533
rect 3918 38502 3928 38505
rect 3835 38490 3862 38502
rect 3918 38490 3945 38502
rect 2992 38438 3008 38449
rect 3060 38438 3792 38449
rect 3844 38438 3860 38490
rect 3918 38449 3928 38490
rect 4001 38449 4028 38505
rect 4084 38449 4111 38505
rect 4167 38449 4194 38505
rect 4250 38449 4276 38505
rect 4332 38449 4358 38505
rect 4414 38449 4440 38505
rect 4496 38449 4522 38505
rect 4578 38449 4604 38505
rect 4660 38449 4686 38505
rect 4764 38502 4768 38505
rect 4832 38502 4848 38554
rect 4906 38533 4932 38589
rect 4988 38533 5195 38589
rect 5251 38533 5276 38589
rect 5332 38533 5357 38589
rect 5413 38533 5438 38589
rect 5494 38533 5519 38589
rect 5575 38533 5600 38589
rect 5752 38567 5762 38589
rect 5820 38567 5843 38589
rect 5656 38554 5681 38567
rect 5737 38554 5762 38567
rect 5818 38554 5843 38567
rect 5752 38533 5762 38554
rect 5820 38533 5843 38554
rect 5899 38533 5924 38589
rect 5980 38533 6005 38589
rect 6061 38533 6086 38589
rect 6142 38533 6167 38589
rect 6223 38533 6248 38589
rect 6304 38533 6329 38589
rect 6385 38533 6410 38589
rect 6466 38533 6491 38589
rect 6547 38567 6552 38589
rect 6547 38554 6572 38567
rect 6628 38554 6653 38567
rect 6709 38554 6734 38567
rect 6547 38533 6552 38554
rect 6790 38533 6815 38589
rect 6871 38533 6896 38589
rect 6952 38533 6977 38589
rect 7033 38533 7058 38589
rect 7114 38533 7139 38589
rect 7195 38533 7221 38589
rect 7277 38533 7303 38589
rect 7359 38567 7472 38589
rect 7524 38567 7540 38619
rect 7592 38567 7608 38619
rect 7660 38567 8392 38619
rect 8444 38567 8460 38619
rect 8512 38567 8528 38619
rect 8580 38567 9312 38619
rect 9364 38567 9380 38619
rect 9432 38567 9448 38619
rect 9500 38567 10232 38619
rect 10284 38567 10300 38619
rect 10352 38567 10368 38619
rect 10420 38567 11152 38619
rect 11204 38567 11220 38619
rect 11272 38567 11288 38619
rect 11340 38567 12072 38619
rect 12124 38567 12140 38619
rect 12192 38567 12208 38619
rect 12260 38573 12992 38619
rect 13044 38573 13060 38625
rect 13112 38573 13128 38625
rect 13180 38573 13440 38625
rect 12260 38567 13440 38573
rect 7359 38560 13440 38567
rect 7359 38554 12992 38560
rect 7359 38533 7472 38554
rect 4900 38505 5632 38533
rect 5684 38505 5700 38533
rect 5752 38505 5768 38533
rect 5820 38505 6552 38533
rect 6604 38505 6620 38533
rect 6672 38505 6688 38533
rect 6740 38505 7472 38533
rect 4742 38490 4768 38502
rect 4824 38490 4850 38502
rect 4764 38449 4768 38490
rect 3912 38438 3928 38449
rect 3980 38438 4712 38449
rect 4764 38438 4780 38449
rect 4832 38438 4848 38490
rect 4906 38449 4932 38505
rect 4988 38449 5195 38505
rect 5251 38449 5276 38505
rect 5332 38449 5357 38505
rect 5413 38449 5438 38505
rect 5494 38449 5519 38505
rect 5575 38449 5600 38505
rect 5752 38502 5762 38505
rect 5820 38502 5843 38505
rect 5656 38490 5681 38502
rect 5737 38490 5762 38502
rect 5818 38490 5843 38502
rect 5752 38449 5762 38490
rect 5820 38449 5843 38490
rect 5899 38449 5924 38505
rect 5980 38449 6005 38505
rect 6061 38449 6086 38505
rect 6142 38449 6167 38505
rect 6223 38449 6248 38505
rect 6304 38449 6329 38505
rect 6385 38449 6410 38505
rect 6466 38449 6491 38505
rect 6547 38502 6552 38505
rect 6547 38490 6572 38502
rect 6628 38490 6653 38502
rect 6709 38490 6734 38502
rect 6547 38449 6552 38490
rect 6790 38449 6815 38505
rect 6871 38449 6896 38505
rect 6952 38449 6977 38505
rect 7033 38449 7058 38505
rect 7114 38449 7139 38505
rect 7195 38449 7221 38505
rect 7277 38449 7303 38505
rect 7359 38502 7472 38505
rect 7524 38502 7540 38554
rect 7592 38502 7608 38554
rect 7660 38502 8392 38554
rect 8444 38502 8460 38554
rect 8512 38502 8528 38554
rect 8580 38502 9312 38554
rect 9364 38502 9380 38554
rect 9432 38502 9448 38554
rect 9500 38502 10232 38554
rect 10284 38502 10300 38554
rect 10352 38502 10368 38554
rect 10420 38502 11152 38554
rect 11204 38502 11220 38554
rect 11272 38502 11288 38554
rect 11340 38502 12072 38554
rect 12124 38502 12140 38554
rect 12192 38502 12208 38554
rect 12260 38508 12992 38554
rect 13044 38508 13060 38560
rect 13112 38508 13128 38560
rect 13180 38508 13440 38560
rect 12260 38502 13440 38508
rect 7359 38495 13440 38502
rect 7359 38490 12992 38495
rect 7359 38449 7472 38490
rect 4900 38438 5632 38449
rect 5684 38438 5700 38449
rect 5752 38438 5768 38449
rect 5820 38438 6552 38449
rect 6604 38438 6620 38449
rect 6672 38438 6688 38449
rect 6740 38438 7472 38449
rect 7524 38438 7540 38490
rect 7592 38438 7608 38490
rect 7660 38438 8392 38490
rect 8444 38438 8460 38490
rect 8512 38438 8528 38490
rect 8580 38438 9312 38490
rect 9364 38438 9380 38490
rect 9432 38438 9448 38490
rect 9500 38438 10232 38490
rect 10284 38438 10300 38490
rect 10352 38438 10368 38490
rect 10420 38438 11152 38490
rect 11204 38438 11220 38490
rect 11272 38438 11288 38490
rect 11340 38438 12072 38490
rect 12124 38438 12140 38490
rect 12192 38438 12208 38490
rect 12260 38443 12992 38490
rect 13044 38443 13060 38495
rect 13112 38443 13128 38495
rect 13180 38443 13440 38495
rect 12260 38438 13440 38443
rect 187 38430 13440 38438
rect 187 38426 12992 38430
rect 187 38421 2872 38426
rect 187 38365 2534 38421
rect 2590 38365 2617 38421
rect 2673 38365 2700 38421
rect 2756 38365 2783 38421
rect 2839 38365 2866 38421
rect 2924 38374 2940 38426
rect 2992 38421 3008 38426
rect 3060 38421 3792 38426
rect 3005 38374 3008 38421
rect 2922 38365 2949 38374
rect 3005 38365 3032 38374
rect 3088 38365 3115 38421
rect 3171 38365 3198 38421
rect 3254 38365 3281 38421
rect 3337 38365 3364 38421
rect 3420 38365 3447 38421
rect 3503 38365 3530 38421
rect 3586 38365 3613 38421
rect 3669 38365 3696 38421
rect 3752 38365 3779 38421
rect 3844 38374 3860 38426
rect 3912 38421 3928 38426
rect 3980 38421 4712 38426
rect 4764 38421 4780 38426
rect 3918 38374 3928 38421
rect 3835 38365 3862 38374
rect 3918 38365 3945 38374
rect 4001 38365 4028 38421
rect 4084 38365 4111 38421
rect 4167 38365 4194 38421
rect 4250 38365 4276 38421
rect 4332 38365 4358 38421
rect 4414 38365 4440 38421
rect 4496 38365 4522 38421
rect 4578 38365 4604 38421
rect 4660 38365 4686 38421
rect 4764 38374 4768 38421
rect 4832 38374 4848 38426
rect 4900 38421 5632 38426
rect 5684 38421 5700 38426
rect 5752 38421 5768 38426
rect 5820 38421 6552 38426
rect 6604 38421 6620 38426
rect 6672 38421 6688 38426
rect 6740 38421 7472 38426
rect 4742 38365 4768 38374
rect 4824 38365 4850 38374
rect 4906 38365 4932 38421
rect 4988 38365 5195 38421
rect 5251 38365 5276 38421
rect 5332 38365 5357 38421
rect 5413 38365 5438 38421
rect 5494 38365 5519 38421
rect 5575 38365 5600 38421
rect 5752 38374 5762 38421
rect 5820 38374 5843 38421
rect 5656 38365 5681 38374
rect 5737 38365 5762 38374
rect 5818 38365 5843 38374
rect 5899 38365 5924 38421
rect 5980 38365 6005 38421
rect 6061 38365 6086 38421
rect 6142 38365 6167 38421
rect 6223 38365 6248 38421
rect 6304 38365 6329 38421
rect 6385 38365 6410 38421
rect 6466 38365 6491 38421
rect 6547 38374 6552 38421
rect 6547 38365 6572 38374
rect 6628 38365 6653 38374
rect 6709 38365 6734 38374
rect 6790 38365 6815 38421
rect 6871 38365 6896 38421
rect 6952 38365 6977 38421
rect 7033 38365 7058 38421
rect 7114 38365 7139 38421
rect 7195 38365 7221 38421
rect 7277 38365 7303 38421
rect 7359 38374 7472 38421
rect 7524 38374 7540 38426
rect 7592 38374 7608 38426
rect 7660 38374 8392 38426
rect 8444 38374 8460 38426
rect 8512 38374 8528 38426
rect 8580 38374 9312 38426
rect 9364 38374 9380 38426
rect 9432 38374 9448 38426
rect 9500 38374 10232 38426
rect 10284 38374 10300 38426
rect 10352 38374 10368 38426
rect 10420 38374 11152 38426
rect 11204 38374 11220 38426
rect 11272 38374 11288 38426
rect 11340 38374 12072 38426
rect 12124 38374 12140 38426
rect 12192 38374 12208 38426
rect 12260 38378 12992 38426
rect 13044 38378 13060 38430
rect 13112 38378 13128 38430
rect 13180 38378 13440 38430
rect 12260 38374 13440 38378
rect 7359 38365 13440 38374
rect 187 38362 12992 38365
rect 187 38337 2872 38362
rect 187 38281 2534 38337
rect 2590 38281 2617 38337
rect 2673 38281 2700 38337
rect 2756 38281 2783 38337
rect 2839 38281 2866 38337
rect 2924 38310 2940 38362
rect 2992 38337 3008 38362
rect 3060 38337 3792 38362
rect 3005 38310 3008 38337
rect 2922 38298 2949 38310
rect 3005 38298 3032 38310
rect 187 38253 2872 38281
rect 187 38197 2534 38253
rect 2590 38197 2617 38253
rect 2673 38197 2700 38253
rect 2756 38197 2783 38253
rect 2839 38197 2866 38253
rect 2924 38246 2940 38298
rect 3005 38281 3008 38298
rect 3088 38281 3115 38337
rect 3171 38281 3198 38337
rect 3254 38281 3281 38337
rect 3337 38281 3364 38337
rect 3420 38281 3447 38337
rect 3503 38281 3530 38337
rect 3586 38281 3613 38337
rect 3669 38281 3696 38337
rect 3752 38281 3779 38337
rect 3844 38310 3860 38362
rect 3912 38337 3928 38362
rect 3980 38337 4712 38362
rect 4764 38337 4780 38362
rect 3918 38310 3928 38337
rect 3835 38298 3862 38310
rect 3918 38298 3945 38310
rect 2992 38253 3008 38281
rect 3060 38253 3792 38281
rect 3005 38246 3008 38253
rect 2922 38234 2949 38246
rect 3005 38234 3032 38246
rect 187 38182 2872 38197
rect 2924 38182 2940 38234
rect 3005 38197 3008 38234
rect 3088 38197 3115 38253
rect 3171 38197 3198 38253
rect 3254 38197 3281 38253
rect 3337 38197 3364 38253
rect 3420 38197 3447 38253
rect 3503 38197 3530 38253
rect 3586 38197 3613 38253
rect 3669 38197 3696 38253
rect 3752 38197 3779 38253
rect 3844 38246 3860 38298
rect 3918 38281 3928 38298
rect 4001 38281 4028 38337
rect 4084 38281 4111 38337
rect 4167 38281 4194 38337
rect 4250 38281 4276 38337
rect 4332 38281 4358 38337
rect 4414 38281 4440 38337
rect 4496 38281 4522 38337
rect 4578 38281 4604 38337
rect 4660 38281 4686 38337
rect 4764 38310 4768 38337
rect 4832 38310 4848 38362
rect 4900 38337 5632 38362
rect 5684 38337 5700 38362
rect 5752 38337 5768 38362
rect 5820 38337 6552 38362
rect 6604 38337 6620 38362
rect 6672 38337 6688 38362
rect 6740 38337 7472 38362
rect 4742 38298 4768 38310
rect 4824 38298 4850 38310
rect 4764 38281 4768 38298
rect 3912 38253 3928 38281
rect 3980 38253 4712 38281
rect 4764 38253 4780 38281
rect 3918 38246 3928 38253
rect 3835 38234 3862 38246
rect 3918 38234 3945 38246
rect 2992 38182 3008 38197
rect 3060 38182 3792 38197
rect 3844 38182 3860 38234
rect 3918 38197 3928 38234
rect 4001 38197 4028 38253
rect 4084 38197 4111 38253
rect 4167 38197 4194 38253
rect 4250 38197 4276 38253
rect 4332 38197 4358 38253
rect 4414 38197 4440 38253
rect 4496 38197 4522 38253
rect 4578 38197 4604 38253
rect 4660 38197 4686 38253
rect 4764 38246 4768 38253
rect 4832 38246 4848 38298
rect 4906 38281 4932 38337
rect 4988 38281 5195 38337
rect 5251 38281 5276 38337
rect 5332 38281 5357 38337
rect 5413 38281 5438 38337
rect 5494 38281 5519 38337
rect 5575 38281 5600 38337
rect 5752 38310 5762 38337
rect 5820 38310 5843 38337
rect 5656 38298 5681 38310
rect 5737 38298 5762 38310
rect 5818 38298 5843 38310
rect 5752 38281 5762 38298
rect 5820 38281 5843 38298
rect 5899 38281 5924 38337
rect 5980 38281 6005 38337
rect 6061 38281 6086 38337
rect 6142 38281 6167 38337
rect 6223 38281 6248 38337
rect 6304 38281 6329 38337
rect 6385 38281 6410 38337
rect 6466 38281 6491 38337
rect 6547 38310 6552 38337
rect 6547 38298 6572 38310
rect 6628 38298 6653 38310
rect 6709 38298 6734 38310
rect 6547 38281 6552 38298
rect 6790 38281 6815 38337
rect 6871 38281 6896 38337
rect 6952 38281 6977 38337
rect 7033 38281 7058 38337
rect 7114 38281 7139 38337
rect 7195 38281 7221 38337
rect 7277 38281 7303 38337
rect 7359 38310 7472 38337
rect 7524 38310 7540 38362
rect 7592 38310 7608 38362
rect 7660 38310 8392 38362
rect 8444 38310 8460 38362
rect 8512 38310 8528 38362
rect 8580 38310 9312 38362
rect 9364 38310 9380 38362
rect 9432 38310 9448 38362
rect 9500 38310 10232 38362
rect 10284 38310 10300 38362
rect 10352 38310 10368 38362
rect 10420 38310 11152 38362
rect 11204 38310 11220 38362
rect 11272 38310 11288 38362
rect 11340 38310 12072 38362
rect 12124 38310 12140 38362
rect 12192 38310 12208 38362
rect 12260 38313 12992 38362
rect 13044 38313 13060 38365
rect 13112 38313 13128 38365
rect 13180 38313 13440 38365
rect 12260 38310 13440 38313
rect 7359 38300 13440 38310
rect 7359 38298 12992 38300
rect 7359 38281 7472 38298
rect 4900 38253 5632 38281
rect 5684 38253 5700 38281
rect 5752 38253 5768 38281
rect 5820 38253 6552 38281
rect 6604 38253 6620 38281
rect 6672 38253 6688 38281
rect 6740 38253 7472 38281
rect 4742 38234 4768 38246
rect 4824 38234 4850 38246
rect 4764 38197 4768 38234
rect 3912 38182 3928 38197
rect 3980 38182 4712 38197
rect 4764 38182 4780 38197
rect 4832 38182 4848 38234
rect 4906 38197 4932 38253
rect 4988 38197 5195 38253
rect 5251 38197 5276 38253
rect 5332 38197 5357 38253
rect 5413 38197 5438 38253
rect 5494 38197 5519 38253
rect 5575 38197 5600 38253
rect 5752 38246 5762 38253
rect 5820 38246 5843 38253
rect 5656 38234 5681 38246
rect 5737 38234 5762 38246
rect 5818 38234 5843 38246
rect 5752 38197 5762 38234
rect 5820 38197 5843 38234
rect 5899 38197 5924 38253
rect 5980 38197 6005 38253
rect 6061 38197 6086 38253
rect 6142 38197 6167 38253
rect 6223 38197 6248 38253
rect 6304 38197 6329 38253
rect 6385 38197 6410 38253
rect 6466 38197 6491 38253
rect 6547 38246 6552 38253
rect 6547 38234 6572 38246
rect 6628 38234 6653 38246
rect 6709 38234 6734 38246
rect 6547 38197 6552 38234
rect 6790 38197 6815 38253
rect 6871 38197 6896 38253
rect 6952 38197 6977 38253
rect 7033 38197 7058 38253
rect 7114 38197 7139 38253
rect 7195 38197 7221 38253
rect 7277 38197 7303 38253
rect 7359 38246 7472 38253
rect 7524 38246 7540 38298
rect 7592 38246 7608 38298
rect 7660 38246 8392 38298
rect 8444 38246 8460 38298
rect 8512 38246 8528 38298
rect 8580 38246 9312 38298
rect 9364 38246 9380 38298
rect 9432 38246 9448 38298
rect 9500 38246 10232 38298
rect 10284 38246 10300 38298
rect 10352 38246 10368 38298
rect 10420 38246 11152 38298
rect 11204 38246 11220 38298
rect 11272 38246 11288 38298
rect 11340 38246 12072 38298
rect 12124 38246 12140 38298
rect 12192 38246 12208 38298
rect 12260 38248 12992 38298
rect 13044 38248 13060 38300
rect 13112 38248 13128 38300
rect 13180 38248 13440 38300
rect 12260 38246 13440 38248
rect 7359 38235 13440 38246
rect 7359 38234 12992 38235
rect 7359 38197 7472 38234
rect 4900 38182 5632 38197
rect 5684 38182 5700 38197
rect 5752 38182 5768 38197
rect 5820 38182 6552 38197
rect 6604 38182 6620 38197
rect 6672 38182 6688 38197
rect 6740 38182 7472 38197
rect 7524 38182 7540 38234
rect 7592 38182 7608 38234
rect 7660 38182 8392 38234
rect 8444 38182 8460 38234
rect 8512 38182 8528 38234
rect 8580 38182 9312 38234
rect 9364 38182 9380 38234
rect 9432 38182 9448 38234
rect 9500 38182 10232 38234
rect 10284 38182 10300 38234
rect 10352 38182 10368 38234
rect 10420 38182 11152 38234
rect 11204 38182 11220 38234
rect 11272 38182 11288 38234
rect 11340 38182 12072 38234
rect 12124 38182 12140 38234
rect 12192 38182 12208 38234
rect 12260 38183 12992 38234
rect 13044 38183 13060 38235
rect 13112 38183 13128 38235
rect 13180 38183 13440 38235
rect 12260 38182 13440 38183
rect 187 38170 13440 38182
rect 187 38169 2872 38170
rect 187 38113 2534 38169
rect 2590 38113 2617 38169
rect 2673 38113 2700 38169
rect 2756 38113 2783 38169
rect 2839 38113 2866 38169
rect 2924 38118 2940 38170
rect 2992 38169 3008 38170
rect 3060 38169 3792 38170
rect 3005 38118 3008 38169
rect 2922 38113 2949 38118
rect 3005 38113 3032 38118
rect 3088 38113 3115 38169
rect 3171 38113 3198 38169
rect 3254 38113 3281 38169
rect 3337 38113 3364 38169
rect 3420 38113 3447 38169
rect 3503 38113 3530 38169
rect 3586 38113 3613 38169
rect 3669 38113 3696 38169
rect 3752 38113 3779 38169
rect 3844 38118 3860 38170
rect 3912 38169 3928 38170
rect 3980 38169 4712 38170
rect 4764 38169 4780 38170
rect 3918 38118 3928 38169
rect 3835 38113 3862 38118
rect 3918 38113 3945 38118
rect 4001 38113 4028 38169
rect 4084 38113 4111 38169
rect 4167 38113 4194 38169
rect 4250 38113 4276 38169
rect 4332 38113 4358 38169
rect 4414 38113 4440 38169
rect 4496 38113 4522 38169
rect 4578 38113 4604 38169
rect 4660 38113 4686 38169
rect 4764 38118 4768 38169
rect 4832 38118 4848 38170
rect 4900 38169 5632 38170
rect 5684 38169 5700 38170
rect 5752 38169 5768 38170
rect 5820 38169 6552 38170
rect 6604 38169 6620 38170
rect 6672 38169 6688 38170
rect 6740 38169 7472 38170
rect 4742 38113 4768 38118
rect 4824 38113 4850 38118
rect 4906 38113 4932 38169
rect 4988 38113 5195 38169
rect 5251 38113 5276 38169
rect 5332 38113 5357 38169
rect 5413 38113 5438 38169
rect 5494 38113 5519 38169
rect 5575 38113 5600 38169
rect 5752 38118 5762 38169
rect 5820 38118 5843 38169
rect 5656 38113 5681 38118
rect 5737 38113 5762 38118
rect 5818 38113 5843 38118
rect 5899 38113 5924 38169
rect 5980 38113 6005 38169
rect 6061 38113 6086 38169
rect 6142 38113 6167 38169
rect 6223 38113 6248 38169
rect 6304 38113 6329 38169
rect 6385 38113 6410 38169
rect 6466 38113 6491 38169
rect 6547 38118 6552 38169
rect 6547 38113 6572 38118
rect 6628 38113 6653 38118
rect 6709 38113 6734 38118
rect 6790 38113 6815 38169
rect 6871 38113 6896 38169
rect 6952 38113 6977 38169
rect 7033 38113 7058 38169
rect 7114 38113 7139 38169
rect 7195 38113 7221 38169
rect 7277 38113 7303 38169
rect 7359 38118 7472 38169
rect 7524 38118 7540 38170
rect 7592 38118 7608 38170
rect 7660 38118 8392 38170
rect 8444 38118 8460 38170
rect 8512 38118 8528 38170
rect 8580 38118 9312 38170
rect 9364 38118 9380 38170
rect 9432 38118 9448 38170
rect 9500 38118 10232 38170
rect 10284 38118 10300 38170
rect 10352 38118 10368 38170
rect 10420 38118 11152 38170
rect 11204 38118 11220 38170
rect 11272 38118 11288 38170
rect 11340 38118 12072 38170
rect 12124 38118 12140 38170
rect 12192 38118 12208 38170
rect 12260 38118 12992 38170
rect 13044 38118 13060 38170
rect 13112 38118 13128 38170
rect 13180 38118 13440 38170
rect 7359 38113 13440 38118
rect 187 38112 13440 38113
rect 187 38073 2824 38112
rect 187 38017 2531 38073
rect 2587 38017 2649 38073
rect 2705 38017 2767 38073
rect 2823 38017 2824 38073
rect 187 37993 2824 38017
rect 187 37941 2231 37993
rect 2283 37941 2335 37993
rect 2387 37988 2824 37993
rect 2387 37941 2531 37988
rect 187 37932 2531 37941
rect 2587 37932 2649 37988
rect 2705 37932 2767 37988
rect 2823 37932 2824 37988
rect 187 37929 2824 37932
rect 187 37877 2231 37929
rect 2283 37877 2335 37929
rect 2387 37903 2824 37929
tri 2824 37917 3019 38112 nw
rect 3124 37997 14858 38003
rect 3124 37945 3361 37997
rect 3413 37945 3439 37997
rect 3491 37945 4281 37997
rect 4333 37945 4359 37997
rect 4411 37945 5201 37997
rect 5253 37945 5279 37997
rect 5331 37945 6121 37997
rect 6173 37945 6199 37997
rect 6251 37945 7041 37997
rect 7093 37945 7119 37997
rect 7171 37945 7961 37997
rect 8013 37945 8039 37997
rect 8091 37945 8881 37997
rect 8933 37945 8959 37997
rect 9011 37945 9801 37997
rect 9853 37945 9879 37997
rect 9931 37945 10721 37997
rect 10773 37945 10799 37997
rect 10851 37945 11641 37997
rect 11693 37945 11719 37997
rect 11771 37945 12561 37997
rect 12613 37945 12639 37997
rect 12691 37945 14858 37997
rect 3124 37929 14858 37945
rect 2387 37877 2531 37903
rect 187 37865 2531 37877
rect 187 37813 2231 37865
rect 2283 37813 2335 37865
rect 2387 37847 2531 37865
rect 2587 37847 2649 37903
rect 2705 37847 2767 37903
rect 2823 37847 2824 37903
rect 2387 37818 2824 37847
rect 2387 37813 2531 37818
rect 187 37801 2531 37813
rect 187 37749 2231 37801
rect 2283 37749 2335 37801
rect 2387 37762 2531 37801
rect 2587 37762 2649 37818
rect 2705 37762 2767 37818
rect 2823 37762 2824 37818
rect 2387 37749 2824 37762
rect 187 37737 2824 37749
rect 187 37685 2231 37737
rect 2283 37685 2335 37737
rect 2387 37733 2824 37737
rect 2387 37685 2531 37733
rect 187 37677 2531 37685
rect 2587 37677 2649 37733
rect 2705 37677 2767 37733
rect 2823 37677 2824 37733
rect 187 37673 2824 37677
rect 187 37621 2231 37673
rect 2283 37621 2335 37673
rect 2387 37648 2824 37673
rect 2387 37621 2531 37648
rect 187 37609 2531 37621
rect 187 37557 2231 37609
rect 2283 37557 2335 37609
rect 2387 37592 2531 37609
rect 2587 37592 2649 37648
rect 2705 37592 2767 37648
rect 2823 37592 2824 37648
rect 2387 37563 2824 37592
rect 2387 37557 2531 37563
rect 187 37545 2531 37557
rect 187 37493 2231 37545
rect 2283 37493 2335 37545
rect 2387 37507 2531 37545
rect 2587 37507 2649 37563
rect 2705 37507 2767 37563
rect 2823 37507 2824 37563
rect 2387 37493 2824 37507
rect 187 37481 2824 37493
rect 187 37429 2231 37481
rect 2283 37429 2335 37481
rect 2387 37478 2824 37481
rect 2387 37429 2531 37478
rect 187 37422 2531 37429
rect 2587 37422 2649 37478
rect 2705 37422 2767 37478
rect 2823 37422 2824 37478
rect 187 37417 2824 37422
rect 187 37365 2231 37417
rect 2283 37365 2335 37417
rect 2387 37393 2824 37417
rect 2387 37365 2531 37393
rect 187 37353 2531 37365
rect 187 37301 2231 37353
rect 2283 37301 2335 37353
rect 2387 37337 2531 37353
rect 2587 37337 2649 37393
rect 2705 37337 2767 37393
rect 2823 37337 2824 37393
rect 2387 37308 2824 37337
rect 2387 37301 2531 37308
rect 187 37289 2531 37301
rect 187 37237 2231 37289
rect 2283 37237 2335 37289
rect 2387 37252 2531 37289
rect 2587 37252 2649 37308
rect 2705 37252 2767 37308
rect 2823 37252 2824 37308
rect 2387 37237 2824 37252
rect 187 37225 2824 37237
rect 187 37173 2231 37225
rect 2283 37173 2335 37225
rect 2387 37222 2824 37225
rect 2387 37173 2531 37222
rect 187 37166 2531 37173
rect 2587 37166 2649 37222
rect 2705 37166 2767 37222
rect 2823 37166 2824 37222
rect 187 37161 2824 37166
rect 187 37109 2231 37161
rect 2283 37109 2335 37161
rect 2387 37136 2824 37161
rect 2387 37109 2531 37136
rect 187 37097 2531 37109
rect 187 37045 2231 37097
rect 2283 37045 2335 37097
rect 2387 37080 2531 37097
rect 2587 37080 2649 37136
rect 2705 37080 2767 37136
rect 2823 37080 2824 37136
rect 2387 37050 2824 37080
rect 3124 37877 3361 37929
rect 3413 37877 3439 37929
rect 3491 37877 4281 37929
rect 4333 37877 4359 37929
rect 4411 37877 5201 37929
rect 5253 37877 5279 37929
rect 5331 37877 6121 37929
rect 6173 37877 6199 37929
rect 6251 37877 7041 37929
rect 7093 37877 7119 37929
rect 7171 37877 7961 37929
rect 8013 37877 8039 37929
rect 8091 37877 8881 37929
rect 8933 37877 8959 37929
rect 9011 37877 9801 37929
rect 9853 37877 9879 37929
rect 9931 37877 10721 37929
rect 10773 37877 10799 37929
rect 10851 37877 11641 37929
rect 11693 37877 11719 37929
rect 11771 37877 12561 37929
rect 12613 37877 12639 37929
rect 12691 37877 14858 37929
rect 3124 37861 14858 37877
rect 3124 37809 3361 37861
rect 3413 37809 3439 37861
rect 3491 37809 4281 37861
rect 4333 37809 4359 37861
rect 4411 37809 5201 37861
rect 5253 37809 5279 37861
rect 5331 37809 6121 37861
rect 6173 37809 6199 37861
rect 6251 37809 7041 37861
rect 7093 37809 7119 37861
rect 7171 37809 7961 37861
rect 8013 37809 8039 37861
rect 8091 37809 8881 37861
rect 8933 37809 8959 37861
rect 9011 37809 9801 37861
rect 9853 37809 9879 37861
rect 9931 37809 10721 37861
rect 10773 37809 10799 37861
rect 10851 37809 11641 37861
rect 11693 37809 11719 37861
rect 11771 37809 12561 37861
rect 12613 37809 12639 37861
rect 12691 37809 14858 37861
rect 3124 37793 14858 37809
rect 3124 37741 3361 37793
rect 3413 37741 3439 37793
rect 3491 37741 4281 37793
rect 4333 37741 4359 37793
rect 4411 37741 5201 37793
rect 5253 37741 5279 37793
rect 5331 37741 6121 37793
rect 6173 37741 6199 37793
rect 6251 37741 7041 37793
rect 7093 37741 7119 37793
rect 7171 37741 7961 37793
rect 8013 37741 8039 37793
rect 8091 37741 8881 37793
rect 8933 37741 8959 37793
rect 9011 37741 9801 37793
rect 9853 37741 9879 37793
rect 9931 37741 10721 37793
rect 10773 37741 10799 37793
rect 10851 37741 11641 37793
rect 11693 37741 11719 37793
rect 11771 37741 12561 37793
rect 12613 37741 12639 37793
rect 12691 37741 14858 37793
rect 3124 37725 14858 37741
rect 3124 37673 3361 37725
rect 3413 37673 3439 37725
rect 3491 37673 4281 37725
rect 4333 37673 4359 37725
rect 4411 37673 5201 37725
rect 5253 37673 5279 37725
rect 5331 37673 6121 37725
rect 6173 37673 6199 37725
rect 6251 37673 7041 37725
rect 7093 37673 7119 37725
rect 7171 37673 7961 37725
rect 8013 37673 8039 37725
rect 8091 37673 8881 37725
rect 8933 37673 8959 37725
rect 9011 37673 9801 37725
rect 9853 37673 9879 37725
rect 9931 37673 10721 37725
rect 10773 37673 10799 37725
rect 10851 37673 11641 37725
rect 11693 37673 11719 37725
rect 11771 37673 12561 37725
rect 12613 37673 12639 37725
rect 12691 37673 14858 37725
rect 3124 37657 14858 37673
rect 3124 37605 3361 37657
rect 3413 37605 3439 37657
rect 3491 37605 4281 37657
rect 4333 37605 4359 37657
rect 4411 37605 5201 37657
rect 5253 37605 5279 37657
rect 5331 37605 6121 37657
rect 6173 37605 6199 37657
rect 6251 37605 7041 37657
rect 7093 37605 7119 37657
rect 7171 37605 7961 37657
rect 8013 37605 8039 37657
rect 8091 37605 8881 37657
rect 8933 37605 8959 37657
rect 9011 37605 9801 37657
rect 9853 37605 9879 37657
rect 9931 37605 10721 37657
rect 10773 37605 10799 37657
rect 10851 37605 11641 37657
rect 11693 37605 11719 37657
rect 11771 37605 12561 37657
rect 12613 37605 12639 37657
rect 12691 37605 14858 37657
rect 3124 37589 14858 37605
rect 3124 37537 3361 37589
rect 3413 37537 3439 37589
rect 3491 37537 4281 37589
rect 4333 37537 4359 37589
rect 4411 37537 5201 37589
rect 5253 37537 5279 37589
rect 5331 37537 6121 37589
rect 6173 37537 6199 37589
rect 6251 37537 7041 37589
rect 7093 37537 7119 37589
rect 7171 37537 7961 37589
rect 8013 37537 8039 37589
rect 8091 37537 8881 37589
rect 8933 37537 8959 37589
rect 9011 37537 9801 37589
rect 9853 37537 9879 37589
rect 9931 37537 10721 37589
rect 10773 37537 10799 37589
rect 10851 37537 11641 37589
rect 11693 37537 11719 37589
rect 11771 37537 12561 37589
rect 12613 37537 12639 37589
rect 12691 37537 14858 37589
rect 3124 37521 14858 37537
rect 3124 37469 3361 37521
rect 3413 37469 3439 37521
rect 3491 37469 4281 37521
rect 4333 37469 4359 37521
rect 4411 37469 5201 37521
rect 5253 37469 5279 37521
rect 5331 37469 6121 37521
rect 6173 37469 6199 37521
rect 6251 37469 7041 37521
rect 7093 37469 7119 37521
rect 7171 37469 7961 37521
rect 8013 37469 8039 37521
rect 8091 37469 8881 37521
rect 8933 37469 8959 37521
rect 9011 37469 9801 37521
rect 9853 37469 9879 37521
rect 9931 37469 10721 37521
rect 10773 37469 10799 37521
rect 10851 37469 11641 37521
rect 11693 37469 11719 37521
rect 11771 37469 12561 37521
rect 12613 37469 12639 37521
rect 12691 37469 14858 37521
rect 3124 37453 14858 37469
rect 3124 37401 3361 37453
rect 3413 37401 3439 37453
rect 3491 37401 4281 37453
rect 4333 37401 4359 37453
rect 4411 37401 5201 37453
rect 5253 37401 5279 37453
rect 5331 37401 6121 37453
rect 6173 37401 6199 37453
rect 6251 37401 7041 37453
rect 7093 37401 7119 37453
rect 7171 37401 7961 37453
rect 8013 37401 8039 37453
rect 8091 37401 8881 37453
rect 8933 37401 8959 37453
rect 9011 37401 9801 37453
rect 9853 37401 9879 37453
rect 9931 37401 10721 37453
rect 10773 37401 10799 37453
rect 10851 37401 11641 37453
rect 11693 37401 11719 37453
rect 11771 37401 12561 37453
rect 12613 37401 12639 37453
rect 12691 37401 14858 37453
rect 3124 37385 14858 37401
rect 3124 37333 3361 37385
rect 3413 37333 3439 37385
rect 3491 37333 4281 37385
rect 4333 37333 4359 37385
rect 4411 37333 5201 37385
rect 5253 37333 5279 37385
rect 5331 37333 6121 37385
rect 6173 37333 6199 37385
rect 6251 37333 7041 37385
rect 7093 37333 7119 37385
rect 7171 37333 7961 37385
rect 8013 37333 8039 37385
rect 8091 37333 8881 37385
rect 8933 37333 8959 37385
rect 9011 37333 9801 37385
rect 9853 37333 9879 37385
rect 9931 37333 10721 37385
rect 10773 37333 10799 37385
rect 10851 37333 11641 37385
rect 11693 37333 11719 37385
rect 11771 37333 12561 37385
rect 12613 37333 12639 37385
rect 12691 37333 14858 37385
rect 3124 37318 14858 37333
rect 3124 37266 3361 37318
rect 3413 37266 3439 37318
rect 3491 37266 4281 37318
rect 4333 37266 4359 37318
rect 4411 37266 5201 37318
rect 5253 37266 5279 37318
rect 5331 37266 6121 37318
rect 6173 37266 6199 37318
rect 6251 37266 7041 37318
rect 7093 37266 7119 37318
rect 7171 37266 7961 37318
rect 8013 37266 8039 37318
rect 8091 37266 8881 37318
rect 8933 37266 8959 37318
rect 9011 37266 9801 37318
rect 9853 37266 9879 37318
rect 9931 37266 10721 37318
rect 10773 37266 10799 37318
rect 10851 37266 11641 37318
rect 11693 37266 11719 37318
rect 11771 37266 12561 37318
rect 12613 37266 12639 37318
rect 12691 37266 14858 37318
rect 3124 37251 14858 37266
rect 3124 37199 3361 37251
rect 3413 37199 3439 37251
rect 3491 37199 4281 37251
rect 4333 37199 4359 37251
rect 4411 37199 5201 37251
rect 5253 37199 5279 37251
rect 5331 37199 6121 37251
rect 6173 37199 6199 37251
rect 6251 37199 7041 37251
rect 7093 37199 7119 37251
rect 7171 37199 7961 37251
rect 8013 37199 8039 37251
rect 8091 37199 8881 37251
rect 8933 37199 8959 37251
rect 9011 37199 9801 37251
rect 9853 37199 9879 37251
rect 9931 37199 10721 37251
rect 10773 37199 10799 37251
rect 10851 37199 11641 37251
rect 11693 37199 11719 37251
rect 11771 37199 12561 37251
rect 12613 37199 12639 37251
rect 12691 37199 14858 37251
rect 3124 37184 14858 37199
rect 3124 37132 3361 37184
rect 3413 37132 3439 37184
rect 3491 37132 4281 37184
rect 4333 37132 4359 37184
rect 4411 37132 5201 37184
rect 5253 37132 5279 37184
rect 5331 37132 6121 37184
rect 6173 37132 6199 37184
rect 6251 37132 7041 37184
rect 7093 37132 7119 37184
rect 7171 37132 7961 37184
rect 8013 37132 8039 37184
rect 8091 37132 8881 37184
rect 8933 37132 8959 37184
rect 9011 37132 9801 37184
rect 9853 37132 9879 37184
rect 9931 37132 10721 37184
rect 10773 37132 10799 37184
rect 10851 37132 11641 37184
rect 11693 37132 11719 37184
rect 11771 37132 12561 37184
rect 12613 37132 12639 37184
rect 12691 37132 14858 37184
rect 3124 37117 14858 37132
rect 3124 37065 3361 37117
rect 3413 37065 3439 37117
rect 3491 37065 4281 37117
rect 4333 37065 4359 37117
rect 4411 37065 5201 37117
rect 5253 37065 5279 37117
rect 5331 37065 6121 37117
rect 6173 37065 6199 37117
rect 6251 37065 7041 37117
rect 7093 37065 7119 37117
rect 7171 37065 7961 37117
rect 8013 37065 8039 37117
rect 8091 37065 8881 37117
rect 8933 37065 8959 37117
rect 9011 37065 9801 37117
rect 9853 37065 9879 37117
rect 9931 37065 10721 37117
rect 10773 37065 10799 37117
rect 10851 37065 11641 37117
rect 11693 37065 11719 37117
rect 11771 37065 12561 37117
rect 12613 37065 12639 37117
rect 12691 37065 14858 37117
rect 3124 37059 14858 37065
rect 2387 37045 2531 37050
rect 187 37033 2531 37045
rect 187 36981 2231 37033
rect 2283 36981 2335 37033
rect 2387 36994 2531 37033
rect 2587 36994 2649 37050
rect 2705 36994 2767 37050
rect 2823 36994 2824 37050
rect 2387 36981 2824 36994
rect 187 36969 2824 36981
rect 187 36917 2231 36969
rect 2283 36917 2335 36969
rect 2387 36964 2824 36969
rect 2387 36917 2531 36964
rect 187 36908 2531 36917
rect 2587 36908 2649 36964
rect 2705 36908 2767 36964
rect 2823 36908 2824 36964
rect 187 36905 2824 36908
rect 187 36853 2231 36905
rect 2283 36853 2335 36905
rect 2387 36878 2824 36905
rect 2387 36853 2531 36878
rect 187 36841 2531 36853
rect 187 36789 2231 36841
rect 2283 36789 2335 36841
rect 2387 36822 2531 36841
rect 2587 36822 2649 36878
rect 2705 36822 2767 36878
rect 2823 36822 2824 36878
rect 2387 36789 2824 36822
rect 187 36781 2824 36789
tri 2824 36781 3054 37011 sw
rect 187 36777 3064 36781
rect 187 36725 2231 36777
rect 2283 36725 2335 36777
rect 2387 36772 3064 36777
rect 2387 36725 2538 36772
rect 187 36716 2538 36725
rect 2594 36716 2632 36772
rect 2688 36716 2726 36772
rect 2782 36716 2820 36772
rect 2876 36716 2914 36772
rect 2970 36716 3008 36772
rect 187 36713 3064 36716
rect 187 36661 2231 36713
rect 2283 36661 2335 36713
rect 2387 36692 3064 36713
rect 2387 36661 2538 36692
rect 187 36649 2538 36661
rect 187 36597 2231 36649
rect 2283 36597 2335 36649
rect 2387 36636 2538 36649
rect 2594 36636 2632 36692
rect 2688 36636 2726 36692
rect 2782 36636 2820 36692
rect 2876 36636 2914 36692
rect 2970 36636 3008 36692
tri 3064 36673 3162 36771 sw
rect 3064 36650 3162 36673
rect 3064 36636 3099 36650
rect 2387 36612 3099 36636
rect 2387 36597 2538 36612
rect 187 36585 2538 36597
rect 187 36533 2231 36585
rect 2283 36533 2335 36585
rect 2387 36556 2538 36585
rect 2594 36556 2632 36612
rect 2688 36556 2726 36612
rect 2782 36556 2820 36612
rect 2876 36556 2914 36612
rect 2970 36556 3008 36612
rect 3064 36594 3099 36612
rect 3155 36594 3162 36650
rect 3064 36571 3162 36594
tri 3162 36571 3264 36673 sw
tri 11739 36576 12222 37059 ne
rect 3064 36562 3264 36571
rect 3064 36556 3112 36562
rect 2387 36533 3112 36556
rect 187 36532 3112 36533
rect 187 36521 2538 36532
rect 187 36469 2231 36521
rect 2283 36469 2335 36521
rect 2387 36476 2538 36521
rect 2594 36476 2632 36532
rect 2688 36476 2726 36532
rect 2782 36476 2820 36532
rect 2876 36476 2914 36532
rect 2970 36476 3008 36532
rect 3064 36506 3112 36532
rect 3168 36506 3206 36562
rect 3262 36506 3264 36562
rect 3064 36476 3264 36506
rect 2387 36469 3112 36476
rect 187 36457 3112 36469
rect 187 36405 2231 36457
rect 2283 36405 2335 36457
rect 2387 36452 3112 36457
rect 2387 36405 2538 36452
rect 187 36396 2538 36405
rect 2594 36396 2632 36452
rect 2688 36396 2726 36452
rect 2782 36396 2820 36452
rect 2876 36396 2914 36452
rect 2970 36396 3008 36452
rect 3064 36420 3112 36452
rect 3168 36420 3206 36476
rect 3262 36445 3264 36476
tri 3264 36445 3390 36571 sw
rect 3262 36420 3390 36445
rect 3064 36415 3390 36420
rect 3064 36396 3321 36415
rect 187 36393 3321 36396
rect 187 36341 2231 36393
rect 2283 36341 2335 36393
rect 2387 36390 3321 36393
rect 2387 36372 3112 36390
rect 2387 36341 2538 36372
rect 187 36329 2538 36341
rect 187 36277 2231 36329
rect 2283 36277 2335 36329
rect 2387 36316 2538 36329
rect 2594 36316 2632 36372
rect 2688 36316 2726 36372
rect 2782 36316 2820 36372
rect 2876 36368 2914 36372
rect 2970 36368 3008 36372
rect 2992 36316 3008 36368
rect 3064 36334 3112 36372
rect 3168 36334 3206 36390
rect 3262 36359 3321 36390
rect 3377 36359 3390 36415
rect 3262 36334 3390 36359
rect 3064 36316 3390 36334
rect 2387 36304 3390 36316
rect 2387 36292 2872 36304
rect 2924 36292 2940 36304
rect 2387 36277 2538 36292
rect 187 36265 2538 36277
rect 187 36213 2231 36265
rect 2283 36213 2335 36265
rect 2387 36236 2538 36265
rect 2594 36236 2632 36292
rect 2688 36236 2726 36292
rect 2782 36236 2820 36292
rect 2992 36252 3008 36304
rect 3060 36296 3390 36304
tri 3390 36296 3539 36445 sw
rect 3060 36294 11592 36296
rect 3060 36292 3109 36294
rect 2876 36239 2914 36252
rect 2970 36239 3008 36252
rect 2387 36213 2872 36236
rect 187 36212 2872 36213
rect 2924 36212 2940 36236
rect 187 36201 2538 36212
rect 187 36149 2231 36201
rect 2283 36149 2335 36201
rect 2387 36156 2538 36201
rect 2594 36156 2632 36212
rect 2688 36156 2726 36212
rect 2782 36156 2820 36212
rect 2992 36187 3008 36239
rect 3064 36238 3109 36292
rect 3165 36238 3193 36294
rect 3249 36238 3277 36294
rect 3333 36238 3360 36294
rect 3416 36238 3443 36294
rect 3499 36238 3526 36294
rect 3582 36238 3609 36294
rect 3665 36238 3692 36294
rect 3748 36238 3775 36294
rect 3831 36290 3858 36294
rect 3914 36290 3941 36294
rect 3844 36238 3858 36290
rect 3914 36238 3928 36290
rect 3997 36238 4024 36294
rect 4080 36238 4107 36294
rect 4163 36238 4190 36294
rect 4246 36238 4273 36294
rect 4329 36238 4356 36294
rect 4412 36238 4439 36294
rect 4495 36238 4522 36294
rect 4578 36238 4605 36294
rect 4661 36238 4688 36294
rect 4744 36290 4771 36294
rect 4827 36290 4854 36294
rect 4764 36238 4771 36290
rect 4832 36238 4848 36290
rect 4910 36238 4937 36294
rect 4993 36238 5195 36294
rect 5251 36238 5277 36294
rect 5333 36238 5359 36294
rect 5415 36238 5441 36294
rect 5497 36238 5523 36294
rect 5579 36238 5605 36294
rect 5661 36290 5687 36294
rect 5743 36290 5769 36294
rect 5684 36238 5687 36290
rect 5752 36238 5768 36290
rect 5825 36238 5851 36294
rect 5907 36238 5933 36294
rect 5989 36238 6015 36294
rect 6071 36238 6097 36294
rect 6153 36238 6179 36294
rect 6235 36238 6261 36294
rect 6317 36238 6343 36294
rect 6399 36238 6425 36294
rect 6481 36238 6507 36294
rect 6563 36290 6589 36294
rect 6645 36290 6671 36294
rect 6727 36290 6753 36294
rect 6740 36238 6753 36290
rect 6809 36290 11592 36294
rect 6809 36278 7472 36290
rect 6809 36238 6853 36278
rect 3064 36236 6853 36238
rect 3060 36226 6853 36236
rect 3060 36214 3792 36226
rect 3844 36214 3860 36226
rect 3912 36214 3928 36226
rect 3980 36214 4712 36226
rect 4764 36214 4780 36226
rect 3060 36212 3109 36214
rect 2876 36174 2914 36187
rect 2970 36174 3008 36187
rect 2387 36149 2872 36156
rect 187 36137 2872 36149
rect 187 36085 2231 36137
rect 2283 36085 2335 36137
rect 2387 36132 2872 36137
rect 2924 36132 2940 36156
rect 2387 36085 2538 36132
rect 187 36076 2538 36085
rect 2594 36076 2632 36132
rect 2688 36076 2726 36132
rect 2782 36076 2820 36132
rect 2992 36122 3008 36174
rect 3064 36158 3109 36212
rect 3165 36158 3193 36214
rect 3249 36158 3277 36214
rect 3333 36158 3360 36214
rect 3416 36158 3443 36214
rect 3499 36158 3526 36214
rect 3582 36158 3609 36214
rect 3665 36158 3692 36214
rect 3748 36158 3775 36214
rect 3844 36174 3858 36214
rect 3914 36174 3928 36214
rect 3831 36162 3858 36174
rect 3914 36162 3941 36174
rect 3844 36158 3858 36162
rect 3914 36158 3928 36162
rect 3997 36158 4024 36214
rect 4080 36158 4107 36214
rect 4163 36158 4190 36214
rect 4246 36158 4273 36214
rect 4329 36158 4356 36214
rect 4412 36158 4439 36214
rect 4495 36158 4522 36214
rect 4578 36158 4605 36214
rect 4661 36158 4688 36214
rect 4764 36174 4771 36214
rect 4832 36174 4848 36226
rect 4900 36214 5632 36226
rect 5684 36214 5700 36226
rect 4744 36162 4771 36174
rect 4827 36162 4854 36174
rect 4764 36158 4771 36162
rect 3064 36156 3792 36158
rect 3060 36134 3792 36156
rect 3844 36134 3860 36158
rect 3912 36134 3928 36158
rect 3980 36134 4712 36158
rect 4764 36134 4780 36158
rect 3060 36132 3109 36134
rect 2876 36109 2914 36122
rect 2970 36109 3008 36122
rect 187 36073 2872 36076
rect 187 36021 2231 36073
rect 2283 36021 2335 36073
rect 2387 36057 2872 36073
rect 2924 36057 2940 36076
rect 2992 36057 3008 36109
rect 3064 36078 3109 36132
rect 3165 36078 3193 36134
rect 3249 36078 3277 36134
rect 3333 36078 3360 36134
rect 3416 36078 3443 36134
rect 3499 36078 3526 36134
rect 3582 36078 3609 36134
rect 3665 36078 3692 36134
rect 3748 36078 3775 36134
rect 3844 36110 3858 36134
rect 3914 36110 3928 36134
rect 3831 36098 3858 36110
rect 3914 36098 3941 36110
rect 3844 36078 3858 36098
rect 3914 36078 3928 36098
rect 3997 36078 4024 36134
rect 4080 36078 4107 36134
rect 4163 36078 4190 36134
rect 4246 36078 4273 36134
rect 4329 36078 4356 36134
rect 4412 36078 4439 36134
rect 4495 36078 4522 36134
rect 4578 36078 4605 36134
rect 4661 36078 4688 36134
rect 4764 36110 4771 36134
rect 4832 36110 4848 36162
rect 4910 36158 4937 36214
rect 4993 36158 5195 36214
rect 5251 36158 5277 36214
rect 5333 36158 5359 36214
rect 5415 36158 5441 36214
rect 5497 36158 5523 36214
rect 5579 36158 5605 36214
rect 5684 36174 5687 36214
rect 5752 36174 5768 36226
rect 5820 36214 6552 36226
rect 6604 36214 6620 36226
rect 6672 36214 6688 36226
rect 6740 36222 6853 36226
rect 6909 36222 6941 36278
rect 6997 36222 7029 36278
rect 7085 36222 7117 36278
rect 7173 36222 7205 36278
rect 7261 36222 7293 36278
rect 7349 36238 7472 36278
rect 7524 36238 7540 36290
rect 7592 36238 7608 36290
rect 7660 36238 8392 36290
rect 8444 36238 8460 36290
rect 8512 36238 8528 36290
rect 8580 36238 9312 36290
rect 9364 36238 9380 36290
rect 9432 36238 9448 36290
rect 9500 36238 10232 36290
rect 10284 36238 10300 36290
rect 10352 36238 10368 36290
rect 10420 36238 11152 36290
rect 11204 36238 11220 36290
rect 11272 36238 11288 36290
rect 11340 36238 11592 36290
rect 7349 36226 11592 36238
rect 7349 36222 7472 36226
rect 6740 36214 7472 36222
rect 5661 36162 5687 36174
rect 5743 36162 5769 36174
rect 5684 36158 5687 36162
rect 4900 36134 5632 36158
rect 5684 36134 5700 36158
rect 4744 36098 4771 36110
rect 4827 36098 4854 36110
rect 4764 36078 4771 36098
rect 3064 36076 3792 36078
rect 3060 36057 3792 36076
rect 2387 36054 3792 36057
rect 3844 36054 3860 36078
rect 3912 36054 3928 36078
rect 3980 36054 4712 36078
rect 4764 36054 4780 36078
rect 2387 36052 3109 36054
rect 2387 36021 2538 36052
rect 187 36009 2538 36021
rect 187 35957 2231 36009
rect 2283 35957 2335 36009
rect 2387 35996 2538 36009
rect 2594 35996 2632 36052
rect 2688 35996 2726 36052
rect 2782 35996 2820 36052
rect 2876 36044 2914 36052
rect 2970 36044 3008 36052
rect 2387 35992 2872 35996
rect 2924 35992 2940 35996
rect 2992 35992 3008 36044
rect 3064 35998 3109 36052
rect 3165 35998 3193 36054
rect 3249 35998 3277 36054
rect 3333 35998 3360 36054
rect 3416 35998 3443 36054
rect 3499 35998 3526 36054
rect 3582 35998 3609 36054
rect 3665 35998 3692 36054
rect 3748 35998 3775 36054
rect 3844 36046 3858 36054
rect 3914 36046 3928 36054
rect 3831 36034 3858 36046
rect 3914 36034 3941 36046
rect 3844 35998 3858 36034
rect 3914 35998 3928 36034
rect 3997 35998 4024 36054
rect 4080 35998 4107 36054
rect 4163 35998 4190 36054
rect 4246 35998 4273 36054
rect 4329 35998 4356 36054
rect 4412 35998 4439 36054
rect 4495 35998 4522 36054
rect 4578 35998 4605 36054
rect 4661 35998 4688 36054
rect 4764 36046 4771 36054
rect 4832 36046 4848 36098
rect 4910 36078 4937 36134
rect 4993 36078 5195 36134
rect 5251 36078 5277 36134
rect 5333 36078 5359 36134
rect 5415 36078 5441 36134
rect 5497 36078 5523 36134
rect 5579 36078 5605 36134
rect 5684 36110 5687 36134
rect 5752 36110 5768 36162
rect 5825 36158 5851 36214
rect 5907 36158 5933 36214
rect 5989 36158 6015 36214
rect 6071 36158 6097 36214
rect 6153 36158 6179 36214
rect 6235 36158 6261 36214
rect 6317 36158 6343 36214
rect 6399 36158 6425 36214
rect 6481 36158 6507 36214
rect 6740 36174 6753 36214
rect 6563 36162 6589 36174
rect 6645 36162 6671 36174
rect 6727 36162 6753 36174
rect 6740 36158 6753 36162
rect 6809 36196 7472 36214
rect 6809 36158 6853 36196
rect 5820 36134 6552 36158
rect 6604 36134 6620 36158
rect 6672 36134 6688 36158
rect 6740 36140 6853 36158
rect 6909 36140 6941 36196
rect 6997 36140 7029 36196
rect 7085 36140 7117 36196
rect 7173 36140 7205 36196
rect 7261 36140 7293 36196
rect 7349 36174 7472 36196
rect 7524 36174 7540 36226
rect 7592 36174 7608 36226
rect 7660 36174 8392 36226
rect 8444 36174 8460 36226
rect 8512 36174 8528 36226
rect 8580 36174 9312 36226
rect 9364 36174 9380 36226
rect 9432 36174 9448 36226
rect 9500 36174 10232 36226
rect 10284 36174 10300 36226
rect 10352 36174 10368 36226
rect 10420 36174 11152 36226
rect 11204 36174 11220 36226
rect 11272 36174 11288 36226
rect 11340 36174 11592 36226
rect 7349 36162 11592 36174
rect 7349 36140 7472 36162
rect 6740 36134 7472 36140
rect 5661 36098 5687 36110
rect 5743 36098 5769 36110
rect 5684 36078 5687 36098
rect 4900 36054 5632 36078
rect 5684 36054 5700 36078
rect 4744 36034 4771 36046
rect 4827 36034 4854 36046
rect 4764 35998 4771 36034
rect 3064 35996 3792 35998
rect 3060 35992 3792 35996
rect 2387 35982 3792 35992
rect 3844 35982 3860 35998
rect 3912 35982 3928 35998
rect 3980 35982 4712 35998
rect 4764 35982 4780 35998
rect 4832 35982 4848 36034
rect 4910 35998 4937 36054
rect 4993 35998 5195 36054
rect 5251 35998 5277 36054
rect 5333 35998 5359 36054
rect 5415 35998 5441 36054
rect 5497 35998 5523 36054
rect 5579 35998 5605 36054
rect 5684 36046 5687 36054
rect 5752 36046 5768 36098
rect 5825 36078 5851 36134
rect 5907 36078 5933 36134
rect 5989 36078 6015 36134
rect 6071 36078 6097 36134
rect 6153 36078 6179 36134
rect 6235 36078 6261 36134
rect 6317 36078 6343 36134
rect 6399 36078 6425 36134
rect 6481 36078 6507 36134
rect 6740 36110 6753 36134
rect 6563 36098 6589 36110
rect 6645 36098 6671 36110
rect 6727 36098 6753 36110
rect 6740 36078 6753 36098
rect 6809 36114 7472 36134
rect 6809 36078 6853 36114
rect 5820 36054 6552 36078
rect 6604 36054 6620 36078
rect 6672 36054 6688 36078
rect 6740 36058 6853 36078
rect 6909 36058 6941 36114
rect 6997 36058 7029 36114
rect 7085 36058 7117 36114
rect 7173 36058 7205 36114
rect 7261 36058 7293 36114
rect 7349 36110 7472 36114
rect 7524 36110 7540 36162
rect 7592 36110 7608 36162
rect 7660 36110 8392 36162
rect 8444 36110 8460 36162
rect 8512 36110 8528 36162
rect 8580 36110 9312 36162
rect 9364 36110 9380 36162
rect 9432 36110 9448 36162
rect 9500 36110 10232 36162
rect 10284 36110 10300 36162
rect 10352 36110 10368 36162
rect 10420 36110 11152 36162
rect 11204 36110 11220 36162
rect 11272 36110 11288 36162
rect 11340 36110 11592 36162
rect 7349 36098 11592 36110
rect 7349 36058 7472 36098
rect 6740 36054 7472 36058
rect 5661 36034 5687 36046
rect 5743 36034 5769 36046
rect 5684 35998 5687 36034
rect 4900 35982 5632 35998
rect 5684 35982 5700 35998
rect 5752 35982 5768 36034
rect 5825 35998 5851 36054
rect 5907 35998 5933 36054
rect 5989 35998 6015 36054
rect 6071 35998 6097 36054
rect 6153 35998 6179 36054
rect 6235 35998 6261 36054
rect 6317 35998 6343 36054
rect 6399 35998 6425 36054
rect 6481 35998 6507 36054
rect 6740 36046 6753 36054
rect 6563 36034 6589 36046
rect 6645 36034 6671 36046
rect 6727 36034 6753 36046
rect 6740 35998 6753 36034
rect 6809 36046 7472 36054
rect 7524 36046 7540 36098
rect 7592 36046 7608 36098
rect 7660 36046 8392 36098
rect 8444 36046 8460 36098
rect 8512 36046 8528 36098
rect 8580 36046 9312 36098
rect 9364 36046 9380 36098
rect 9432 36046 9448 36098
rect 9500 36046 10232 36098
rect 10284 36046 10300 36098
rect 10352 36046 10368 36098
rect 10420 36046 11152 36098
rect 11204 36046 11220 36098
rect 11272 36046 11288 36098
rect 11340 36046 11592 36098
rect 6809 36034 11592 36046
rect 6809 36032 7472 36034
rect 6809 35998 6853 36032
rect 5820 35982 6552 35998
rect 6604 35982 6620 35998
rect 6672 35982 6688 35998
rect 6740 35982 6853 35998
rect 2387 35979 6853 35982
rect 2387 35972 2872 35979
rect 2924 35972 2940 35979
rect 2387 35957 2538 35972
rect 187 35945 2538 35957
rect 187 35893 2231 35945
rect 2283 35893 2335 35945
rect 2387 35916 2538 35945
rect 2594 35916 2632 35972
rect 2688 35916 2726 35972
rect 2782 35916 2820 35972
rect 2992 35927 3008 35979
rect 3060 35976 6853 35979
rect 6909 35976 6941 36032
rect 6997 35976 7029 36032
rect 7085 35976 7117 36032
rect 7173 35976 7205 36032
rect 7261 35976 7293 36032
rect 7349 35982 7472 36032
rect 7524 35982 7540 36034
rect 7592 35982 7608 36034
rect 7660 35982 8392 36034
rect 8444 35982 8460 36034
rect 8512 35982 8528 36034
rect 8580 35982 9312 36034
rect 9364 35982 9380 36034
rect 9432 35982 9448 36034
rect 9500 35982 10232 36034
rect 10284 35982 10300 36034
rect 10352 35982 10368 36034
rect 10420 35982 11152 36034
rect 11204 35982 11220 36034
rect 11272 35982 11288 36034
rect 11340 35982 11592 36034
rect 7349 35976 11592 35982
rect 3060 35974 11592 35976
rect 3060 35972 3109 35974
rect 2876 35916 2914 35927
rect 2970 35916 3008 35927
rect 3064 35918 3109 35972
rect 3165 35918 3193 35974
rect 3249 35918 3277 35974
rect 3333 35918 3360 35974
rect 3416 35918 3443 35974
rect 3499 35918 3526 35974
rect 3582 35918 3609 35974
rect 3665 35918 3692 35974
rect 3748 35918 3775 35974
rect 3831 35970 3858 35974
rect 3914 35970 3941 35974
rect 3844 35918 3858 35970
rect 3914 35918 3928 35970
rect 3997 35918 4024 35974
rect 4080 35918 4107 35974
rect 4163 35918 4190 35974
rect 4246 35918 4273 35974
rect 4329 35918 4356 35974
rect 4412 35918 4439 35974
rect 4495 35918 4522 35974
rect 4578 35918 4605 35974
rect 4661 35918 4688 35974
rect 4744 35970 4771 35974
rect 4827 35970 4854 35974
rect 4764 35918 4771 35970
rect 4832 35918 4848 35970
rect 4910 35918 4937 35974
rect 4993 35918 5195 35974
rect 5251 35918 5277 35974
rect 5333 35918 5359 35974
rect 5415 35918 5441 35974
rect 5497 35918 5523 35974
rect 5579 35918 5605 35974
rect 5661 35970 5687 35974
rect 5743 35970 5769 35974
rect 5684 35918 5687 35970
rect 5752 35918 5768 35970
rect 5825 35918 5851 35974
rect 5907 35918 5933 35974
rect 5989 35918 6015 35974
rect 6071 35918 6097 35974
rect 6153 35918 6179 35974
rect 6235 35918 6261 35974
rect 6317 35918 6343 35974
rect 6399 35918 6425 35974
rect 6481 35918 6507 35974
rect 6563 35970 6589 35974
rect 6645 35970 6671 35974
rect 6727 35970 6753 35974
rect 6740 35918 6753 35970
rect 6809 35970 11592 35974
rect 6809 35950 7472 35970
rect 6809 35918 6853 35950
rect 3064 35916 6853 35918
rect 2387 35914 6853 35916
rect 2387 35893 2872 35914
rect 187 35892 2872 35893
rect 2924 35892 2940 35914
rect 187 35881 2538 35892
rect 187 35829 2231 35881
rect 2283 35829 2335 35881
rect 2387 35836 2538 35881
rect 2594 35836 2632 35892
rect 2688 35836 2726 35892
rect 2782 35836 2820 35892
rect 2992 35862 3008 35914
rect 3060 35906 6853 35914
rect 3060 35894 3792 35906
rect 3844 35894 3860 35906
rect 3912 35894 3928 35906
rect 3980 35894 4712 35906
rect 4764 35894 4780 35906
rect 3060 35892 3109 35894
rect 2876 35849 2914 35862
rect 2970 35849 3008 35862
rect 2387 35829 2872 35836
rect 187 35817 2872 35829
rect 187 35765 2231 35817
rect 2283 35765 2335 35817
rect 2387 35812 2872 35817
rect 2924 35812 2940 35836
rect 2387 35765 2538 35812
rect 187 35756 2538 35765
rect 2594 35756 2632 35812
rect 2688 35756 2726 35812
rect 2782 35756 2820 35812
rect 2992 35797 3008 35849
rect 3064 35838 3109 35892
rect 3165 35838 3193 35894
rect 3249 35838 3277 35894
rect 3333 35838 3360 35894
rect 3416 35838 3443 35894
rect 3499 35838 3526 35894
rect 3582 35838 3609 35894
rect 3665 35838 3692 35894
rect 3748 35838 3775 35894
rect 3844 35854 3858 35894
rect 3914 35854 3928 35894
rect 3831 35842 3858 35854
rect 3914 35842 3941 35854
rect 3844 35838 3858 35842
rect 3914 35838 3928 35842
rect 3997 35838 4024 35894
rect 4080 35838 4107 35894
rect 4163 35838 4190 35894
rect 4246 35838 4273 35894
rect 4329 35838 4356 35894
rect 4412 35838 4439 35894
rect 4495 35838 4522 35894
rect 4578 35838 4605 35894
rect 4661 35838 4688 35894
rect 4764 35854 4771 35894
rect 4832 35854 4848 35906
rect 4900 35894 5632 35906
rect 5684 35894 5700 35906
rect 4744 35842 4771 35854
rect 4827 35842 4854 35854
rect 4764 35838 4771 35842
rect 3064 35836 3792 35838
rect 3060 35814 3792 35836
rect 3844 35814 3860 35838
rect 3912 35814 3928 35838
rect 3980 35814 4712 35838
rect 4764 35814 4780 35838
rect 3060 35812 3109 35814
rect 2876 35784 2914 35797
rect 2970 35784 3008 35797
rect 187 35753 2872 35756
rect 187 35701 2231 35753
rect 2283 35701 2335 35753
rect 2387 35732 2872 35753
rect 2924 35732 2940 35756
rect 2992 35732 3008 35784
rect 3064 35758 3109 35812
rect 3165 35758 3193 35814
rect 3249 35758 3277 35814
rect 3333 35758 3360 35814
rect 3416 35758 3443 35814
rect 3499 35758 3526 35814
rect 3582 35758 3609 35814
rect 3665 35758 3692 35814
rect 3748 35758 3775 35814
rect 3844 35790 3858 35814
rect 3914 35790 3928 35814
rect 3831 35778 3858 35790
rect 3914 35778 3941 35790
rect 3844 35758 3858 35778
rect 3914 35758 3928 35778
rect 3997 35758 4024 35814
rect 4080 35758 4107 35814
rect 4163 35758 4190 35814
rect 4246 35758 4273 35814
rect 4329 35758 4356 35814
rect 4412 35758 4439 35814
rect 4495 35758 4522 35814
rect 4578 35758 4605 35814
rect 4661 35758 4688 35814
rect 4764 35790 4771 35814
rect 4832 35790 4848 35842
rect 4910 35838 4937 35894
rect 4993 35838 5195 35894
rect 5251 35838 5277 35894
rect 5333 35838 5359 35894
rect 5415 35838 5441 35894
rect 5497 35838 5523 35894
rect 5579 35838 5605 35894
rect 5684 35854 5687 35894
rect 5752 35854 5768 35906
rect 5820 35894 6552 35906
rect 6604 35894 6620 35906
rect 6672 35894 6688 35906
rect 6740 35894 6853 35906
rect 6909 35894 6941 35950
rect 6997 35894 7029 35950
rect 7085 35894 7117 35950
rect 7173 35894 7205 35950
rect 7261 35894 7293 35950
rect 7349 35918 7472 35950
rect 7524 35918 7540 35970
rect 7592 35918 7608 35970
rect 7660 35918 8392 35970
rect 8444 35918 8460 35970
rect 8512 35918 8528 35970
rect 8580 35918 9312 35970
rect 9364 35918 9380 35970
rect 9432 35918 9448 35970
rect 9500 35918 10232 35970
rect 10284 35918 10300 35970
rect 10352 35918 10368 35970
rect 10420 35918 11152 35970
rect 11204 35918 11220 35970
rect 11272 35918 11288 35970
rect 11340 35918 11592 35970
rect 7349 35906 11592 35918
rect 7349 35894 7472 35906
rect 5661 35842 5687 35854
rect 5743 35842 5769 35854
rect 5684 35838 5687 35842
rect 4900 35814 5632 35838
rect 5684 35814 5700 35838
rect 4744 35778 4771 35790
rect 4827 35778 4854 35790
rect 4764 35758 4771 35778
rect 3064 35756 3792 35758
rect 3060 35734 3792 35756
rect 3844 35734 3860 35758
rect 3912 35734 3928 35758
rect 3980 35734 4712 35758
rect 4764 35734 4780 35758
rect 3060 35732 3109 35734
rect 2387 35701 2538 35732
rect 187 35689 2538 35701
rect 187 35637 2231 35689
rect 2283 35637 2335 35689
rect 2387 35676 2538 35689
rect 2594 35676 2632 35732
rect 2688 35676 2726 35732
rect 2782 35676 2820 35732
rect 2876 35719 2914 35732
rect 2970 35719 3008 35732
rect 2387 35667 2872 35676
rect 2924 35667 2940 35676
rect 2992 35667 3008 35719
rect 3064 35678 3109 35732
rect 3165 35678 3193 35734
rect 3249 35678 3277 35734
rect 3333 35678 3360 35734
rect 3416 35678 3443 35734
rect 3499 35678 3526 35734
rect 3582 35678 3609 35734
rect 3665 35678 3692 35734
rect 3748 35678 3775 35734
rect 3844 35726 3858 35734
rect 3914 35726 3928 35734
rect 3831 35714 3858 35726
rect 3914 35714 3941 35726
rect 3844 35678 3858 35714
rect 3914 35678 3928 35714
rect 3997 35678 4024 35734
rect 4080 35678 4107 35734
rect 4163 35678 4190 35734
rect 4246 35678 4273 35734
rect 4329 35678 4356 35734
rect 4412 35678 4439 35734
rect 4495 35678 4522 35734
rect 4578 35678 4605 35734
rect 4661 35678 4688 35734
rect 4764 35726 4771 35734
rect 4832 35726 4848 35778
rect 4910 35758 4937 35814
rect 4993 35758 5195 35814
rect 5251 35758 5277 35814
rect 5333 35758 5359 35814
rect 5415 35758 5441 35814
rect 5497 35758 5523 35814
rect 5579 35758 5605 35814
rect 5684 35790 5687 35814
rect 5752 35790 5768 35842
rect 5825 35838 5851 35894
rect 5907 35838 5933 35894
rect 5989 35838 6015 35894
rect 6071 35838 6097 35894
rect 6153 35838 6179 35894
rect 6235 35838 6261 35894
rect 6317 35838 6343 35894
rect 6399 35838 6425 35894
rect 6481 35838 6507 35894
rect 6740 35854 6753 35894
rect 6563 35842 6589 35854
rect 6645 35842 6671 35854
rect 6727 35842 6753 35854
rect 6740 35838 6753 35842
rect 6809 35868 7472 35894
rect 6809 35838 6853 35868
rect 5820 35814 6552 35838
rect 6604 35814 6620 35838
rect 6672 35814 6688 35838
rect 6740 35814 6853 35838
rect 5661 35778 5687 35790
rect 5743 35778 5769 35790
rect 5684 35758 5687 35778
rect 4900 35734 5632 35758
rect 5684 35734 5700 35758
rect 4744 35714 4771 35726
rect 4827 35714 4854 35726
rect 4764 35678 4771 35714
rect 3064 35676 3792 35678
rect 3060 35667 3792 35676
rect 2387 35662 3792 35667
rect 3844 35662 3860 35678
rect 3912 35662 3928 35678
rect 3980 35662 4712 35678
rect 4764 35662 4780 35678
rect 4832 35662 4848 35714
rect 4910 35678 4937 35734
rect 4993 35678 5195 35734
rect 5251 35678 5277 35734
rect 5333 35678 5359 35734
rect 5415 35678 5441 35734
rect 5497 35678 5523 35734
rect 5579 35678 5605 35734
rect 5684 35726 5687 35734
rect 5752 35726 5768 35778
rect 5825 35758 5851 35814
rect 5907 35758 5933 35814
rect 5989 35758 6015 35814
rect 6071 35758 6097 35814
rect 6153 35758 6179 35814
rect 6235 35758 6261 35814
rect 6317 35758 6343 35814
rect 6399 35758 6425 35814
rect 6481 35758 6507 35814
rect 6740 35790 6753 35814
rect 6563 35778 6589 35790
rect 6645 35778 6671 35790
rect 6727 35778 6753 35790
rect 6740 35758 6753 35778
rect 6809 35812 6853 35814
rect 6909 35812 6941 35868
rect 6997 35812 7029 35868
rect 7085 35812 7117 35868
rect 7173 35812 7205 35868
rect 7261 35812 7293 35868
rect 7349 35854 7472 35868
rect 7524 35854 7540 35906
rect 7592 35854 7608 35906
rect 7660 35854 8392 35906
rect 8444 35854 8460 35906
rect 8512 35854 8528 35906
rect 8580 35854 9312 35906
rect 9364 35854 9380 35906
rect 9432 35854 9448 35906
rect 9500 35854 10232 35906
rect 10284 35854 10300 35906
rect 10352 35854 10368 35906
rect 10420 35854 11152 35906
rect 11204 35854 11220 35906
rect 11272 35854 11288 35906
rect 11340 35854 11592 35906
rect 7349 35842 11592 35854
rect 7349 35812 7472 35842
rect 6809 35790 7472 35812
rect 7524 35790 7540 35842
rect 7592 35790 7608 35842
rect 7660 35790 8392 35842
rect 8444 35790 8460 35842
rect 8512 35790 8528 35842
rect 8580 35790 9312 35842
rect 9364 35790 9380 35842
rect 9432 35790 9448 35842
rect 9500 35790 10232 35842
rect 10284 35790 10300 35842
rect 10352 35790 10368 35842
rect 10420 35790 11152 35842
rect 11204 35790 11220 35842
rect 11272 35790 11288 35842
rect 11340 35790 11592 35842
rect 6809 35786 11592 35790
rect 6809 35758 6853 35786
rect 5820 35734 6552 35758
rect 6604 35734 6620 35758
rect 6672 35734 6688 35758
rect 6740 35734 6853 35758
rect 5661 35714 5687 35726
rect 5743 35714 5769 35726
rect 5684 35678 5687 35714
rect 4900 35662 5632 35678
rect 5684 35662 5700 35678
rect 5752 35662 5768 35714
rect 5825 35678 5851 35734
rect 5907 35678 5933 35734
rect 5989 35678 6015 35734
rect 6071 35678 6097 35734
rect 6153 35678 6179 35734
rect 6235 35678 6261 35734
rect 6317 35678 6343 35734
rect 6399 35678 6425 35734
rect 6481 35678 6507 35734
rect 6740 35726 6753 35734
rect 6563 35714 6589 35726
rect 6645 35714 6671 35726
rect 6727 35714 6753 35726
rect 6740 35678 6753 35714
rect 6809 35730 6853 35734
rect 6909 35730 6941 35786
rect 6997 35730 7029 35786
rect 7085 35730 7117 35786
rect 7173 35730 7205 35786
rect 7261 35730 7293 35786
rect 7349 35778 11592 35786
rect 7349 35730 7472 35778
rect 6809 35726 7472 35730
rect 7524 35726 7540 35778
rect 7592 35726 7608 35778
rect 7660 35726 8392 35778
rect 8444 35726 8460 35778
rect 8512 35726 8528 35778
rect 8580 35726 9312 35778
rect 9364 35726 9380 35778
rect 9432 35726 9448 35778
rect 9500 35726 10232 35778
rect 10284 35726 10300 35778
rect 10352 35726 10368 35778
rect 10420 35726 11152 35778
rect 11204 35726 11220 35778
rect 11272 35726 11288 35778
rect 11340 35726 11592 35778
rect 6809 35714 11592 35726
rect 6809 35704 7472 35714
rect 6809 35678 6853 35704
rect 5820 35662 6552 35678
rect 6604 35662 6620 35678
rect 6672 35662 6688 35678
rect 6740 35662 6853 35678
rect 2387 35654 6853 35662
rect 2387 35652 2872 35654
rect 2924 35652 2940 35654
rect 2387 35637 2538 35652
rect 187 35625 2538 35637
rect 187 35573 2231 35625
rect 2283 35573 2335 35625
rect 2387 35596 2538 35625
rect 2594 35596 2632 35652
rect 2688 35596 2726 35652
rect 2782 35596 2820 35652
rect 2992 35602 3008 35654
rect 3060 35652 3109 35654
rect 2876 35596 2914 35602
rect 2970 35596 3008 35602
rect 3064 35598 3109 35652
rect 3165 35598 3193 35654
rect 3249 35598 3277 35654
rect 3333 35598 3360 35654
rect 3416 35598 3443 35654
rect 3499 35598 3526 35654
rect 3582 35598 3609 35654
rect 3665 35598 3692 35654
rect 3748 35598 3775 35654
rect 3831 35650 3858 35654
rect 3914 35650 3941 35654
rect 3844 35598 3858 35650
rect 3914 35598 3928 35650
rect 3997 35598 4024 35654
rect 4080 35598 4107 35654
rect 4163 35598 4190 35654
rect 4246 35598 4273 35654
rect 4329 35598 4356 35654
rect 4412 35598 4439 35654
rect 4495 35598 4522 35654
rect 4578 35598 4605 35654
rect 4661 35598 4688 35654
rect 4744 35650 4771 35654
rect 4827 35650 4854 35654
rect 4764 35598 4771 35650
rect 4832 35598 4848 35650
rect 4910 35598 4937 35654
rect 4993 35598 5195 35654
rect 5251 35598 5277 35654
rect 5333 35598 5359 35654
rect 5415 35598 5441 35654
rect 5497 35598 5523 35654
rect 5579 35598 5605 35654
rect 5661 35650 5687 35654
rect 5743 35650 5769 35654
rect 5684 35598 5687 35650
rect 5752 35598 5768 35650
rect 5825 35598 5851 35654
rect 5907 35598 5933 35654
rect 5989 35598 6015 35654
rect 6071 35598 6097 35654
rect 6153 35598 6179 35654
rect 6235 35598 6261 35654
rect 6317 35598 6343 35654
rect 6399 35598 6425 35654
rect 6481 35598 6507 35654
rect 6563 35650 6589 35654
rect 6645 35650 6671 35654
rect 6727 35650 6753 35654
rect 6740 35598 6753 35650
rect 6809 35648 6853 35654
rect 6909 35648 6941 35704
rect 6997 35648 7029 35704
rect 7085 35648 7117 35704
rect 7173 35648 7205 35704
rect 7261 35648 7293 35704
rect 7349 35662 7472 35704
rect 7524 35662 7540 35714
rect 7592 35662 7608 35714
rect 7660 35662 8392 35714
rect 8444 35662 8460 35714
rect 8512 35662 8528 35714
rect 8580 35662 9312 35714
rect 9364 35662 9380 35714
rect 9432 35662 9448 35714
rect 9500 35662 10232 35714
rect 10284 35662 10300 35714
rect 10352 35662 10368 35714
rect 10420 35662 11152 35714
rect 11204 35662 11220 35714
rect 11272 35662 11288 35714
rect 11340 35662 11592 35714
rect 7349 35650 11592 35662
rect 7349 35648 7472 35650
rect 6809 35622 7472 35648
rect 6809 35598 6853 35622
rect 3064 35596 6853 35598
rect 2387 35589 6853 35596
rect 2387 35573 2872 35589
rect 187 35572 2872 35573
rect 2924 35572 2940 35589
rect 187 35561 2538 35572
rect 187 35509 2231 35561
rect 2283 35509 2335 35561
rect 2387 35516 2538 35561
rect 2594 35516 2632 35572
rect 2688 35516 2726 35572
rect 2782 35516 2820 35572
rect 2992 35537 3008 35589
rect 3060 35586 6853 35589
rect 3060 35574 3792 35586
rect 3844 35574 3860 35586
rect 3912 35574 3928 35586
rect 3980 35574 4712 35586
rect 4764 35574 4780 35586
rect 3060 35572 3109 35574
rect 2876 35524 2914 35537
rect 2970 35524 3008 35537
rect 2387 35509 2872 35516
rect 187 35497 2872 35509
rect 187 35445 2231 35497
rect 2283 35445 2335 35497
rect 2387 35491 2872 35497
rect 2924 35491 2940 35516
rect 2387 35445 2538 35491
rect 187 35435 2538 35445
rect 2594 35435 2632 35491
rect 2688 35435 2726 35491
rect 2782 35435 2820 35491
rect 2992 35472 3008 35524
rect 3064 35518 3109 35572
rect 3165 35518 3193 35574
rect 3249 35518 3277 35574
rect 3333 35518 3360 35574
rect 3416 35518 3443 35574
rect 3499 35518 3526 35574
rect 3582 35518 3609 35574
rect 3665 35518 3692 35574
rect 3748 35518 3775 35574
rect 3844 35534 3858 35574
rect 3914 35534 3928 35574
rect 3831 35522 3858 35534
rect 3914 35522 3941 35534
rect 3844 35518 3858 35522
rect 3914 35518 3928 35522
rect 3997 35518 4024 35574
rect 4080 35518 4107 35574
rect 4163 35518 4190 35574
rect 4246 35518 4273 35574
rect 4329 35518 4356 35574
rect 4412 35518 4439 35574
rect 4495 35518 4522 35574
rect 4578 35518 4605 35574
rect 4661 35518 4688 35574
rect 4764 35534 4771 35574
rect 4832 35534 4848 35586
rect 4900 35574 5632 35586
rect 5684 35574 5700 35586
rect 4744 35522 4771 35534
rect 4827 35522 4854 35534
rect 4764 35518 4771 35522
rect 3064 35516 3792 35518
rect 3060 35494 3792 35516
rect 3844 35494 3860 35518
rect 3912 35494 3928 35518
rect 3980 35494 4712 35518
rect 4764 35494 4780 35518
rect 3060 35491 3109 35494
rect 2876 35459 2914 35472
rect 2970 35459 3008 35472
rect 187 35433 2872 35435
rect 187 35381 2231 35433
rect 2283 35381 2335 35433
rect 2387 35410 2872 35433
rect 2924 35410 2940 35435
rect 2387 35381 2538 35410
rect 187 35369 2538 35381
rect 187 35317 2231 35369
rect 2283 35317 2335 35369
rect 2387 35354 2538 35369
rect 2594 35354 2632 35410
rect 2688 35354 2726 35410
rect 2782 35354 2820 35410
rect 2992 35407 3008 35459
rect 3064 35438 3109 35491
rect 3165 35438 3193 35494
rect 3249 35438 3277 35494
rect 3333 35438 3360 35494
rect 3416 35438 3443 35494
rect 3499 35438 3526 35494
rect 3582 35438 3609 35494
rect 3665 35438 3692 35494
rect 3748 35438 3775 35494
rect 3844 35470 3858 35494
rect 3914 35470 3928 35494
rect 3831 35458 3858 35470
rect 3914 35458 3941 35470
rect 3844 35438 3858 35458
rect 3914 35438 3928 35458
rect 3997 35438 4024 35494
rect 4080 35438 4107 35494
rect 4163 35438 4190 35494
rect 4246 35438 4273 35494
rect 4329 35438 4356 35494
rect 4412 35438 4439 35494
rect 4495 35438 4522 35494
rect 4578 35438 4605 35494
rect 4661 35438 4688 35494
rect 4764 35470 4771 35494
rect 4832 35470 4848 35522
rect 4910 35518 4937 35574
rect 4993 35518 5195 35574
rect 5251 35518 5277 35574
rect 5333 35518 5359 35574
rect 5415 35518 5441 35574
rect 5497 35518 5523 35574
rect 5579 35518 5605 35574
rect 5684 35534 5687 35574
rect 5752 35534 5768 35586
rect 5820 35574 6552 35586
rect 6604 35574 6620 35586
rect 6672 35574 6688 35586
rect 6740 35574 6853 35586
rect 5661 35522 5687 35534
rect 5743 35522 5769 35534
rect 5684 35518 5687 35522
rect 4900 35494 5632 35518
rect 5684 35494 5700 35518
rect 4744 35458 4771 35470
rect 4827 35458 4854 35470
rect 4764 35438 4771 35458
rect 3064 35435 3792 35438
rect 3060 35414 3792 35435
rect 3844 35414 3860 35438
rect 3912 35414 3928 35438
rect 3980 35414 4712 35438
rect 4764 35414 4780 35438
rect 3060 35410 3109 35414
rect 2876 35394 2914 35407
rect 2970 35394 3008 35407
rect 2387 35342 2872 35354
rect 2924 35342 2940 35354
rect 2992 35342 3008 35394
rect 3064 35358 3109 35410
rect 3165 35358 3193 35414
rect 3249 35358 3277 35414
rect 3333 35358 3360 35414
rect 3416 35358 3443 35414
rect 3499 35358 3526 35414
rect 3582 35358 3609 35414
rect 3665 35358 3692 35414
rect 3748 35358 3775 35414
rect 3844 35406 3858 35414
rect 3914 35406 3928 35414
rect 3831 35394 3858 35406
rect 3914 35394 3941 35406
rect 3844 35358 3858 35394
rect 3914 35358 3928 35394
rect 3997 35358 4024 35414
rect 4080 35358 4107 35414
rect 4163 35358 4190 35414
rect 4246 35358 4273 35414
rect 4329 35358 4356 35414
rect 4412 35358 4439 35414
rect 4495 35358 4522 35414
rect 4578 35358 4605 35414
rect 4661 35358 4688 35414
rect 4764 35406 4771 35414
rect 4832 35406 4848 35458
rect 4910 35438 4937 35494
rect 4993 35438 5195 35494
rect 5251 35438 5277 35494
rect 5333 35438 5359 35494
rect 5415 35438 5441 35494
rect 5497 35438 5523 35494
rect 5579 35438 5605 35494
rect 5684 35470 5687 35494
rect 5752 35470 5768 35522
rect 5825 35518 5851 35574
rect 5907 35518 5933 35574
rect 5989 35518 6015 35574
rect 6071 35518 6097 35574
rect 6153 35518 6179 35574
rect 6235 35518 6261 35574
rect 6317 35518 6343 35574
rect 6399 35518 6425 35574
rect 6481 35518 6507 35574
rect 6740 35534 6753 35574
rect 6563 35522 6589 35534
rect 6645 35522 6671 35534
rect 6727 35522 6753 35534
rect 6740 35518 6753 35522
rect 6809 35566 6853 35574
rect 6909 35566 6941 35622
rect 6997 35566 7029 35622
rect 7085 35566 7117 35622
rect 7173 35566 7205 35622
rect 7261 35566 7293 35622
rect 7349 35598 7472 35622
rect 7524 35598 7540 35650
rect 7592 35598 7608 35650
rect 7660 35598 8392 35650
rect 8444 35598 8460 35650
rect 8512 35598 8528 35650
rect 8580 35598 9312 35650
rect 9364 35598 9380 35650
rect 9432 35598 9448 35650
rect 9500 35598 10232 35650
rect 10284 35598 10300 35650
rect 10352 35598 10368 35650
rect 10420 35598 11152 35650
rect 11204 35598 11220 35650
rect 11272 35598 11288 35650
rect 11340 35598 11592 35650
rect 7349 35586 11592 35598
rect 7349 35566 7472 35586
rect 6809 35539 7472 35566
rect 6809 35518 6853 35539
rect 5820 35494 6552 35518
rect 6604 35494 6620 35518
rect 6672 35494 6688 35518
rect 6740 35494 6853 35518
rect 5661 35458 5687 35470
rect 5743 35458 5769 35470
rect 5684 35438 5687 35458
rect 4900 35414 5632 35438
rect 5684 35414 5700 35438
rect 4744 35394 4771 35406
rect 4827 35394 4854 35406
rect 4764 35358 4771 35394
rect 3064 35354 3792 35358
rect 3060 35342 3792 35354
rect 3844 35342 3860 35358
rect 3912 35342 3928 35358
rect 3980 35342 4712 35358
rect 4764 35342 4780 35358
rect 4832 35342 4848 35394
rect 4910 35358 4937 35414
rect 4993 35358 5195 35414
rect 5251 35358 5277 35414
rect 5333 35358 5359 35414
rect 5415 35358 5441 35414
rect 5497 35358 5523 35414
rect 5579 35358 5605 35414
rect 5684 35406 5687 35414
rect 5752 35406 5768 35458
rect 5825 35438 5851 35494
rect 5907 35438 5933 35494
rect 5989 35438 6015 35494
rect 6071 35438 6097 35494
rect 6153 35438 6179 35494
rect 6235 35438 6261 35494
rect 6317 35438 6343 35494
rect 6399 35438 6425 35494
rect 6481 35438 6507 35494
rect 6740 35470 6753 35494
rect 6563 35458 6589 35470
rect 6645 35458 6671 35470
rect 6727 35458 6753 35470
rect 6740 35438 6753 35458
rect 6809 35483 6853 35494
rect 6909 35483 6941 35539
rect 6997 35483 7029 35539
rect 7085 35483 7117 35539
rect 7173 35483 7205 35539
rect 7261 35483 7293 35539
rect 7349 35534 7472 35539
rect 7524 35534 7540 35586
rect 7592 35534 7608 35586
rect 7660 35534 8392 35586
rect 8444 35534 8460 35586
rect 8512 35534 8528 35586
rect 8580 35534 9312 35586
rect 9364 35534 9380 35586
rect 9432 35534 9448 35586
rect 9500 35534 10232 35586
rect 10284 35534 10300 35586
rect 10352 35534 10368 35586
rect 10420 35534 11152 35586
rect 11204 35534 11220 35586
rect 11272 35534 11288 35586
rect 11340 35534 11592 35586
rect 7349 35522 11592 35534
rect 7349 35483 7472 35522
rect 6809 35470 7472 35483
rect 7524 35470 7540 35522
rect 7592 35470 7608 35522
rect 7660 35470 8392 35522
rect 8444 35470 8460 35522
rect 8512 35470 8528 35522
rect 8580 35470 9312 35522
rect 9364 35470 9380 35522
rect 9432 35470 9448 35522
rect 9500 35470 10232 35522
rect 10284 35470 10300 35522
rect 10352 35470 10368 35522
rect 10420 35470 11152 35522
rect 11204 35470 11220 35522
rect 11272 35470 11288 35522
rect 11340 35470 11592 35522
rect 6809 35458 11592 35470
rect 6809 35456 7472 35458
rect 6809 35438 6853 35456
rect 5820 35414 6552 35438
rect 6604 35414 6620 35438
rect 6672 35414 6688 35438
rect 6740 35414 6853 35438
rect 5661 35394 5687 35406
rect 5743 35394 5769 35406
rect 5684 35358 5687 35394
rect 4900 35342 5632 35358
rect 5684 35342 5700 35358
rect 5752 35342 5768 35394
rect 5825 35358 5851 35414
rect 5907 35358 5933 35414
rect 5989 35358 6015 35414
rect 6071 35358 6097 35414
rect 6153 35358 6179 35414
rect 6235 35358 6261 35414
rect 6317 35358 6343 35414
rect 6399 35358 6425 35414
rect 6481 35358 6507 35414
rect 6740 35406 6753 35414
rect 6563 35394 6589 35406
rect 6645 35394 6671 35406
rect 6727 35394 6753 35406
rect 6740 35358 6753 35394
rect 6809 35400 6853 35414
rect 6909 35400 6941 35456
rect 6997 35400 7029 35456
rect 7085 35400 7117 35456
rect 7173 35400 7205 35456
rect 7261 35400 7293 35456
rect 7349 35406 7472 35456
rect 7524 35406 7540 35458
rect 7592 35406 7608 35458
rect 7660 35406 8392 35458
rect 8444 35406 8460 35458
rect 8512 35406 8528 35458
rect 8580 35406 9312 35458
rect 9364 35406 9380 35458
rect 9432 35406 9448 35458
rect 9500 35406 10232 35458
rect 10284 35406 10300 35458
rect 10352 35406 10368 35458
rect 10420 35406 11152 35458
rect 11204 35406 11220 35458
rect 11272 35406 11288 35458
rect 11340 35406 11592 35458
rect 7349 35400 11592 35406
rect 6809 35394 11592 35400
rect 6809 35373 7472 35394
rect 6809 35358 6853 35373
rect 5820 35342 6552 35358
rect 6604 35342 6620 35358
rect 6672 35342 6688 35358
rect 6740 35342 6853 35358
rect 2387 35334 6853 35342
rect 2387 35329 3109 35334
rect 2387 35317 2538 35329
rect 187 35305 2538 35317
rect 187 35253 2231 35305
rect 2283 35253 2335 35305
rect 2387 35273 2538 35305
rect 2594 35273 2632 35329
rect 2688 35273 2726 35329
rect 2782 35273 2820 35329
rect 2992 35277 3008 35329
rect 3064 35278 3109 35329
rect 3165 35278 3193 35334
rect 3249 35278 3277 35334
rect 3333 35278 3360 35334
rect 3416 35278 3443 35334
rect 3499 35278 3526 35334
rect 3582 35278 3609 35334
rect 3665 35278 3692 35334
rect 3748 35278 3775 35334
rect 3831 35329 3858 35334
rect 3914 35329 3941 35334
rect 3844 35278 3858 35329
rect 3914 35278 3928 35329
rect 3997 35278 4024 35334
rect 4080 35278 4107 35334
rect 4163 35278 4190 35334
rect 4246 35278 4273 35334
rect 4329 35278 4356 35334
rect 4412 35278 4439 35334
rect 4495 35278 4522 35334
rect 4578 35278 4605 35334
rect 4661 35278 4688 35334
rect 4744 35329 4771 35334
rect 4827 35329 4854 35334
rect 4764 35278 4771 35329
rect 3064 35277 3792 35278
rect 3844 35277 3860 35278
rect 3912 35277 3928 35278
rect 3980 35277 4712 35278
rect 4764 35277 4780 35278
rect 4832 35277 4848 35329
rect 4910 35278 4937 35334
rect 4993 35278 5195 35334
rect 5251 35278 5277 35334
rect 5333 35278 5359 35334
rect 5415 35278 5441 35334
rect 5497 35278 5523 35334
rect 5579 35278 5605 35334
rect 5661 35329 5687 35334
rect 5743 35329 5769 35334
rect 5684 35278 5687 35329
rect 4900 35277 5632 35278
rect 5684 35277 5700 35278
rect 5752 35277 5768 35329
rect 5825 35278 5851 35334
rect 5907 35278 5933 35334
rect 5989 35278 6015 35334
rect 6071 35278 6097 35334
rect 6153 35278 6179 35334
rect 6235 35278 6261 35334
rect 6317 35278 6343 35334
rect 6399 35278 6425 35334
rect 6481 35278 6507 35334
rect 6563 35329 6589 35334
rect 6645 35329 6671 35334
rect 6727 35329 6753 35334
rect 6740 35278 6753 35329
rect 6809 35317 6853 35334
rect 6909 35317 6941 35373
rect 6997 35317 7029 35373
rect 7085 35317 7117 35373
rect 7173 35317 7205 35373
rect 7261 35317 7293 35373
rect 7349 35342 7472 35373
rect 7524 35342 7540 35394
rect 7592 35342 7608 35394
rect 7660 35342 8392 35394
rect 8444 35342 8460 35394
rect 8512 35342 8528 35394
rect 8580 35342 9312 35394
rect 9364 35342 9380 35394
rect 9432 35342 9448 35394
rect 9500 35342 10232 35394
rect 10284 35342 10300 35394
rect 10352 35342 10368 35394
rect 10420 35342 11152 35394
rect 11204 35342 11220 35394
rect 11272 35342 11288 35394
rect 11340 35342 11592 35394
rect 7349 35329 11592 35342
rect 7349 35317 7472 35329
rect 6809 35290 7472 35317
rect 6809 35278 6853 35290
rect 5820 35277 6552 35278
rect 6604 35277 6620 35278
rect 6672 35277 6688 35278
rect 6740 35277 6853 35278
rect 2876 35273 2914 35277
rect 2970 35273 3008 35277
rect 3064 35273 6853 35277
rect 2387 35264 6853 35273
rect 2387 35253 2872 35264
rect 187 35248 2872 35253
rect 2924 35248 2940 35264
rect 187 35241 2538 35248
rect 187 35189 2231 35241
rect 2283 35189 2335 35241
rect 2387 35192 2538 35241
rect 2594 35192 2632 35248
rect 2688 35192 2726 35248
rect 2782 35192 2820 35248
rect 2992 35212 3008 35264
rect 3060 35254 3792 35264
rect 3844 35254 3860 35264
rect 3912 35254 3928 35264
rect 3980 35254 4712 35264
rect 4764 35254 4780 35264
rect 3060 35248 3109 35254
rect 2876 35199 2914 35212
rect 2970 35199 3008 35212
rect 2387 35189 2872 35192
rect 187 35176 2872 35189
rect 187 35124 2231 35176
rect 2283 35124 2335 35176
rect 2387 35150 2872 35176
rect 2924 35150 2940 35192
rect 2992 35150 3008 35199
rect 3064 35198 3109 35248
rect 3165 35198 3193 35254
rect 3249 35198 3277 35254
rect 3333 35198 3360 35254
rect 3416 35198 3443 35254
rect 3499 35198 3526 35254
rect 3582 35198 3609 35254
rect 3665 35198 3692 35254
rect 3748 35198 3775 35254
rect 3844 35212 3858 35254
rect 3914 35212 3928 35254
rect 3831 35199 3858 35212
rect 3914 35199 3941 35212
rect 3844 35198 3858 35199
rect 3914 35198 3928 35199
rect 3997 35198 4024 35254
rect 4080 35198 4107 35254
rect 4163 35198 4190 35254
rect 4246 35198 4273 35254
rect 4329 35198 4356 35254
rect 4412 35198 4439 35254
rect 4495 35198 4522 35254
rect 4578 35198 4605 35254
rect 4661 35198 4688 35254
rect 4764 35212 4771 35254
rect 4832 35212 4848 35264
rect 4900 35254 5632 35264
rect 5684 35254 5700 35264
rect 4744 35199 4771 35212
rect 4827 35199 4854 35212
rect 4764 35198 4771 35199
rect 3064 35192 3792 35198
rect 3060 35174 3792 35192
rect 3844 35174 3860 35198
rect 3912 35174 3928 35198
rect 3980 35174 4712 35198
rect 4764 35174 4780 35198
rect 3060 35150 3109 35174
rect 2387 35139 2821 35150
rect 2992 35147 3006 35150
rect 2387 35124 2675 35139
rect 187 35111 2675 35124
rect 187 35059 2231 35111
rect 2283 35059 2335 35111
rect 2387 35083 2675 35111
rect 2731 35094 2821 35139
rect 2877 35134 2914 35147
rect 2970 35134 3006 35147
rect 2992 35094 3006 35134
rect 3062 35118 3109 35150
rect 3165 35118 3193 35174
rect 3249 35118 3277 35174
rect 3333 35118 3360 35174
rect 3416 35118 3443 35174
rect 3499 35118 3526 35174
rect 3582 35118 3609 35174
rect 3665 35118 3692 35174
rect 3748 35118 3775 35174
rect 3844 35147 3858 35174
rect 3914 35147 3928 35174
rect 3831 35134 3858 35147
rect 3914 35134 3941 35147
rect 3844 35118 3858 35134
rect 3914 35118 3928 35134
rect 3997 35118 4024 35174
rect 4080 35118 4107 35174
rect 4163 35118 4190 35174
rect 4246 35118 4273 35174
rect 4329 35118 4356 35174
rect 4412 35118 4439 35174
rect 4495 35118 4522 35174
rect 4578 35118 4605 35174
rect 4661 35118 4688 35174
rect 4764 35147 4771 35174
rect 4832 35147 4848 35199
rect 4910 35198 4937 35254
rect 4993 35198 5195 35254
rect 5251 35198 5277 35254
rect 5333 35198 5359 35254
rect 5415 35198 5441 35254
rect 5497 35198 5523 35254
rect 5579 35198 5605 35254
rect 5684 35212 5687 35254
rect 5752 35212 5768 35264
rect 5820 35254 6552 35264
rect 6604 35254 6620 35264
rect 6672 35254 6688 35264
rect 6740 35254 6853 35264
rect 5661 35199 5687 35212
rect 5743 35199 5769 35212
rect 5684 35198 5687 35199
rect 4900 35174 5632 35198
rect 5684 35174 5700 35198
rect 4744 35134 4771 35147
rect 4827 35134 4854 35147
rect 4764 35118 4771 35134
rect 3062 35094 3792 35118
rect 3844 35094 3860 35118
rect 3912 35094 3928 35118
rect 3980 35094 4712 35118
rect 4764 35094 4780 35118
rect 2731 35083 2872 35094
rect 2387 35082 2872 35083
rect 2924 35082 2940 35094
rect 2992 35082 3008 35094
rect 3060 35082 3109 35094
rect 2387 35069 3109 35082
rect 2387 35059 2872 35069
rect 187 35058 2872 35059
rect 2924 35058 2940 35069
rect 2992 35058 3008 35069
rect 3060 35058 3109 35069
rect 187 35046 2821 35058
rect 187 34994 2231 35046
rect 2283 34994 2335 35046
rect 2387 35002 2821 35046
rect 2992 35017 3006 35058
rect 3062 35038 3109 35058
rect 3165 35038 3193 35094
rect 3249 35038 3277 35094
rect 3333 35038 3360 35094
rect 3416 35038 3443 35094
rect 3499 35038 3526 35094
rect 3582 35038 3609 35094
rect 3665 35038 3692 35094
rect 3748 35038 3775 35094
rect 3844 35082 3858 35094
rect 3914 35082 3928 35094
rect 3831 35069 3858 35082
rect 3914 35069 3941 35082
rect 3844 35038 3858 35069
rect 3914 35038 3928 35069
rect 3997 35038 4024 35094
rect 4080 35038 4107 35094
rect 4163 35038 4190 35094
rect 4246 35038 4273 35094
rect 4329 35038 4356 35094
rect 4412 35038 4439 35094
rect 4495 35038 4522 35094
rect 4578 35038 4605 35094
rect 4661 35038 4688 35094
rect 4764 35082 4771 35094
rect 4832 35082 4848 35134
rect 4910 35118 4937 35174
rect 4993 35118 5195 35174
rect 5251 35118 5277 35174
rect 5333 35118 5359 35174
rect 5415 35118 5441 35174
rect 5497 35118 5523 35174
rect 5579 35118 5605 35174
rect 5684 35147 5687 35174
rect 5752 35147 5768 35199
rect 5825 35198 5851 35254
rect 5907 35198 5933 35254
rect 5989 35198 6015 35254
rect 6071 35198 6097 35254
rect 6153 35198 6179 35254
rect 6235 35198 6261 35254
rect 6317 35198 6343 35254
rect 6399 35198 6425 35254
rect 6481 35198 6507 35254
rect 6740 35212 6753 35254
rect 6563 35199 6589 35212
rect 6645 35199 6671 35212
rect 6727 35199 6753 35212
rect 6740 35198 6753 35199
rect 6809 35234 6853 35254
rect 6909 35234 6941 35290
rect 6997 35234 7029 35290
rect 7085 35234 7117 35290
rect 7173 35234 7205 35290
rect 7261 35234 7293 35290
rect 7349 35277 7472 35290
rect 7524 35277 7540 35329
rect 7592 35277 7608 35329
rect 7660 35277 8392 35329
rect 8444 35277 8460 35329
rect 8512 35277 8528 35329
rect 8580 35277 9312 35329
rect 9364 35277 9380 35329
rect 9432 35277 9448 35329
rect 9500 35277 10232 35329
rect 10284 35277 10300 35329
rect 10352 35277 10368 35329
rect 10420 35277 11152 35329
rect 11204 35277 11220 35329
rect 11272 35277 11288 35329
rect 11340 35277 11592 35329
rect 7349 35264 11592 35277
rect 7349 35234 7472 35264
rect 6809 35212 7472 35234
rect 7524 35212 7540 35264
rect 7592 35212 7608 35264
rect 7660 35212 8392 35264
rect 8444 35212 8460 35264
rect 8512 35212 8528 35264
rect 8580 35212 9312 35264
rect 9364 35212 9380 35264
rect 9432 35212 9448 35264
rect 9500 35212 10232 35264
rect 10284 35212 10300 35264
rect 10352 35212 10368 35264
rect 10420 35212 11152 35264
rect 11204 35212 11220 35264
rect 11272 35212 11288 35264
rect 11340 35212 11592 35264
rect 6809 35207 11592 35212
rect 6809 35198 6853 35207
rect 5820 35174 6552 35198
rect 6604 35174 6620 35198
rect 6672 35174 6688 35198
rect 6740 35174 6853 35198
rect 5661 35134 5687 35147
rect 5743 35134 5769 35147
rect 5684 35118 5687 35134
rect 4900 35094 5632 35118
rect 5684 35094 5700 35118
rect 4744 35069 4771 35082
rect 4827 35069 4854 35082
rect 4764 35038 4771 35069
rect 3062 35017 3792 35038
rect 3844 35017 3860 35038
rect 3912 35017 3928 35038
rect 3980 35017 4712 35038
rect 4764 35017 4780 35038
rect 4832 35017 4848 35069
rect 4910 35038 4937 35094
rect 4993 35038 5195 35094
rect 5251 35038 5277 35094
rect 5333 35038 5359 35094
rect 5415 35038 5441 35094
rect 5497 35038 5523 35094
rect 5579 35038 5605 35094
rect 5684 35082 5687 35094
rect 5752 35082 5768 35134
rect 5825 35118 5851 35174
rect 5907 35118 5933 35174
rect 5989 35118 6015 35174
rect 6071 35118 6097 35174
rect 6153 35118 6179 35174
rect 6235 35118 6261 35174
rect 6317 35118 6343 35174
rect 6399 35118 6425 35174
rect 6481 35118 6507 35174
rect 6740 35147 6753 35174
rect 6563 35134 6589 35147
rect 6645 35134 6671 35147
rect 6727 35134 6753 35147
rect 6740 35118 6753 35134
rect 6809 35151 6853 35174
rect 6909 35151 6941 35207
rect 6997 35151 7029 35207
rect 7085 35151 7117 35207
rect 7173 35151 7205 35207
rect 7261 35151 7293 35207
rect 7349 35199 11592 35207
rect 7349 35151 7472 35199
rect 6809 35147 7472 35151
rect 7524 35147 7540 35199
rect 7592 35147 7608 35199
rect 7660 35147 8392 35199
rect 8444 35147 8460 35199
rect 8512 35147 8528 35199
rect 8580 35147 9312 35199
rect 9364 35147 9380 35199
rect 9432 35147 9448 35199
rect 9500 35147 10232 35199
rect 10284 35147 10300 35199
rect 10352 35147 10368 35199
rect 10420 35147 11152 35199
rect 11204 35147 11220 35199
rect 11272 35147 11288 35199
rect 11340 35147 11592 35199
rect 6809 35134 11592 35147
rect 6809 35124 7472 35134
rect 6809 35118 6853 35124
rect 5820 35094 6552 35118
rect 6604 35094 6620 35118
rect 6672 35094 6688 35118
rect 6740 35094 6853 35118
rect 5661 35069 5687 35082
rect 5743 35069 5769 35082
rect 5684 35038 5687 35069
rect 4900 35017 5632 35038
rect 5684 35017 5700 35038
rect 5752 35017 5768 35069
rect 5825 35038 5851 35094
rect 5907 35038 5933 35094
rect 5989 35038 6015 35094
rect 6071 35038 6097 35094
rect 6153 35038 6179 35094
rect 6235 35038 6261 35094
rect 6317 35038 6343 35094
rect 6399 35038 6425 35094
rect 6481 35038 6507 35094
rect 6740 35082 6753 35094
rect 6563 35069 6589 35082
rect 6645 35069 6671 35082
rect 6727 35069 6753 35082
rect 6740 35038 6753 35069
rect 6809 35068 6853 35094
rect 6909 35068 6941 35124
rect 6997 35068 7029 35124
rect 7085 35068 7117 35124
rect 7173 35068 7205 35124
rect 7261 35068 7293 35124
rect 7349 35082 7472 35124
rect 7524 35082 7540 35134
rect 7592 35082 7608 35134
rect 7660 35082 8392 35134
rect 8444 35082 8460 35134
rect 8512 35082 8528 35134
rect 8580 35082 9312 35134
rect 9364 35082 9380 35134
rect 9432 35082 9448 35134
rect 9500 35082 10232 35134
rect 10284 35082 10300 35134
rect 10352 35082 10368 35134
rect 10420 35082 11152 35134
rect 11204 35082 11220 35134
rect 11272 35082 11288 35134
rect 11340 35082 11592 35134
rect 7349 35069 11592 35082
rect 7349 35068 7472 35069
rect 6809 35038 7472 35068
rect 5820 35017 6552 35038
rect 6604 35017 6620 35038
rect 6672 35017 6688 35038
rect 6740 35017 7472 35038
rect 7524 35017 7540 35069
rect 7592 35017 7608 35069
rect 7660 35017 8392 35069
rect 8444 35017 8460 35069
rect 8512 35017 8528 35069
rect 8580 35017 9312 35069
rect 9364 35017 9380 35069
rect 9432 35017 9448 35069
rect 9500 35017 10232 35069
rect 10284 35017 10300 35069
rect 10352 35017 10368 35069
rect 10420 35017 11152 35069
rect 11204 35017 11220 35069
rect 11272 35017 11288 35069
rect 11340 35017 11592 35069
rect 2877 35004 2914 35017
rect 2970 35004 3006 35017
rect 3062 35014 11592 35017
rect 2992 35002 3006 35004
rect 3062 35002 3109 35014
rect 2387 34994 2872 35002
rect 187 34981 2872 34994
rect 187 34929 2231 34981
rect 2283 34929 2335 34981
rect 2387 34966 2872 34981
rect 2924 34966 2940 35002
rect 2992 34966 3008 35002
rect 3060 34966 3109 35002
rect 2387 34929 2821 34966
rect 2992 34952 3006 34966
rect 3062 34958 3109 34966
rect 3165 34958 3193 35014
rect 3249 34958 3277 35014
rect 3333 34958 3360 35014
rect 3416 34958 3443 35014
rect 3499 34958 3526 35014
rect 3582 34958 3609 35014
rect 3665 34958 3692 35014
rect 3748 34958 3775 35014
rect 3831 35004 3858 35014
rect 3914 35004 3941 35014
rect 3844 34958 3858 35004
rect 3914 34958 3928 35004
rect 3997 34958 4024 35014
rect 4080 34958 4107 35014
rect 4163 34958 4190 35014
rect 4246 34958 4273 35014
rect 4329 34958 4356 35014
rect 4412 34958 4439 35014
rect 4495 34958 4522 35014
rect 4578 34958 4605 35014
rect 4661 34958 4688 35014
rect 4744 35004 4771 35014
rect 4827 35004 4854 35014
rect 4764 34958 4771 35004
rect 3062 34952 3792 34958
rect 3844 34952 3860 34958
rect 3912 34952 3928 34958
rect 3980 34952 4712 34958
rect 4764 34952 4780 34958
rect 4832 34952 4848 35004
rect 4910 34958 4937 35014
rect 4993 34958 5195 35014
rect 5251 34958 5277 35014
rect 5333 34958 5359 35014
rect 5415 34958 5441 35014
rect 5497 34958 5523 35014
rect 5579 34958 5605 35014
rect 5661 35004 5687 35014
rect 5743 35004 5769 35014
rect 5684 34958 5687 35004
rect 4900 34952 5632 34958
rect 5684 34952 5700 34958
rect 5752 34952 5768 35004
rect 5825 34958 5851 35014
rect 5907 34958 5933 35014
rect 5989 34958 6015 35014
rect 6071 34958 6097 35014
rect 6153 34958 6179 35014
rect 6235 34958 6261 35014
rect 6317 34958 6343 35014
rect 6399 34958 6425 35014
rect 6481 34958 6507 35014
rect 6563 35004 6589 35014
rect 6645 35004 6671 35014
rect 6727 35004 6753 35014
rect 6740 34958 6753 35004
rect 6809 35010 11592 35014
rect 6809 34958 6847 35010
rect 5820 34952 6552 34958
rect 6604 34952 6620 34958
rect 6672 34952 6688 34958
rect 6740 34954 6847 34958
rect 6903 34954 6989 35010
rect 7045 35004 11592 35010
rect 7045 34980 7472 35004
rect 7045 34954 7102 34980
rect 6740 34952 7102 34954
rect 2877 34939 2914 34952
rect 2970 34939 3006 34952
rect 3062 34939 7102 34952
rect 187 34916 2821 34929
rect 187 34864 2231 34916
rect 2283 34864 2335 34916
rect 2387 34910 2821 34916
rect 2992 34910 3006 34939
rect 3062 34934 3792 34939
rect 3844 34934 3860 34939
rect 3912 34934 3928 34939
rect 3980 34934 4712 34939
rect 4764 34934 4780 34939
rect 3062 34910 3109 34934
rect 2387 34887 2872 34910
rect 2924 34887 2940 34910
rect 2992 34887 3008 34910
rect 3060 34887 3109 34910
rect 2387 34878 3109 34887
rect 3165 34878 3193 34934
rect 3249 34878 3277 34934
rect 3333 34878 3360 34934
rect 3416 34878 3443 34934
rect 3499 34878 3526 34934
rect 3582 34878 3609 34934
rect 3665 34878 3692 34934
rect 3748 34878 3775 34934
rect 3844 34887 3858 34934
rect 3914 34887 3928 34934
rect 3831 34878 3858 34887
rect 3914 34878 3941 34887
rect 3997 34878 4024 34934
rect 4080 34878 4107 34934
rect 4163 34878 4190 34934
rect 4246 34878 4273 34934
rect 4329 34878 4356 34934
rect 4412 34878 4439 34934
rect 4495 34878 4522 34934
rect 4578 34878 4605 34934
rect 4661 34878 4688 34934
rect 4764 34887 4771 34934
rect 4832 34887 4848 34939
rect 4900 34934 5632 34939
rect 5684 34934 5700 34939
rect 4744 34878 4771 34887
rect 4827 34878 4854 34887
rect 4910 34878 4937 34934
rect 4993 34878 5195 34934
rect 5251 34878 5277 34934
rect 5333 34878 5359 34934
rect 5415 34878 5441 34934
rect 5497 34878 5523 34934
rect 5579 34878 5605 34934
rect 5684 34887 5687 34934
rect 5752 34887 5768 34939
rect 5820 34934 6552 34939
rect 6604 34934 6620 34939
rect 6672 34934 6688 34939
rect 6740 34934 7102 34939
rect 5661 34878 5687 34887
rect 5743 34878 5769 34887
rect 5825 34878 5851 34934
rect 5907 34878 5933 34934
rect 5989 34878 6015 34934
rect 6071 34878 6097 34934
rect 6153 34878 6179 34934
rect 6235 34878 6261 34934
rect 6317 34878 6343 34934
rect 6399 34878 6425 34934
rect 6481 34878 6507 34934
rect 6740 34887 6753 34934
rect 6563 34878 6589 34887
rect 6645 34878 6671 34887
rect 6727 34878 6753 34887
rect 6809 34924 7102 34934
rect 7158 34952 7472 34980
rect 7524 34952 7540 35004
rect 7592 34952 7608 35004
rect 7660 34952 8392 35004
rect 8444 34952 8460 35004
rect 8512 34952 8528 35004
rect 8580 34952 9312 35004
rect 9364 34952 9380 35004
rect 9432 34952 9448 35004
rect 9500 34952 10232 35004
rect 10284 34952 10300 35004
rect 10352 34952 10368 35004
rect 10420 34952 11152 35004
rect 11204 34952 11220 35004
rect 11272 34952 11288 35004
rect 11340 34952 11592 35004
rect 7158 34939 11592 34952
rect 7158 34924 7472 34939
rect 6809 34923 7472 34924
rect 6809 34878 6847 34923
rect 2387 34874 6847 34878
rect 2387 34864 2872 34874
rect 187 34851 2872 34864
rect 187 34799 2231 34851
rect 2283 34799 2335 34851
rect 2387 34822 2872 34851
rect 2924 34822 2940 34874
rect 2992 34851 3008 34874
rect 3060 34854 3792 34874
rect 3844 34854 3860 34874
rect 3912 34854 3928 34874
rect 3980 34854 4712 34874
rect 4764 34854 4780 34874
rect 3060 34822 3109 34854
rect 2387 34809 2963 34822
rect 3019 34809 3109 34822
rect 2387 34799 2872 34809
rect 187 34786 2872 34799
rect 187 34734 2231 34786
rect 2283 34734 2335 34786
rect 2387 34757 2872 34786
rect 2924 34757 2940 34809
rect 3060 34798 3109 34809
rect 3165 34798 3193 34854
rect 3249 34798 3277 34854
rect 3333 34798 3360 34854
rect 3416 34798 3443 34854
rect 3499 34798 3526 34854
rect 3582 34798 3609 34854
rect 3665 34798 3692 34854
rect 3748 34798 3775 34854
rect 3844 34822 3858 34854
rect 3914 34822 3928 34854
rect 3831 34809 3858 34822
rect 3914 34809 3941 34822
rect 3844 34798 3858 34809
rect 3914 34798 3928 34809
rect 3997 34798 4024 34854
rect 4080 34798 4107 34854
rect 4163 34798 4190 34854
rect 4246 34798 4273 34854
rect 4329 34798 4356 34854
rect 4412 34798 4439 34854
rect 4495 34798 4522 34854
rect 4578 34798 4605 34854
rect 4661 34798 4688 34854
rect 4764 34822 4771 34854
rect 4832 34822 4848 34874
rect 4900 34854 5632 34874
rect 5684 34854 5700 34874
rect 4744 34809 4771 34822
rect 4827 34809 4854 34822
rect 4764 34798 4771 34809
rect 2992 34757 3008 34795
rect 3060 34774 3792 34798
rect 3844 34774 3860 34798
rect 3912 34774 3928 34798
rect 3980 34774 4712 34798
rect 4764 34774 4780 34798
rect 3060 34757 3109 34774
rect 2387 34744 3109 34757
rect 2387 34734 2872 34744
rect 187 34721 2872 34734
rect 187 34669 2231 34721
rect 2283 34669 2335 34721
rect 2387 34692 2872 34721
rect 2924 34692 2940 34744
rect 2992 34692 3008 34744
rect 3060 34718 3109 34744
rect 3165 34718 3193 34774
rect 3249 34718 3277 34774
rect 3333 34718 3360 34774
rect 3416 34718 3443 34774
rect 3499 34718 3526 34774
rect 3582 34718 3609 34774
rect 3665 34718 3692 34774
rect 3748 34718 3775 34774
rect 3844 34757 3858 34774
rect 3914 34757 3928 34774
rect 3831 34744 3858 34757
rect 3914 34744 3941 34757
rect 3844 34718 3858 34744
rect 3914 34718 3928 34744
rect 3997 34718 4024 34774
rect 4080 34718 4107 34774
rect 4163 34718 4190 34774
rect 4246 34718 4273 34774
rect 4329 34718 4356 34774
rect 4412 34718 4439 34774
rect 4495 34718 4522 34774
rect 4578 34718 4605 34774
rect 4661 34718 4688 34774
rect 4764 34757 4771 34774
rect 4832 34757 4848 34809
rect 4910 34798 4937 34854
rect 4993 34798 5195 34854
rect 5251 34798 5277 34854
rect 5333 34798 5359 34854
rect 5415 34798 5441 34854
rect 5497 34798 5523 34854
rect 5579 34798 5605 34854
rect 5684 34822 5687 34854
rect 5752 34822 5768 34874
rect 5820 34854 6552 34874
rect 6604 34854 6620 34874
rect 6672 34854 6688 34874
rect 6740 34867 6847 34874
rect 6903 34867 6989 34923
rect 7045 34887 7472 34923
rect 7524 34887 7540 34939
rect 7592 34887 7608 34939
rect 7660 34887 8392 34939
rect 8444 34887 8460 34939
rect 8512 34887 8528 34939
rect 8580 34887 9312 34939
rect 9364 34887 9380 34939
rect 9432 34887 9448 34939
rect 9500 34887 10232 34939
rect 10284 34887 10300 34939
rect 10352 34887 10368 34939
rect 10420 34887 11152 34939
rect 11204 34887 11220 34939
rect 11272 34887 11288 34939
rect 11340 34887 11592 34939
rect 7045 34874 11592 34887
rect 7045 34867 7472 34874
rect 6740 34854 7472 34867
rect 5661 34809 5687 34822
rect 5743 34809 5769 34822
rect 5684 34798 5687 34809
rect 4900 34774 5632 34798
rect 5684 34774 5700 34798
rect 4744 34744 4771 34757
rect 4827 34744 4854 34757
rect 4764 34718 4771 34744
rect 3060 34694 3792 34718
rect 3844 34694 3860 34718
rect 3912 34694 3928 34718
rect 3980 34694 4712 34718
rect 4764 34694 4780 34718
rect 3060 34692 3109 34694
rect 2387 34679 3109 34692
rect 2387 34669 2872 34679
rect 187 34656 2872 34669
rect 187 34604 2231 34656
rect 2283 34604 2335 34656
rect 2387 34627 2872 34656
rect 2924 34627 2940 34679
rect 2992 34627 3008 34679
rect 3060 34638 3109 34679
rect 3165 34638 3193 34694
rect 3249 34638 3277 34694
rect 3333 34638 3360 34694
rect 3416 34638 3443 34694
rect 3499 34638 3526 34694
rect 3582 34638 3609 34694
rect 3665 34638 3692 34694
rect 3748 34638 3775 34694
rect 3844 34692 3858 34694
rect 3914 34692 3928 34694
rect 3831 34679 3858 34692
rect 3914 34679 3941 34692
rect 3844 34638 3858 34679
rect 3914 34638 3928 34679
rect 3997 34638 4024 34694
rect 4080 34638 4107 34694
rect 4163 34638 4190 34694
rect 4246 34638 4273 34694
rect 4329 34638 4356 34694
rect 4412 34638 4439 34694
rect 4495 34638 4522 34694
rect 4578 34638 4605 34694
rect 4661 34638 4688 34694
rect 4764 34692 4771 34694
rect 4832 34692 4848 34744
rect 4910 34718 4937 34774
rect 4993 34718 5195 34774
rect 5251 34718 5277 34774
rect 5333 34718 5359 34774
rect 5415 34718 5441 34774
rect 5497 34718 5523 34774
rect 5579 34718 5605 34774
rect 5684 34757 5687 34774
rect 5752 34757 5768 34809
rect 5825 34798 5851 34854
rect 5907 34798 5933 34854
rect 5989 34798 6015 34854
rect 6071 34798 6097 34854
rect 6153 34798 6179 34854
rect 6235 34798 6261 34854
rect 6317 34798 6343 34854
rect 6399 34798 6425 34854
rect 6481 34798 6507 34854
rect 6740 34822 6753 34854
rect 6563 34809 6589 34822
rect 6645 34809 6671 34822
rect 6727 34809 6753 34822
rect 6740 34798 6753 34809
rect 6809 34835 7472 34854
rect 6809 34798 6847 34835
rect 5820 34774 6552 34798
rect 6604 34774 6620 34798
rect 6672 34774 6688 34798
rect 6740 34779 6847 34798
rect 6903 34779 6989 34835
rect 7045 34822 7472 34835
rect 7524 34822 7540 34874
rect 7592 34822 7608 34874
rect 7660 34822 8392 34874
rect 8444 34822 8460 34874
rect 8512 34822 8528 34874
rect 8580 34822 9312 34874
rect 9364 34822 9380 34874
rect 9432 34822 9448 34874
rect 9500 34822 10232 34874
rect 10284 34822 10300 34874
rect 10352 34822 10368 34874
rect 10420 34822 11152 34874
rect 11204 34822 11220 34874
rect 11272 34822 11288 34874
rect 11340 34822 11592 34874
rect 7045 34809 11592 34822
rect 7045 34779 7472 34809
rect 6740 34774 7472 34779
rect 5661 34744 5687 34757
rect 5743 34744 5769 34757
rect 5684 34718 5687 34744
rect 4900 34694 5632 34718
rect 5684 34694 5700 34718
rect 4744 34679 4771 34692
rect 4827 34679 4854 34692
rect 4764 34638 4771 34679
rect 3060 34627 3792 34638
rect 3844 34627 3860 34638
rect 3912 34627 3928 34638
rect 3980 34627 4712 34638
rect 4764 34627 4780 34638
rect 4832 34627 4848 34679
rect 4910 34638 4937 34694
rect 4993 34638 5195 34694
rect 5251 34638 5277 34694
rect 5333 34638 5359 34694
rect 5415 34638 5441 34694
rect 5497 34638 5523 34694
rect 5579 34638 5605 34694
rect 5684 34692 5687 34694
rect 5752 34692 5768 34744
rect 5825 34718 5851 34774
rect 5907 34718 5933 34774
rect 5989 34718 6015 34774
rect 6071 34718 6097 34774
rect 6153 34718 6179 34774
rect 6235 34718 6261 34774
rect 6317 34718 6343 34774
rect 6399 34718 6425 34774
rect 6481 34718 6507 34774
rect 6740 34757 6753 34774
rect 6563 34744 6589 34757
rect 6645 34744 6671 34757
rect 6727 34744 6753 34757
rect 6740 34718 6753 34744
rect 6809 34757 7472 34774
rect 7524 34757 7540 34809
rect 7592 34757 7608 34809
rect 7660 34757 8392 34809
rect 8444 34757 8460 34809
rect 8512 34757 8528 34809
rect 8580 34757 9312 34809
rect 9364 34757 9380 34809
rect 9432 34757 9448 34809
rect 9500 34757 10232 34809
rect 10284 34757 10300 34809
rect 10352 34757 10368 34809
rect 10420 34757 11152 34809
rect 11204 34757 11220 34809
rect 11272 34757 11288 34809
rect 11340 34757 11592 34809
rect 6809 34744 11592 34757
rect 6809 34718 7472 34744
rect 5820 34694 6552 34718
rect 6604 34694 6620 34718
rect 6672 34694 6688 34718
rect 6740 34695 7472 34718
rect 6740 34694 6847 34695
rect 5661 34679 5687 34692
rect 5743 34679 5769 34692
rect 5684 34638 5687 34679
rect 4900 34627 5632 34638
rect 5684 34627 5700 34638
rect 5752 34627 5768 34679
rect 5825 34638 5851 34694
rect 5907 34638 5933 34694
rect 5989 34638 6015 34694
rect 6071 34638 6097 34694
rect 6153 34638 6179 34694
rect 6235 34638 6261 34694
rect 6317 34638 6343 34694
rect 6399 34638 6425 34694
rect 6481 34638 6507 34694
rect 6740 34692 6753 34694
rect 6563 34679 6589 34692
rect 6645 34679 6671 34692
rect 6727 34679 6753 34692
rect 6740 34638 6753 34679
rect 6809 34639 6847 34694
rect 6903 34692 7472 34695
rect 7524 34692 7540 34744
rect 7592 34692 7608 34744
rect 7660 34692 8392 34744
rect 8444 34692 8460 34744
rect 8512 34692 8528 34744
rect 8580 34692 9312 34744
rect 9364 34692 9380 34744
rect 9432 34692 9448 34744
rect 9500 34692 10232 34744
rect 10284 34692 10300 34744
rect 10352 34692 10368 34744
rect 10420 34692 11152 34744
rect 11204 34692 11220 34744
rect 11272 34692 11288 34744
rect 11340 34692 11592 34744
rect 6903 34679 11592 34692
rect 6903 34639 7472 34679
rect 6809 34638 7472 34639
rect 5820 34627 6552 34638
rect 6604 34627 6620 34638
rect 6672 34627 6688 34638
rect 6740 34627 7472 34638
rect 7524 34627 7540 34679
rect 7592 34627 7608 34679
rect 7660 34627 8392 34679
rect 8444 34627 8460 34679
rect 8512 34627 8528 34679
rect 8580 34627 9312 34679
rect 9364 34627 9380 34679
rect 9432 34627 9448 34679
rect 9500 34627 10232 34679
rect 10284 34627 10300 34679
rect 10352 34627 10368 34679
rect 10420 34627 11152 34679
rect 11204 34627 11220 34679
rect 11272 34627 11288 34679
rect 11340 34627 11592 34679
rect 2387 34614 11592 34627
rect 2387 34604 2872 34614
rect 187 34591 2872 34604
rect 187 34539 2231 34591
rect 2283 34539 2335 34591
rect 2387 34562 2872 34591
rect 2924 34562 2940 34614
rect 2992 34562 3008 34614
rect 3060 34562 3109 34614
rect 2387 34558 3109 34562
rect 3165 34558 3193 34614
rect 3249 34558 3277 34614
rect 3333 34558 3360 34614
rect 3416 34558 3443 34614
rect 3499 34558 3526 34614
rect 3582 34558 3609 34614
rect 3665 34558 3692 34614
rect 3748 34558 3775 34614
rect 3844 34562 3858 34614
rect 3914 34562 3928 34614
rect 3831 34558 3858 34562
rect 3914 34558 3941 34562
rect 3997 34558 4024 34614
rect 4080 34558 4107 34614
rect 4163 34558 4190 34614
rect 4246 34558 4273 34614
rect 4329 34558 4356 34614
rect 4412 34558 4439 34614
rect 4495 34558 4522 34614
rect 4578 34558 4605 34614
rect 4661 34558 4688 34614
rect 4764 34562 4771 34614
rect 4832 34562 4848 34614
rect 4744 34558 4771 34562
rect 4827 34558 4854 34562
rect 4910 34558 4937 34614
rect 4993 34558 5195 34614
rect 5251 34558 5277 34614
rect 5333 34558 5359 34614
rect 5415 34558 5441 34614
rect 5497 34558 5523 34614
rect 5579 34558 5605 34614
rect 5684 34562 5687 34614
rect 5752 34562 5768 34614
rect 5661 34558 5687 34562
rect 5743 34558 5769 34562
rect 5825 34558 5851 34614
rect 5907 34558 5933 34614
rect 5989 34558 6015 34614
rect 6071 34558 6097 34614
rect 6153 34558 6179 34614
rect 6235 34558 6261 34614
rect 6317 34558 6343 34614
rect 6399 34558 6425 34614
rect 6481 34558 6507 34614
rect 6740 34562 6753 34614
rect 6563 34558 6589 34562
rect 6645 34558 6671 34562
rect 6727 34558 6753 34562
rect 6809 34562 7472 34614
rect 7524 34562 7540 34614
rect 7592 34562 7608 34614
rect 7660 34562 8392 34614
rect 8444 34562 8460 34614
rect 8512 34562 8528 34614
rect 8580 34562 9312 34614
rect 9364 34562 9380 34614
rect 9432 34562 9448 34614
rect 9500 34562 10232 34614
rect 10284 34562 10300 34614
rect 10352 34562 10368 34614
rect 10420 34562 11152 34614
rect 11204 34562 11220 34614
rect 11272 34562 11288 34614
rect 11340 34562 11592 34614
rect 6809 34558 11592 34562
rect 2387 34556 11592 34558
tri 11838 34556 12222 34940 se
rect 12222 34556 14858 37059
rect 2387 34539 3342 34556
rect 187 34526 3342 34539
rect 187 34474 2231 34526
rect 2283 34474 2335 34526
rect 2387 34474 3342 34526
rect 187 34461 3342 34474
rect 187 34409 2231 34461
rect 2283 34409 2335 34461
rect 2387 34409 3342 34461
rect 187 34396 3342 34409
rect 187 34344 2231 34396
rect 2283 34344 2335 34396
rect 2387 34362 3342 34396
tri 3342 34362 3536 34556 nw
rect 2387 34344 2824 34362
rect 187 34331 2824 34344
rect 187 34279 2231 34331
rect 2283 34279 2335 34331
rect 2387 34279 2824 34331
rect 187 34266 2824 34279
rect 187 34214 2231 34266
rect 2283 34214 2335 34266
rect 2387 34214 2824 34266
rect 187 31774 2824 34214
tri 2824 33844 3342 34362 nw
tri 11513 34231 11838 34556 se
rect 11838 34231 14858 34556
rect 3361 34229 14858 34231
rect 3361 34225 8580 34229
rect 3413 34173 3439 34225
rect 3491 34173 4281 34225
rect 4333 34173 4359 34225
rect 4411 34173 5201 34225
rect 5253 34173 5279 34225
rect 5331 34173 6121 34225
rect 6173 34173 6199 34225
rect 6251 34173 7041 34225
rect 7093 34173 7119 34225
rect 7171 34173 7961 34225
rect 8013 34173 8039 34225
rect 8091 34173 8580 34225
rect 8636 34173 8661 34229
rect 8717 34173 8742 34229
rect 8798 34173 8823 34229
rect 8879 34225 8904 34229
rect 8960 34225 8985 34229
rect 8879 34173 8881 34225
rect 9041 34173 9066 34229
rect 3361 34161 9066 34173
rect 3413 34109 3439 34161
rect 3491 34109 4281 34161
rect 4333 34109 4359 34161
rect 4411 34109 5201 34161
rect 5253 34109 5279 34161
rect 5331 34109 6121 34161
rect 6173 34109 6199 34161
rect 6251 34109 7041 34161
rect 7093 34109 7119 34161
rect 7171 34109 7961 34161
rect 8013 34109 8039 34161
rect 8091 34149 8881 34161
rect 8933 34149 8959 34161
rect 9011 34149 9066 34161
rect 8091 34109 8580 34149
rect 3361 34097 8580 34109
rect 3413 34045 3439 34097
rect 3491 34045 4281 34097
rect 4333 34045 4359 34097
rect 4411 34045 5201 34097
rect 5253 34045 5279 34097
rect 5331 34045 6121 34097
rect 6173 34045 6199 34097
rect 6251 34045 7041 34097
rect 7093 34045 7119 34097
rect 7171 34045 7961 34097
rect 8013 34045 8039 34097
rect 8091 34093 8580 34097
rect 8636 34093 8661 34149
rect 8717 34093 8742 34149
rect 8798 34093 8823 34149
rect 8879 34109 8881 34149
rect 8879 34097 8904 34109
rect 8960 34097 8985 34109
rect 8879 34093 8881 34097
rect 9041 34093 9066 34149
rect 8091 34069 8881 34093
rect 8933 34069 8959 34093
rect 9011 34069 9066 34093
rect 8091 34045 8580 34069
rect 3361 34033 8580 34045
rect 3413 33981 3439 34033
rect 3491 33981 4281 34033
rect 4333 33981 4359 34033
rect 4411 33981 5201 34033
rect 5253 33981 5279 34033
rect 5331 33981 6121 34033
rect 6173 33981 6199 34033
rect 6251 33981 7041 34033
rect 7093 33981 7119 34033
rect 7171 33981 7961 34033
rect 8013 33981 8039 34033
rect 8091 34013 8580 34033
rect 8636 34013 8661 34069
rect 8717 34013 8742 34069
rect 8798 34013 8823 34069
rect 8879 34045 8881 34069
rect 8879 34033 8904 34045
rect 8960 34033 8985 34045
rect 8879 34013 8881 34033
rect 9041 34013 9066 34069
rect 8091 33989 8881 34013
rect 8933 33989 8959 34013
rect 9011 33989 9066 34013
rect 8091 33981 8580 33989
rect 3361 33969 8580 33981
rect 3413 33917 3439 33969
rect 3491 33917 4281 33969
rect 4333 33917 4359 33969
rect 4411 33917 5201 33969
rect 5253 33917 5279 33969
rect 5331 33917 6121 33969
rect 6173 33917 6199 33969
rect 6251 33917 7041 33969
rect 7093 33917 7119 33969
rect 7171 33917 7961 33969
rect 8013 33917 8039 33969
rect 8091 33933 8580 33969
rect 8636 33933 8661 33989
rect 8717 33933 8742 33989
rect 8798 33933 8823 33989
rect 8879 33981 8881 33989
rect 8879 33969 8904 33981
rect 8960 33969 8985 33981
rect 8879 33933 8881 33969
rect 9041 33933 9066 33989
rect 8091 33917 8881 33933
rect 8933 33917 8959 33933
rect 9011 33917 9066 33933
rect 3361 33909 9066 33917
rect 3361 33905 8580 33909
rect 3413 33853 3439 33905
rect 3491 33853 4281 33905
rect 4333 33853 4359 33905
rect 4411 33853 5201 33905
rect 5253 33853 5279 33905
rect 5331 33853 6121 33905
rect 6173 33853 6199 33905
rect 6251 33853 7041 33905
rect 7093 33853 7119 33905
rect 7171 33853 7961 33905
rect 8013 33853 8039 33905
rect 8091 33853 8580 33905
rect 8636 33853 8661 33909
rect 8717 33853 8742 33909
rect 8798 33853 8823 33909
rect 8879 33905 8904 33909
rect 8960 33905 8985 33909
rect 8879 33853 8881 33905
rect 9041 33853 9066 33909
rect 3361 33841 9066 33853
rect 3413 33789 3439 33841
rect 3491 33789 4281 33841
rect 4333 33789 4359 33841
rect 4411 33789 5201 33841
rect 5253 33789 5279 33841
rect 5331 33789 6121 33841
rect 6173 33789 6199 33841
rect 6251 33789 7041 33841
rect 7093 33789 7119 33841
rect 7171 33789 7961 33841
rect 8013 33789 8039 33841
rect 8091 33829 8881 33841
rect 8933 33829 8959 33841
rect 9011 33829 9066 33841
rect 8091 33789 8580 33829
rect 3361 33777 8580 33789
rect 3413 33725 3439 33777
rect 3491 33725 4281 33777
rect 4333 33725 4359 33777
rect 4411 33725 5201 33777
rect 5253 33725 5279 33777
rect 5331 33725 6121 33777
rect 6173 33725 6199 33777
rect 6251 33725 7041 33777
rect 7093 33725 7119 33777
rect 7171 33725 7961 33777
rect 8013 33725 8039 33777
rect 8091 33773 8580 33777
rect 8636 33773 8661 33829
rect 8717 33773 8742 33829
rect 8798 33773 8823 33829
rect 8879 33789 8881 33829
rect 8879 33777 8904 33789
rect 8960 33777 8985 33789
rect 8879 33773 8881 33777
rect 9041 33773 9066 33829
rect 8091 33749 8881 33773
rect 8933 33749 8959 33773
rect 9011 33749 9066 33773
rect 8091 33725 8580 33749
rect 3361 33713 8580 33725
rect 3413 33661 3439 33713
rect 3491 33661 4281 33713
rect 4333 33661 4359 33713
rect 4411 33661 5201 33713
rect 5253 33661 5279 33713
rect 5331 33661 6121 33713
rect 6173 33661 6199 33713
rect 6251 33661 7041 33713
rect 7093 33661 7119 33713
rect 7171 33661 7961 33713
rect 8013 33661 8039 33713
rect 8091 33693 8580 33713
rect 8636 33693 8661 33749
rect 8717 33693 8742 33749
rect 8798 33693 8823 33749
rect 8879 33725 8881 33749
rect 8879 33713 8904 33725
rect 8960 33713 8985 33725
rect 8879 33693 8881 33713
rect 9041 33693 9066 33749
rect 8091 33669 8881 33693
rect 8933 33669 8959 33693
rect 9011 33669 9066 33693
rect 8091 33661 8580 33669
rect 3361 33649 8580 33661
rect 3413 33597 3439 33649
rect 3491 33597 4281 33649
rect 4333 33597 4359 33649
rect 4411 33597 5201 33649
rect 5253 33597 5279 33649
rect 5331 33597 6121 33649
rect 6173 33597 6199 33649
rect 6251 33597 7041 33649
rect 7093 33597 7119 33649
rect 7171 33597 7961 33649
rect 8013 33597 8039 33649
rect 8091 33613 8580 33649
rect 8636 33613 8661 33669
rect 8717 33613 8742 33669
rect 8798 33613 8823 33669
rect 8879 33661 8881 33669
rect 8879 33649 8904 33661
rect 8960 33649 8985 33661
rect 8879 33613 8881 33649
rect 9041 33613 9066 33669
rect 8091 33597 8881 33613
rect 8933 33597 8959 33613
rect 9011 33597 9066 33613
rect 3361 33589 9066 33597
rect 3361 33585 8580 33589
rect 3413 33533 3439 33585
rect 3491 33533 4281 33585
rect 4333 33533 4359 33585
rect 4411 33533 5201 33585
rect 5253 33533 5279 33585
rect 5331 33533 6121 33585
rect 6173 33533 6199 33585
rect 6251 33533 7041 33585
rect 7093 33533 7119 33585
rect 7171 33533 7961 33585
rect 8013 33533 8039 33585
rect 8091 33533 8580 33585
rect 8636 33533 8661 33589
rect 8717 33533 8742 33589
rect 8798 33533 8823 33589
rect 8879 33585 8904 33589
rect 8960 33585 8985 33589
rect 8879 33533 8881 33585
rect 9041 33533 9066 33589
rect 3361 33521 9066 33533
rect 3413 33469 3439 33521
rect 3491 33469 4281 33521
rect 4333 33469 4359 33521
rect 4411 33469 5201 33521
rect 5253 33469 5279 33521
rect 5331 33469 6121 33521
rect 6173 33469 6199 33521
rect 6251 33469 7041 33521
rect 7093 33469 7119 33521
rect 7171 33469 7961 33521
rect 8013 33469 8039 33521
rect 8091 33509 8881 33521
rect 8933 33509 8959 33521
rect 9011 33509 9066 33521
rect 8091 33469 8580 33509
rect 3361 33457 8580 33469
rect 3413 33405 3439 33457
rect 3491 33405 4281 33457
rect 4333 33405 4359 33457
rect 4411 33405 5201 33457
rect 5253 33405 5279 33457
rect 5331 33405 6121 33457
rect 6173 33405 6199 33457
rect 6251 33405 7041 33457
rect 7093 33405 7119 33457
rect 7171 33405 7961 33457
rect 8013 33405 8039 33457
rect 8091 33453 8580 33457
rect 8636 33453 8661 33509
rect 8717 33453 8742 33509
rect 8798 33453 8823 33509
rect 8879 33469 8881 33509
rect 8879 33457 8904 33469
rect 8960 33457 8985 33469
rect 8879 33453 8881 33457
rect 9041 33453 9066 33509
rect 8091 33429 8881 33453
rect 8933 33429 8959 33453
rect 9011 33429 9066 33453
rect 8091 33405 8580 33429
rect 3361 33393 8580 33405
rect 3413 33341 3439 33393
rect 3491 33341 4281 33393
rect 4333 33341 4359 33393
rect 4411 33341 5201 33393
rect 5253 33341 5279 33393
rect 5331 33341 6121 33393
rect 6173 33341 6199 33393
rect 6251 33341 7041 33393
rect 7093 33341 7119 33393
rect 7171 33341 7961 33393
rect 8013 33341 8039 33393
rect 8091 33373 8580 33393
rect 8636 33373 8661 33429
rect 8717 33373 8742 33429
rect 8798 33373 8823 33429
rect 8879 33405 8881 33429
rect 8879 33393 8904 33405
rect 8960 33393 8985 33405
rect 8879 33373 8881 33393
rect 9041 33373 9066 33429
rect 8091 33349 8881 33373
rect 8933 33349 8959 33373
rect 9011 33349 9066 33373
rect 8091 33341 8580 33349
rect 3361 33329 8580 33341
rect 3413 33277 3439 33329
rect 3491 33277 4281 33329
rect 4333 33277 4359 33329
rect 4411 33277 5201 33329
rect 5253 33277 5279 33329
rect 5331 33277 6121 33329
rect 6173 33277 6199 33329
rect 6251 33277 7041 33329
rect 7093 33277 7119 33329
rect 7171 33277 7961 33329
rect 8013 33277 8039 33329
rect 8091 33293 8580 33329
rect 8636 33293 8661 33349
rect 8717 33293 8742 33349
rect 8798 33293 8823 33349
rect 8879 33341 8881 33349
rect 8879 33329 8904 33341
rect 8960 33329 8985 33341
rect 8879 33293 8881 33329
rect 9041 33293 9066 33349
rect 8091 33277 8881 33293
rect 8933 33277 8959 33293
rect 9011 33277 9066 33293
rect 3361 33269 9066 33277
rect 3361 33264 8580 33269
rect 3413 33212 3439 33264
rect 3491 33212 4281 33264
rect 4333 33212 4359 33264
rect 4411 33212 5201 33264
rect 5253 33212 5279 33264
rect 5331 33212 6121 33264
rect 6173 33212 6199 33264
rect 6251 33212 7041 33264
rect 7093 33212 7119 33264
rect 7171 33212 7961 33264
rect 8013 33212 8039 33264
rect 8091 33213 8580 33264
rect 8636 33213 8661 33269
rect 8717 33213 8742 33269
rect 8798 33213 8823 33269
rect 8879 33264 8904 33269
rect 8960 33264 8985 33269
rect 8879 33213 8881 33264
rect 9041 33213 9066 33269
rect 8091 33212 8881 33213
rect 8933 33212 8959 33213
rect 9011 33212 9066 33213
rect 3361 33199 9066 33212
rect 3413 33147 3439 33199
rect 3491 33147 4281 33199
rect 4333 33147 4359 33199
rect 4411 33147 5201 33199
rect 5253 33147 5279 33199
rect 5331 33147 6121 33199
rect 6173 33147 6199 33199
rect 6251 33147 7041 33199
rect 7093 33147 7119 33199
rect 7171 33147 7961 33199
rect 8013 33147 8039 33199
rect 8091 33189 8881 33199
rect 8933 33189 8959 33199
rect 9011 33189 9066 33199
rect 8091 33147 8580 33189
rect 3361 33134 8580 33147
rect 3413 33082 3439 33134
rect 3491 33082 4281 33134
rect 4333 33082 4359 33134
rect 4411 33082 5201 33134
rect 5253 33082 5279 33134
rect 5331 33082 6121 33134
rect 6173 33082 6199 33134
rect 6251 33082 7041 33134
rect 7093 33082 7119 33134
rect 7171 33082 7961 33134
rect 8013 33082 8039 33134
rect 8091 33133 8580 33134
rect 8636 33133 8661 33189
rect 8717 33133 8742 33189
rect 8798 33133 8823 33189
rect 8879 33147 8881 33189
rect 8879 33134 8904 33147
rect 8960 33134 8985 33147
rect 8879 33133 8881 33134
rect 9041 33133 9066 33189
rect 8091 33109 8881 33133
rect 8933 33109 8959 33133
rect 9011 33109 9066 33133
rect 8091 33082 8580 33109
rect 3361 33069 8580 33082
rect 3413 33017 3439 33069
rect 3491 33017 4281 33069
rect 4333 33017 4359 33069
rect 4411 33017 5201 33069
rect 5253 33017 5279 33069
rect 5331 33017 6121 33069
rect 6173 33017 6199 33069
rect 6251 33017 7041 33069
rect 7093 33017 7119 33069
rect 7171 33017 7961 33069
rect 8013 33017 8039 33069
rect 8091 33053 8580 33069
rect 8636 33053 8661 33109
rect 8717 33053 8742 33109
rect 8798 33053 8823 33109
rect 8879 33082 8881 33109
rect 8879 33069 8904 33082
rect 8960 33069 8985 33082
rect 8879 33053 8881 33069
rect 9041 33053 9066 33109
rect 8091 33029 8881 33053
rect 8933 33029 8959 33053
rect 9011 33029 9066 33053
rect 8091 33017 8580 33029
rect 3361 33004 8580 33017
rect 3413 32952 3439 33004
rect 3491 32952 4281 33004
rect 4333 32952 4359 33004
rect 4411 32952 5201 33004
rect 5253 32952 5279 33004
rect 5331 32952 6121 33004
rect 6173 32952 6199 33004
rect 6251 32952 7041 33004
rect 7093 32952 7119 33004
rect 7171 32952 7961 33004
rect 8013 32952 8039 33004
rect 8091 32973 8580 33004
rect 8636 32973 8661 33029
rect 8717 32973 8742 33029
rect 8798 32973 8823 33029
rect 8879 33017 8881 33029
rect 8879 33004 8904 33017
rect 8960 33004 8985 33017
rect 8879 32973 8881 33004
rect 9041 32973 9066 33029
rect 8091 32952 8881 32973
rect 8933 32952 8959 32973
rect 9011 32952 9066 32973
rect 3361 32949 9066 32952
rect 3361 32939 8580 32949
rect 3413 32887 3439 32939
rect 3491 32887 4281 32939
rect 4333 32887 4359 32939
rect 4411 32887 5201 32939
rect 5253 32887 5279 32939
rect 5331 32887 6121 32939
rect 6173 32887 6199 32939
rect 6251 32887 7041 32939
rect 7093 32887 7119 32939
rect 7171 32887 7961 32939
rect 8013 32887 8039 32939
rect 8091 32893 8580 32939
rect 8636 32893 8661 32949
rect 8717 32893 8742 32949
rect 8798 32893 8823 32949
rect 8879 32939 8904 32949
rect 8960 32939 8985 32949
rect 8879 32893 8881 32939
rect 9041 32893 9066 32949
rect 8091 32887 8881 32893
rect 8933 32887 8959 32893
rect 9011 32887 9066 32893
rect 3361 32874 9066 32887
rect 3413 32822 3439 32874
rect 3491 32822 4281 32874
rect 4333 32822 4359 32874
rect 4411 32822 5201 32874
rect 5253 32822 5279 32874
rect 5331 32822 6121 32874
rect 6173 32822 6199 32874
rect 6251 32822 7041 32874
rect 7093 32822 7119 32874
rect 7171 32822 7961 32874
rect 8013 32822 8039 32874
rect 8091 32869 8881 32874
rect 8933 32869 8959 32874
rect 9011 32869 9066 32874
rect 8091 32822 8580 32869
rect 3361 32813 8580 32822
rect 8636 32813 8661 32869
rect 8717 32813 8742 32869
rect 8798 32813 8823 32869
rect 8879 32822 8881 32869
rect 8879 32813 8904 32822
rect 8960 32813 8985 32822
rect 9041 32813 9066 32869
rect 3361 32809 9066 32813
rect 3413 32757 3439 32809
rect 3491 32757 4281 32809
rect 4333 32757 4359 32809
rect 4411 32757 5201 32809
rect 5253 32757 5279 32809
rect 5331 32757 6121 32809
rect 6173 32757 6199 32809
rect 6251 32757 7041 32809
rect 7093 32757 7119 32809
rect 7171 32757 7961 32809
rect 8013 32757 8039 32809
rect 8091 32789 8881 32809
rect 8933 32789 8959 32809
rect 9011 32789 9066 32809
rect 8091 32757 8580 32789
rect 3361 32744 8580 32757
rect 3413 32692 3439 32744
rect 3491 32692 4281 32744
rect 4333 32692 4359 32744
rect 4411 32692 5201 32744
rect 5253 32692 5279 32744
rect 5331 32692 6121 32744
rect 6173 32692 6199 32744
rect 6251 32692 7041 32744
rect 7093 32692 7119 32744
rect 7171 32692 7961 32744
rect 8013 32692 8039 32744
rect 8091 32733 8580 32744
rect 8636 32733 8661 32789
rect 8717 32733 8742 32789
rect 8798 32733 8823 32789
rect 8879 32757 8881 32789
rect 8879 32744 8904 32757
rect 8960 32744 8985 32757
rect 8879 32733 8881 32744
rect 9041 32733 9066 32789
rect 8091 32709 8881 32733
rect 8933 32709 8959 32733
rect 9011 32709 9066 32733
rect 8091 32692 8580 32709
rect 3361 32679 8580 32692
rect 3413 32627 3439 32679
rect 3491 32627 4281 32679
rect 4333 32627 4359 32679
rect 4411 32627 5201 32679
rect 5253 32627 5279 32679
rect 5331 32627 6121 32679
rect 6173 32627 6199 32679
rect 6251 32627 7041 32679
rect 7093 32627 7119 32679
rect 7171 32627 7961 32679
rect 8013 32627 8039 32679
rect 8091 32653 8580 32679
rect 8636 32653 8661 32709
rect 8717 32653 8742 32709
rect 8798 32653 8823 32709
rect 8879 32692 8881 32709
rect 8879 32679 8904 32692
rect 8960 32679 8985 32692
rect 8879 32653 8881 32679
rect 9041 32653 9066 32709
rect 8091 32629 8881 32653
rect 8933 32629 8959 32653
rect 9011 32629 9066 32653
rect 8091 32627 8580 32629
rect 3361 32614 8580 32627
rect 3413 32562 3439 32614
rect 3491 32562 4281 32614
rect 4333 32562 4359 32614
rect 4411 32562 5201 32614
rect 5253 32562 5279 32614
rect 5331 32562 6121 32614
rect 6173 32562 6199 32614
rect 6251 32562 7041 32614
rect 7093 32562 7119 32614
rect 7171 32562 7961 32614
rect 8013 32562 8039 32614
rect 8091 32573 8580 32614
rect 8636 32573 8661 32629
rect 8717 32573 8742 32629
rect 8798 32573 8823 32629
rect 8879 32627 8881 32629
rect 8879 32614 8904 32627
rect 8960 32614 8985 32627
rect 8879 32573 8881 32614
rect 9041 32573 9066 32629
rect 8091 32562 8881 32573
rect 8933 32562 8959 32573
rect 9011 32562 9066 32573
rect 3361 32549 9066 32562
rect 3413 32497 3439 32549
rect 3491 32497 4281 32549
rect 4333 32497 4359 32549
rect 4411 32497 5201 32549
rect 5253 32497 5279 32549
rect 5331 32497 6121 32549
rect 6173 32497 6199 32549
rect 6251 32497 7041 32549
rect 7093 32497 7119 32549
rect 7171 32497 7961 32549
rect 8013 32497 8039 32549
rect 8091 32497 8580 32549
rect 3361 32493 8580 32497
rect 8636 32493 8661 32549
rect 8717 32493 8742 32549
rect 8798 32493 8823 32549
rect 8879 32497 8881 32549
rect 8879 32493 8904 32497
rect 8960 32493 8985 32497
rect 9041 32493 9066 32549
rect 9762 34225 10666 34229
rect 10722 34225 10747 34229
rect 10803 34225 10828 34229
rect 9762 34173 9801 34225
rect 9853 34173 9879 34225
rect 9931 34173 10666 34225
rect 10884 34173 10909 34229
rect 10965 34173 10990 34229
rect 11046 34173 11071 34229
rect 11127 34173 11152 34229
rect 11848 34225 14858 34229
rect 11848 34173 12561 34225
rect 12613 34173 12639 34225
rect 12691 34173 14858 34225
rect 9762 34161 11152 34173
rect 11848 34161 14858 34173
rect 9762 34109 9801 34161
rect 9853 34109 9879 34161
rect 9931 34149 10721 34161
rect 10773 34149 10799 34161
rect 10851 34149 11152 34161
rect 9931 34109 10666 34149
rect 9762 34097 10666 34109
rect 10722 34097 10747 34109
rect 10803 34097 10828 34109
rect 9762 34045 9801 34097
rect 9853 34045 9879 34097
rect 9931 34093 10666 34097
rect 10884 34093 10909 34149
rect 10965 34093 10990 34149
rect 11046 34093 11071 34149
rect 11127 34093 11152 34149
rect 11848 34109 12561 34161
rect 12613 34109 12639 34161
rect 12691 34109 14858 34161
rect 11848 34097 14858 34109
rect 9931 34069 10721 34093
rect 10773 34069 10799 34093
rect 10851 34069 11152 34093
rect 9931 34045 10666 34069
rect 9762 34033 10666 34045
rect 10722 34033 10747 34045
rect 10803 34033 10828 34045
rect 9762 33981 9801 34033
rect 9853 33981 9879 34033
rect 9931 34013 10666 34033
rect 10884 34013 10909 34069
rect 10965 34013 10990 34069
rect 11046 34013 11071 34069
rect 11127 34013 11152 34069
rect 11848 34045 12561 34097
rect 12613 34045 12639 34097
rect 12691 34045 14858 34097
rect 11848 34033 14858 34045
rect 9931 33989 10721 34013
rect 10773 33989 10799 34013
rect 10851 33989 11152 34013
rect 9931 33981 10666 33989
rect 9762 33969 10666 33981
rect 10722 33969 10747 33981
rect 10803 33969 10828 33981
rect 9762 33917 9801 33969
rect 9853 33917 9879 33969
rect 9931 33933 10666 33969
rect 10884 33933 10909 33989
rect 10965 33933 10990 33989
rect 11046 33933 11071 33989
rect 11127 33933 11152 33989
rect 11848 33981 12561 34033
rect 12613 33981 12639 34033
rect 12691 33981 14858 34033
rect 11848 33969 14858 33981
rect 9931 33917 10721 33933
rect 10773 33917 10799 33933
rect 10851 33917 11152 33933
rect 11848 33917 12561 33969
rect 12613 33917 12639 33969
rect 12691 33917 14858 33969
rect 9762 33909 11152 33917
rect 9762 33905 10666 33909
rect 10722 33905 10747 33909
rect 10803 33905 10828 33909
rect 9762 33853 9801 33905
rect 9853 33853 9879 33905
rect 9931 33853 10666 33905
rect 10884 33853 10909 33909
rect 10965 33853 10990 33909
rect 11046 33853 11071 33909
rect 11127 33853 11152 33909
rect 11848 33905 14858 33917
rect 11848 33853 12561 33905
rect 12613 33853 12639 33905
rect 12691 33853 14858 33905
rect 9762 33841 11152 33853
rect 11848 33841 14858 33853
rect 9762 33789 9801 33841
rect 9853 33789 9879 33841
rect 9931 33829 10721 33841
rect 10773 33829 10799 33841
rect 10851 33829 11152 33841
rect 9931 33789 10666 33829
rect 9762 33777 10666 33789
rect 10722 33777 10747 33789
rect 10803 33777 10828 33789
rect 9762 33725 9801 33777
rect 9853 33725 9879 33777
rect 9931 33773 10666 33777
rect 10884 33773 10909 33829
rect 10965 33773 10990 33829
rect 11046 33773 11071 33829
rect 11127 33773 11152 33829
rect 11848 33789 12561 33841
rect 12613 33789 12639 33841
rect 12691 33789 14858 33841
rect 11848 33777 14858 33789
rect 9931 33749 10721 33773
rect 10773 33749 10799 33773
rect 10851 33749 11152 33773
rect 9931 33725 10666 33749
rect 9762 33713 10666 33725
rect 10722 33713 10747 33725
rect 10803 33713 10828 33725
rect 9762 33661 9801 33713
rect 9853 33661 9879 33713
rect 9931 33693 10666 33713
rect 10884 33693 10909 33749
rect 10965 33693 10990 33749
rect 11046 33693 11071 33749
rect 11127 33693 11152 33749
rect 11848 33725 12561 33777
rect 12613 33725 12639 33777
rect 12691 33725 14858 33777
rect 11848 33713 14858 33725
rect 9931 33669 10721 33693
rect 10773 33669 10799 33693
rect 10851 33669 11152 33693
rect 9931 33661 10666 33669
rect 9762 33649 10666 33661
rect 10722 33649 10747 33661
rect 10803 33649 10828 33661
rect 9762 33597 9801 33649
rect 9853 33597 9879 33649
rect 9931 33613 10666 33649
rect 10884 33613 10909 33669
rect 10965 33613 10990 33669
rect 11046 33613 11071 33669
rect 11127 33613 11152 33669
rect 11848 33661 12561 33713
rect 12613 33661 12639 33713
rect 12691 33661 14858 33713
rect 11848 33649 14858 33661
rect 9931 33597 10721 33613
rect 10773 33597 10799 33613
rect 10851 33597 11152 33613
rect 11848 33597 12561 33649
rect 12613 33597 12639 33649
rect 12691 33597 14858 33649
rect 9762 33589 11152 33597
rect 9762 33585 10666 33589
rect 10722 33585 10747 33589
rect 10803 33585 10828 33589
rect 9762 33533 9801 33585
rect 9853 33533 9879 33585
rect 9931 33533 10666 33585
rect 10884 33533 10909 33589
rect 10965 33533 10990 33589
rect 11046 33533 11071 33589
rect 11127 33533 11152 33589
rect 11848 33585 14858 33597
rect 11848 33533 12561 33585
rect 12613 33533 12639 33585
rect 12691 33533 14858 33585
rect 9762 33521 11152 33533
rect 11848 33521 14858 33533
rect 9762 33469 9801 33521
rect 9853 33469 9879 33521
rect 9931 33509 10721 33521
rect 10773 33509 10799 33521
rect 10851 33509 11152 33521
rect 9931 33469 10666 33509
rect 9762 33457 10666 33469
rect 10722 33457 10747 33469
rect 10803 33457 10828 33469
rect 9762 33405 9801 33457
rect 9853 33405 9879 33457
rect 9931 33453 10666 33457
rect 10884 33453 10909 33509
rect 10965 33453 10990 33509
rect 11046 33453 11071 33509
rect 11127 33453 11152 33509
rect 11848 33469 12561 33521
rect 12613 33469 12639 33521
rect 12691 33469 14858 33521
rect 11848 33457 14858 33469
rect 9931 33429 10721 33453
rect 10773 33429 10799 33453
rect 10851 33429 11152 33453
rect 9931 33405 10666 33429
rect 9762 33393 10666 33405
rect 10722 33393 10747 33405
rect 10803 33393 10828 33405
rect 9762 33341 9801 33393
rect 9853 33341 9879 33393
rect 9931 33373 10666 33393
rect 10884 33373 10909 33429
rect 10965 33373 10990 33429
rect 11046 33373 11071 33429
rect 11127 33373 11152 33429
rect 11848 33405 12561 33457
rect 12613 33405 12639 33457
rect 12691 33405 14858 33457
rect 11848 33393 14858 33405
rect 9931 33349 10721 33373
rect 10773 33349 10799 33373
rect 10851 33349 11152 33373
rect 9931 33341 10666 33349
rect 9762 33329 10666 33341
rect 10722 33329 10747 33341
rect 10803 33329 10828 33341
rect 9762 33277 9801 33329
rect 9853 33277 9879 33329
rect 9931 33293 10666 33329
rect 10884 33293 10909 33349
rect 10965 33293 10990 33349
rect 11046 33293 11071 33349
rect 11127 33293 11152 33349
rect 11848 33341 12561 33393
rect 12613 33341 12639 33393
rect 12691 33341 14858 33393
rect 11848 33329 14858 33341
rect 9931 33277 10721 33293
rect 10773 33277 10799 33293
rect 10851 33277 11152 33293
rect 11848 33277 12561 33329
rect 12613 33277 12639 33329
rect 12691 33277 14858 33329
rect 9762 33269 11152 33277
rect 9762 33264 10666 33269
rect 10722 33264 10747 33269
rect 10803 33264 10828 33269
rect 9762 33212 9801 33264
rect 9853 33212 9879 33264
rect 9931 33213 10666 33264
rect 10884 33213 10909 33269
rect 10965 33213 10990 33269
rect 11046 33213 11071 33269
rect 11127 33213 11152 33269
rect 11848 33264 14858 33277
rect 9931 33212 10721 33213
rect 10773 33212 10799 33213
rect 10851 33212 11152 33213
rect 11848 33212 12561 33264
rect 12613 33212 12639 33264
rect 12691 33212 14858 33264
rect 9762 33199 11152 33212
rect 11848 33199 14858 33212
rect 9762 33147 9801 33199
rect 9853 33147 9879 33199
rect 9931 33189 10721 33199
rect 10773 33189 10799 33199
rect 10851 33189 11152 33199
rect 9931 33147 10666 33189
rect 9762 33134 10666 33147
rect 10722 33134 10747 33147
rect 10803 33134 10828 33147
rect 9762 33082 9801 33134
rect 9853 33082 9879 33134
rect 9931 33133 10666 33134
rect 10884 33133 10909 33189
rect 10965 33133 10990 33189
rect 11046 33133 11071 33189
rect 11127 33133 11152 33189
rect 11848 33147 12561 33199
rect 12613 33147 12639 33199
rect 12691 33147 14858 33199
rect 11848 33134 14858 33147
rect 9931 33109 10721 33133
rect 10773 33109 10799 33133
rect 10851 33109 11152 33133
rect 9931 33082 10666 33109
rect 9762 33069 10666 33082
rect 10722 33069 10747 33082
rect 10803 33069 10828 33082
rect 9762 33017 9801 33069
rect 9853 33017 9879 33069
rect 9931 33053 10666 33069
rect 10884 33053 10909 33109
rect 10965 33053 10990 33109
rect 11046 33053 11071 33109
rect 11127 33053 11152 33109
rect 11848 33082 12561 33134
rect 12613 33082 12639 33134
rect 12691 33082 14858 33134
rect 11848 33069 14858 33082
rect 9931 33029 10721 33053
rect 10773 33029 10799 33053
rect 10851 33029 11152 33053
rect 9931 33017 10666 33029
rect 9762 33004 10666 33017
rect 10722 33004 10747 33017
rect 10803 33004 10828 33017
rect 9762 32952 9801 33004
rect 9853 32952 9879 33004
rect 9931 32973 10666 33004
rect 10884 32973 10909 33029
rect 10965 32973 10990 33029
rect 11046 32973 11071 33029
rect 11127 32973 11152 33029
rect 11848 33017 12561 33069
rect 12613 33017 12639 33069
rect 12691 33017 14858 33069
rect 11848 33004 14858 33017
rect 9931 32952 10721 32973
rect 10773 32952 10799 32973
rect 10851 32952 11152 32973
rect 11848 32952 12561 33004
rect 12613 32952 12639 33004
rect 12691 32952 14858 33004
rect 9762 32949 11152 32952
rect 9762 32939 10666 32949
rect 10722 32939 10747 32949
rect 10803 32939 10828 32949
rect 9762 32887 9801 32939
rect 9853 32887 9879 32939
rect 9931 32893 10666 32939
rect 10884 32893 10909 32949
rect 10965 32893 10990 32949
rect 11046 32893 11071 32949
rect 11127 32893 11152 32949
rect 11848 32939 14858 32952
rect 9931 32887 10721 32893
rect 10773 32887 10799 32893
rect 10851 32887 11152 32893
rect 11848 32887 12561 32939
rect 12613 32887 12639 32939
rect 12691 32887 14858 32939
rect 9762 32874 11152 32887
rect 11848 32874 14858 32887
rect 9762 32822 9801 32874
rect 9853 32822 9879 32874
rect 9931 32869 10721 32874
rect 10773 32869 10799 32874
rect 10851 32869 11152 32874
rect 9931 32822 10666 32869
rect 9762 32813 10666 32822
rect 10722 32813 10747 32822
rect 10803 32813 10828 32822
rect 10884 32813 10909 32869
rect 10965 32813 10990 32869
rect 11046 32813 11071 32869
rect 11127 32813 11152 32869
rect 11848 32822 12561 32874
rect 12613 32822 12639 32874
rect 12691 32822 14858 32874
rect 9762 32809 11152 32813
rect 11848 32809 14858 32822
rect 9762 32757 9801 32809
rect 9853 32757 9879 32809
rect 9931 32789 10721 32809
rect 10773 32789 10799 32809
rect 10851 32789 11152 32809
rect 9931 32757 10666 32789
rect 9762 32744 10666 32757
rect 10722 32744 10747 32757
rect 10803 32744 10828 32757
rect 9762 32692 9801 32744
rect 9853 32692 9879 32744
rect 9931 32733 10666 32744
rect 10884 32733 10909 32789
rect 10965 32733 10990 32789
rect 11046 32733 11071 32789
rect 11127 32733 11152 32789
rect 11848 32757 12561 32809
rect 12613 32757 12639 32809
rect 12691 32757 14858 32809
rect 11848 32744 14858 32757
rect 9931 32709 10721 32733
rect 10773 32709 10799 32733
rect 10851 32709 11152 32733
rect 9931 32692 10666 32709
rect 9762 32679 10666 32692
rect 10722 32679 10747 32692
rect 10803 32679 10828 32692
rect 9762 32627 9801 32679
rect 9853 32627 9879 32679
rect 9931 32653 10666 32679
rect 10884 32653 10909 32709
rect 10965 32653 10990 32709
rect 11046 32653 11071 32709
rect 11127 32653 11152 32709
rect 11848 32692 12561 32744
rect 12613 32692 12639 32744
rect 12691 32692 14858 32744
rect 11848 32679 14858 32692
rect 9931 32629 10721 32653
rect 10773 32629 10799 32653
rect 10851 32629 11152 32653
rect 9931 32627 10666 32629
rect 9762 32614 10666 32627
rect 10722 32614 10747 32627
rect 10803 32614 10828 32627
rect 9762 32562 9801 32614
rect 9853 32562 9879 32614
rect 9931 32573 10666 32614
rect 10884 32573 10909 32629
rect 10965 32573 10990 32629
rect 11046 32573 11071 32629
rect 11127 32573 11152 32629
rect 11848 32627 12561 32679
rect 12613 32627 12639 32679
rect 12691 32627 14858 32679
rect 11848 32614 14858 32627
rect 9931 32562 10721 32573
rect 10773 32562 10799 32573
rect 10851 32562 11152 32573
rect 11848 32562 12561 32614
rect 12613 32562 12639 32614
rect 12691 32562 14858 32614
rect 9762 32549 11152 32562
rect 11848 32549 14858 32562
rect 9762 32497 9801 32549
rect 9853 32497 9879 32549
rect 9931 32497 10666 32549
rect 9762 32493 10666 32497
rect 10722 32493 10747 32497
rect 10803 32493 10828 32497
rect 10884 32493 10909 32549
rect 10965 32493 10990 32549
rect 11046 32493 11071 32549
rect 11127 32493 11152 32549
rect 11848 32497 12561 32549
rect 12613 32497 12639 32549
rect 12691 32497 14858 32549
rect 11848 32493 14858 32497
rect 3361 32491 14858 32493
tri 2824 31774 3466 32416 sw
tri 11505 31774 12222 32491 ne
rect 187 31768 3466 31774
rect 187 31716 2872 31768
rect 2924 31716 2940 31768
rect 2992 31716 3008 31768
rect 3060 31716 3466 31768
rect 187 31704 3466 31716
rect 187 31652 2872 31704
rect 2924 31652 2940 31704
rect 2992 31652 3008 31704
rect 3060 31696 3466 31704
tri 3466 31696 3544 31774 sw
rect 3060 31694 11341 31696
rect 3060 31652 3109 31694
rect 187 31639 3109 31652
rect 187 31587 2872 31639
rect 2924 31587 2940 31639
rect 2992 31587 3008 31639
rect 3060 31638 3109 31639
rect 3165 31638 3190 31694
rect 3246 31638 3271 31694
rect 3327 31638 3352 31694
rect 3408 31638 3433 31694
rect 3489 31638 3514 31694
rect 4290 31690 5195 31694
rect 4290 31638 4712 31690
rect 4764 31638 4780 31690
rect 4832 31638 4848 31690
rect 4900 31638 5195 31690
rect 5251 31638 5276 31694
rect 5332 31638 5357 31694
rect 5413 31638 5438 31694
rect 5494 31638 5519 31694
rect 5575 31638 5600 31694
rect 6376 31690 11341 31694
rect 6376 31638 6552 31690
rect 6604 31638 6620 31690
rect 6672 31638 6688 31690
rect 6740 31638 7472 31690
rect 7524 31638 7540 31690
rect 7592 31638 7608 31690
rect 7660 31638 8392 31690
rect 8444 31638 8460 31690
rect 8512 31638 8528 31690
rect 8580 31638 9312 31690
rect 9364 31638 9380 31690
rect 9432 31638 9448 31690
rect 9500 31638 10232 31690
rect 10284 31638 10300 31690
rect 10352 31638 10368 31690
rect 10420 31638 11152 31690
rect 11204 31638 11220 31690
rect 11272 31638 11288 31690
rect 11340 31638 11341 31690
rect 3060 31614 3514 31638
rect 4290 31626 5600 31638
rect 6376 31626 11341 31638
rect 3060 31587 3109 31614
rect 187 31574 3109 31587
rect 187 31522 2872 31574
rect 2924 31522 2940 31574
rect 2992 31522 3008 31574
rect 3060 31558 3109 31574
rect 3165 31558 3190 31614
rect 3246 31558 3271 31614
rect 3327 31558 3352 31614
rect 3408 31558 3433 31614
rect 3489 31558 3514 31614
rect 4290 31574 4712 31626
rect 4764 31574 4780 31626
rect 4832 31574 4848 31626
rect 4900 31614 5600 31626
rect 4900 31574 5195 31614
rect 4290 31562 5195 31574
rect 3060 31534 3514 31558
rect 3060 31522 3109 31534
rect 187 31509 3109 31522
rect 187 31457 2872 31509
rect 2924 31457 2940 31509
rect 2992 31457 3008 31509
rect 3060 31478 3109 31509
rect 3165 31478 3190 31534
rect 3246 31478 3271 31534
rect 3327 31478 3352 31534
rect 3408 31478 3433 31534
rect 3489 31478 3514 31534
rect 4290 31510 4712 31562
rect 4764 31510 4780 31562
rect 4832 31510 4848 31562
rect 4900 31558 5195 31562
rect 5251 31558 5276 31614
rect 5332 31558 5357 31614
rect 5413 31558 5438 31614
rect 5494 31558 5519 31614
rect 5575 31558 5600 31614
rect 6376 31574 6552 31626
rect 6604 31574 6620 31626
rect 6672 31574 6688 31626
rect 6740 31574 7472 31626
rect 7524 31574 7540 31626
rect 7592 31574 7608 31626
rect 7660 31574 8392 31626
rect 8444 31574 8460 31626
rect 8512 31574 8528 31626
rect 8580 31574 9312 31626
rect 9364 31574 9380 31626
rect 9432 31574 9448 31626
rect 9500 31574 10232 31626
rect 10284 31574 10300 31626
rect 10352 31574 10368 31626
rect 10420 31574 11152 31626
rect 11204 31574 11220 31626
rect 11272 31574 11288 31626
rect 11340 31574 11341 31626
rect 6376 31562 11341 31574
rect 4900 31534 5600 31558
rect 4900 31510 5195 31534
rect 4290 31498 5195 31510
rect 3060 31457 3514 31478
rect 187 31454 3514 31457
rect 187 31444 3109 31454
rect 187 31392 2872 31444
rect 2924 31392 2940 31444
rect 2992 31392 3008 31444
rect 3060 31398 3109 31444
rect 3165 31398 3190 31454
rect 3246 31398 3271 31454
rect 3327 31398 3352 31454
rect 3408 31398 3433 31454
rect 3489 31398 3514 31454
rect 4290 31446 4712 31498
rect 4764 31446 4780 31498
rect 4832 31446 4848 31498
rect 4900 31478 5195 31498
rect 5251 31478 5276 31534
rect 5332 31478 5357 31534
rect 5413 31478 5438 31534
rect 5494 31478 5519 31534
rect 5575 31478 5600 31534
rect 6376 31510 6552 31562
rect 6604 31510 6620 31562
rect 6672 31510 6688 31562
rect 6740 31510 7472 31562
rect 7524 31510 7540 31562
rect 7592 31510 7608 31562
rect 7660 31510 8392 31562
rect 8444 31510 8460 31562
rect 8512 31510 8528 31562
rect 8580 31510 9312 31562
rect 9364 31510 9380 31562
rect 9432 31510 9448 31562
rect 9500 31510 10232 31562
rect 10284 31510 10300 31562
rect 10352 31510 10368 31562
rect 10420 31510 11152 31562
rect 11204 31510 11220 31562
rect 11272 31510 11288 31562
rect 11340 31510 11341 31562
rect 6376 31498 11341 31510
rect 4900 31454 5600 31478
rect 4900 31446 5195 31454
rect 4290 31434 5195 31446
rect 3060 31392 3514 31398
rect 187 31379 3514 31392
rect 4290 31382 4712 31434
rect 4764 31382 4780 31434
rect 4832 31382 4848 31434
rect 4900 31398 5195 31434
rect 5251 31398 5276 31454
rect 5332 31398 5357 31454
rect 5413 31398 5438 31454
rect 5494 31398 5519 31454
rect 5575 31398 5600 31454
rect 6376 31446 6552 31498
rect 6604 31446 6620 31498
rect 6672 31446 6688 31498
rect 6740 31446 7472 31498
rect 7524 31446 7540 31498
rect 7592 31446 7608 31498
rect 7660 31446 8392 31498
rect 8444 31446 8460 31498
rect 8512 31446 8528 31498
rect 8580 31446 9312 31498
rect 9364 31446 9380 31498
rect 9432 31446 9448 31498
rect 9500 31446 10232 31498
rect 10284 31446 10300 31498
rect 10352 31446 10368 31498
rect 10420 31446 11152 31498
rect 11204 31446 11220 31498
rect 11272 31446 11288 31498
rect 11340 31446 11341 31498
rect 6376 31434 11341 31446
rect 4900 31382 5600 31398
rect 6376 31382 6552 31434
rect 6604 31382 6620 31434
rect 6672 31382 6688 31434
rect 6740 31382 7472 31434
rect 7524 31382 7540 31434
rect 7592 31382 7608 31434
rect 7660 31382 8392 31434
rect 8444 31382 8460 31434
rect 8512 31382 8528 31434
rect 8580 31382 9312 31434
rect 9364 31382 9380 31434
rect 9432 31382 9448 31434
rect 9500 31382 10232 31434
rect 10284 31382 10300 31434
rect 10352 31382 10368 31434
rect 10420 31382 11152 31434
rect 11204 31382 11220 31434
rect 11272 31382 11288 31434
rect 11340 31382 11341 31434
rect 187 31327 2872 31379
rect 2924 31327 2940 31379
rect 2992 31327 3008 31379
rect 3060 31374 3514 31379
rect 3060 31327 3109 31374
rect 187 31318 3109 31327
rect 3165 31318 3190 31374
rect 3246 31318 3271 31374
rect 3327 31318 3352 31374
rect 3408 31318 3433 31374
rect 3489 31318 3514 31374
rect 4290 31374 5600 31382
rect 4290 31370 5195 31374
rect 4290 31318 4712 31370
rect 4764 31318 4780 31370
rect 4832 31318 4848 31370
rect 4900 31318 5195 31370
rect 5251 31318 5276 31374
rect 5332 31318 5357 31374
rect 5413 31318 5438 31374
rect 5494 31318 5519 31374
rect 5575 31318 5600 31374
rect 6376 31370 11341 31382
rect 6376 31318 6552 31370
rect 6604 31318 6620 31370
rect 6672 31318 6688 31370
rect 6740 31318 7472 31370
rect 7524 31318 7540 31370
rect 7592 31318 7608 31370
rect 7660 31318 8392 31370
rect 8444 31318 8460 31370
rect 8512 31318 8528 31370
rect 8580 31318 9312 31370
rect 9364 31318 9380 31370
rect 9432 31318 9448 31370
rect 9500 31318 10232 31370
rect 10284 31318 10300 31370
rect 10352 31318 10368 31370
rect 10420 31318 11152 31370
rect 11204 31318 11220 31370
rect 11272 31318 11288 31370
rect 11340 31318 11341 31370
rect 187 31314 3514 31318
rect 187 31262 2872 31314
rect 2924 31262 2940 31314
rect 2992 31262 3008 31314
rect 3060 31294 3514 31314
rect 4290 31306 5600 31318
rect 6376 31306 11341 31318
rect 3060 31262 3109 31294
rect 187 31249 3109 31262
rect 187 31197 2872 31249
rect 2924 31197 2940 31249
rect 2992 31197 3008 31249
rect 3060 31238 3109 31249
rect 3165 31238 3190 31294
rect 3246 31238 3271 31294
rect 3327 31238 3352 31294
rect 3408 31238 3433 31294
rect 3489 31238 3514 31294
rect 4290 31254 4712 31306
rect 4764 31254 4780 31306
rect 4832 31254 4848 31306
rect 4900 31294 5600 31306
rect 4900 31254 5195 31294
rect 4290 31242 5195 31254
rect 3060 31214 3514 31238
rect 3060 31197 3109 31214
rect 187 31184 3109 31197
rect 187 31132 2872 31184
rect 2924 31132 2940 31184
rect 2992 31132 3008 31184
rect 3060 31158 3109 31184
rect 3165 31158 3190 31214
rect 3246 31158 3271 31214
rect 3327 31158 3352 31214
rect 3408 31158 3433 31214
rect 3489 31158 3514 31214
rect 4290 31190 4712 31242
rect 4764 31190 4780 31242
rect 4832 31190 4848 31242
rect 4900 31238 5195 31242
rect 5251 31238 5276 31294
rect 5332 31238 5357 31294
rect 5413 31238 5438 31294
rect 5494 31238 5519 31294
rect 5575 31238 5600 31294
rect 6376 31254 6552 31306
rect 6604 31254 6620 31306
rect 6672 31254 6688 31306
rect 6740 31254 7472 31306
rect 7524 31254 7540 31306
rect 7592 31254 7608 31306
rect 7660 31254 8392 31306
rect 8444 31254 8460 31306
rect 8512 31254 8528 31306
rect 8580 31254 9312 31306
rect 9364 31254 9380 31306
rect 9432 31254 9448 31306
rect 9500 31254 10232 31306
rect 10284 31254 10300 31306
rect 10352 31254 10368 31306
rect 10420 31254 11152 31306
rect 11204 31254 11220 31306
rect 11272 31254 11288 31306
rect 11340 31254 11341 31306
rect 6376 31242 11341 31254
rect 4900 31214 5600 31238
rect 4900 31190 5195 31214
rect 4290 31178 5195 31190
rect 3060 31134 3514 31158
rect 3060 31132 3109 31134
rect 187 31119 3109 31132
rect 187 31067 2872 31119
rect 2924 31067 2940 31119
rect 2992 31067 3008 31119
rect 3060 31078 3109 31119
rect 3165 31078 3190 31134
rect 3246 31078 3271 31134
rect 3327 31078 3352 31134
rect 3408 31078 3433 31134
rect 3489 31078 3514 31134
rect 4290 31126 4712 31178
rect 4764 31126 4780 31178
rect 4832 31126 4848 31178
rect 4900 31158 5195 31178
rect 5251 31158 5276 31214
rect 5332 31158 5357 31214
rect 5413 31158 5438 31214
rect 5494 31158 5519 31214
rect 5575 31158 5600 31214
rect 6376 31190 6552 31242
rect 6604 31190 6620 31242
rect 6672 31190 6688 31242
rect 6740 31190 7472 31242
rect 7524 31190 7540 31242
rect 7592 31190 7608 31242
rect 7660 31190 8392 31242
rect 8444 31190 8460 31242
rect 8512 31190 8528 31242
rect 8580 31190 9312 31242
rect 9364 31190 9380 31242
rect 9432 31190 9448 31242
rect 9500 31190 10232 31242
rect 10284 31190 10300 31242
rect 10352 31190 10368 31242
rect 10420 31190 11152 31242
rect 11204 31190 11220 31242
rect 11272 31190 11288 31242
rect 11340 31190 11341 31242
rect 6376 31178 11341 31190
rect 4900 31134 5600 31158
rect 4900 31126 5195 31134
rect 4290 31114 5195 31126
rect 3060 31067 3514 31078
rect 187 31054 3514 31067
rect 4290 31062 4712 31114
rect 4764 31062 4780 31114
rect 4832 31062 4848 31114
rect 4900 31078 5195 31114
rect 5251 31078 5276 31134
rect 5332 31078 5357 31134
rect 5413 31078 5438 31134
rect 5494 31078 5519 31134
rect 5575 31078 5600 31134
rect 6376 31126 6552 31178
rect 6604 31126 6620 31178
rect 6672 31126 6688 31178
rect 6740 31126 7472 31178
rect 7524 31126 7540 31178
rect 7592 31126 7608 31178
rect 7660 31126 8392 31178
rect 8444 31126 8460 31178
rect 8512 31126 8528 31178
rect 8580 31126 9312 31178
rect 9364 31126 9380 31178
rect 9432 31126 9448 31178
rect 9500 31126 10232 31178
rect 10284 31126 10300 31178
rect 10352 31126 10368 31178
rect 10420 31126 11152 31178
rect 11204 31126 11220 31178
rect 11272 31126 11288 31178
rect 11340 31126 11341 31178
rect 6376 31114 11341 31126
rect 4900 31062 5600 31078
rect 6376 31062 6552 31114
rect 6604 31062 6620 31114
rect 6672 31062 6688 31114
rect 6740 31062 7472 31114
rect 7524 31062 7540 31114
rect 7592 31062 7608 31114
rect 7660 31062 8392 31114
rect 8444 31062 8460 31114
rect 8512 31062 8528 31114
rect 8580 31062 9312 31114
rect 9364 31062 9380 31114
rect 9432 31062 9448 31114
rect 9500 31062 10232 31114
rect 10284 31062 10300 31114
rect 10352 31062 10368 31114
rect 10420 31062 11152 31114
rect 11204 31062 11220 31114
rect 11272 31062 11288 31114
rect 11340 31062 11341 31114
rect 187 31002 2872 31054
rect 2924 31002 2940 31054
rect 2992 31002 3008 31054
rect 3060 31002 3109 31054
rect 187 30998 3109 31002
rect 3165 30998 3190 31054
rect 3246 30998 3271 31054
rect 3327 30998 3352 31054
rect 3408 30998 3433 31054
rect 3489 30998 3514 31054
rect 4290 31054 5600 31062
rect 4290 31050 5195 31054
rect 4290 30998 4712 31050
rect 4764 30998 4780 31050
rect 4832 30998 4848 31050
rect 4900 30998 5195 31050
rect 5251 30998 5276 31054
rect 5332 30998 5357 31054
rect 5413 30998 5438 31054
rect 5494 30998 5519 31054
rect 5575 30998 5600 31054
rect 6376 31050 11341 31062
rect 6376 30998 6552 31050
rect 6604 30998 6620 31050
rect 6672 30998 6688 31050
rect 6740 30998 7472 31050
rect 7524 30998 7540 31050
rect 7592 30998 7608 31050
rect 7660 30998 8392 31050
rect 8444 30998 8460 31050
rect 8512 30998 8528 31050
rect 8580 30998 9312 31050
rect 9364 30998 9380 31050
rect 9432 30998 9448 31050
rect 9500 30998 10232 31050
rect 10284 30998 10300 31050
rect 10352 30998 10368 31050
rect 10420 30998 11152 31050
rect 11204 30998 11220 31050
rect 11272 30998 11288 31050
rect 11340 30998 11341 31050
rect 187 30989 3514 30998
rect 187 30937 2872 30989
rect 2924 30937 2940 30989
rect 2992 30937 3008 30989
rect 3060 30974 3514 30989
rect 4290 30986 5600 30998
rect 6376 30986 11341 30998
rect 3060 30937 3109 30974
rect 187 30924 3109 30937
rect 187 30872 2872 30924
rect 2924 30872 2940 30924
rect 2992 30872 3008 30924
rect 3060 30918 3109 30924
rect 3165 30918 3190 30974
rect 3246 30918 3271 30974
rect 3327 30918 3352 30974
rect 3408 30918 3433 30974
rect 3489 30918 3514 30974
rect 4290 30934 4712 30986
rect 4764 30934 4780 30986
rect 4832 30934 4848 30986
rect 4900 30974 5600 30986
rect 4900 30934 5195 30974
rect 4290 30922 5195 30934
rect 3060 30894 3514 30918
rect 3060 30872 3109 30894
rect 187 30859 3109 30872
rect 187 30807 2872 30859
rect 2924 30807 2940 30859
rect 2992 30807 3008 30859
rect 3060 30838 3109 30859
rect 3165 30838 3190 30894
rect 3246 30838 3271 30894
rect 3327 30838 3352 30894
rect 3408 30838 3433 30894
rect 3489 30838 3514 30894
rect 4290 30870 4712 30922
rect 4764 30870 4780 30922
rect 4832 30870 4848 30922
rect 4900 30918 5195 30922
rect 5251 30918 5276 30974
rect 5332 30918 5357 30974
rect 5413 30918 5438 30974
rect 5494 30918 5519 30974
rect 5575 30918 5600 30974
rect 6376 30934 6552 30986
rect 6604 30934 6620 30986
rect 6672 30934 6688 30986
rect 6740 30934 7472 30986
rect 7524 30934 7540 30986
rect 7592 30934 7608 30986
rect 7660 30934 8392 30986
rect 8444 30934 8460 30986
rect 8512 30934 8528 30986
rect 8580 30934 9312 30986
rect 9364 30934 9380 30986
rect 9432 30934 9448 30986
rect 9500 30934 10232 30986
rect 10284 30934 10300 30986
rect 10352 30934 10368 30986
rect 10420 30934 11152 30986
rect 11204 30934 11220 30986
rect 11272 30934 11288 30986
rect 11340 30934 11341 30986
rect 6376 30922 11341 30934
rect 4900 30894 5600 30918
rect 4900 30870 5195 30894
rect 4290 30858 5195 30870
rect 3060 30814 3514 30838
rect 3060 30807 3109 30814
rect 187 30794 3109 30807
rect 187 30742 2872 30794
rect 2924 30742 2940 30794
rect 2992 30742 3008 30794
rect 3060 30758 3109 30794
rect 3165 30758 3190 30814
rect 3246 30758 3271 30814
rect 3327 30758 3352 30814
rect 3408 30758 3433 30814
rect 3489 30758 3514 30814
rect 4290 30806 4712 30858
rect 4764 30806 4780 30858
rect 4832 30806 4848 30858
rect 4900 30838 5195 30858
rect 5251 30838 5276 30894
rect 5332 30838 5357 30894
rect 5413 30838 5438 30894
rect 5494 30838 5519 30894
rect 5575 30838 5600 30894
rect 6376 30870 6552 30922
rect 6604 30870 6620 30922
rect 6672 30870 6688 30922
rect 6740 30870 7472 30922
rect 7524 30870 7540 30922
rect 7592 30870 7608 30922
rect 7660 30870 8392 30922
rect 8444 30870 8460 30922
rect 8512 30870 8528 30922
rect 8580 30870 9312 30922
rect 9364 30870 9380 30922
rect 9432 30870 9448 30922
rect 9500 30870 10232 30922
rect 10284 30870 10300 30922
rect 10352 30870 10368 30922
rect 10420 30870 11152 30922
rect 11204 30870 11220 30922
rect 11272 30870 11288 30922
rect 11340 30870 11341 30922
rect 6376 30858 11341 30870
rect 4900 30814 5600 30838
rect 4900 30806 5195 30814
rect 4290 30794 5195 30806
rect 3060 30742 3514 30758
rect 4290 30742 4712 30794
rect 4764 30742 4780 30794
rect 4832 30742 4848 30794
rect 4900 30758 5195 30794
rect 5251 30758 5276 30814
rect 5332 30758 5357 30814
rect 5413 30758 5438 30814
rect 5494 30758 5519 30814
rect 5575 30758 5600 30814
rect 6376 30806 6552 30858
rect 6604 30806 6620 30858
rect 6672 30806 6688 30858
rect 6740 30806 7472 30858
rect 7524 30806 7540 30858
rect 7592 30806 7608 30858
rect 7660 30806 8392 30858
rect 8444 30806 8460 30858
rect 8512 30806 8528 30858
rect 8580 30806 9312 30858
rect 9364 30806 9380 30858
rect 9432 30806 9448 30858
rect 9500 30806 10232 30858
rect 10284 30806 10300 30858
rect 10352 30806 10368 30858
rect 10420 30806 11152 30858
rect 11204 30806 11220 30858
rect 11272 30806 11288 30858
rect 11340 30806 11341 30858
rect 6376 30794 11341 30806
rect 4900 30742 5600 30758
rect 6376 30742 6552 30794
rect 6604 30742 6620 30794
rect 6672 30742 6688 30794
rect 6740 30742 7472 30794
rect 7524 30742 7540 30794
rect 7592 30742 7608 30794
rect 7660 30742 8392 30794
rect 8444 30742 8460 30794
rect 8512 30742 8528 30794
rect 8580 30742 9312 30794
rect 9364 30742 9380 30794
rect 9432 30742 9448 30794
rect 9500 30742 10232 30794
rect 10284 30742 10300 30794
rect 10352 30742 10368 30794
rect 10420 30742 11152 30794
rect 11204 30742 11220 30794
rect 11272 30742 11288 30794
rect 11340 30742 11341 30794
rect 187 30734 3514 30742
rect 187 30729 3109 30734
rect 187 30677 2872 30729
rect 2924 30677 2940 30729
rect 2992 30677 3008 30729
rect 3060 30678 3109 30729
rect 3165 30678 3190 30734
rect 3246 30678 3271 30734
rect 3327 30678 3352 30734
rect 3408 30678 3433 30734
rect 3489 30678 3514 30734
rect 4290 30734 5600 30742
rect 4290 30729 5195 30734
rect 3060 30677 3514 30678
rect 4290 30677 4712 30729
rect 4764 30677 4780 30729
rect 4832 30677 4848 30729
rect 4900 30678 5195 30729
rect 5251 30678 5276 30734
rect 5332 30678 5357 30734
rect 5413 30678 5438 30734
rect 5494 30678 5519 30734
rect 5575 30678 5600 30734
rect 6376 30729 11341 30742
rect 4900 30677 5600 30678
rect 6376 30677 6552 30729
rect 6604 30677 6620 30729
rect 6672 30677 6688 30729
rect 6740 30677 7472 30729
rect 7524 30677 7540 30729
rect 7592 30677 7608 30729
rect 7660 30677 8392 30729
rect 8444 30677 8460 30729
rect 8512 30677 8528 30729
rect 8580 30677 9312 30729
rect 9364 30677 9380 30729
rect 9432 30677 9448 30729
rect 9500 30677 10232 30729
rect 10284 30677 10300 30729
rect 10352 30677 10368 30729
rect 10420 30677 11152 30729
rect 11204 30677 11220 30729
rect 11272 30677 11288 30729
rect 11340 30677 11341 30729
rect 187 30664 3514 30677
rect 4290 30664 5600 30677
rect 6376 30664 11341 30677
rect 187 30612 2872 30664
rect 2924 30612 2940 30664
rect 2992 30612 3008 30664
rect 3060 30654 3514 30664
rect 3060 30612 3109 30654
rect 187 30599 3109 30612
rect 187 30547 2872 30599
rect 2924 30547 2940 30599
rect 2992 30547 3008 30599
rect 3060 30598 3109 30599
rect 3165 30598 3190 30654
rect 3246 30598 3271 30654
rect 3327 30598 3352 30654
rect 3408 30598 3433 30654
rect 3489 30598 3514 30654
rect 4290 30612 4712 30664
rect 4764 30612 4780 30664
rect 4832 30612 4848 30664
rect 4900 30654 5600 30664
rect 4900 30612 5195 30654
rect 4290 30599 5195 30612
rect 3060 30574 3514 30598
rect 3060 30547 3109 30574
rect 187 30534 3109 30547
rect 187 30482 2872 30534
rect 2924 30482 2940 30534
rect 2992 30482 3008 30534
rect 3060 30518 3109 30534
rect 3165 30518 3190 30574
rect 3246 30518 3271 30574
rect 3327 30518 3352 30574
rect 3408 30518 3433 30574
rect 3489 30518 3514 30574
rect 4290 30547 4712 30599
rect 4764 30547 4780 30599
rect 4832 30547 4848 30599
rect 4900 30598 5195 30599
rect 5251 30598 5276 30654
rect 5332 30598 5357 30654
rect 5413 30598 5438 30654
rect 5494 30598 5519 30654
rect 5575 30598 5600 30654
rect 6376 30612 6552 30664
rect 6604 30612 6620 30664
rect 6672 30612 6688 30664
rect 6740 30612 7472 30664
rect 7524 30612 7540 30664
rect 7592 30612 7608 30664
rect 7660 30612 8392 30664
rect 8444 30612 8460 30664
rect 8512 30612 8528 30664
rect 8580 30612 9312 30664
rect 9364 30612 9380 30664
rect 9432 30612 9448 30664
rect 9500 30612 10232 30664
rect 10284 30612 10300 30664
rect 10352 30612 10368 30664
rect 10420 30612 11152 30664
rect 11204 30612 11220 30664
rect 11272 30612 11288 30664
rect 11340 30612 11341 30664
rect 6376 30599 11341 30612
rect 4900 30574 5600 30598
rect 4900 30547 5195 30574
rect 4290 30534 5195 30547
rect 3060 30494 3514 30518
rect 3060 30482 3109 30494
rect 187 30469 3109 30482
rect 187 30417 2872 30469
rect 2924 30417 2940 30469
rect 2992 30417 3008 30469
rect 3060 30438 3109 30469
rect 3165 30438 3190 30494
rect 3246 30438 3271 30494
rect 3327 30438 3352 30494
rect 3408 30438 3433 30494
rect 3489 30438 3514 30494
rect 4290 30482 4712 30534
rect 4764 30482 4780 30534
rect 4832 30482 4848 30534
rect 4900 30518 5195 30534
rect 5251 30518 5276 30574
rect 5332 30518 5357 30574
rect 5413 30518 5438 30574
rect 5494 30518 5519 30574
rect 5575 30518 5600 30574
rect 6376 30547 6552 30599
rect 6604 30547 6620 30599
rect 6672 30547 6688 30599
rect 6740 30547 7472 30599
rect 7524 30547 7540 30599
rect 7592 30547 7608 30599
rect 7660 30547 8392 30599
rect 8444 30547 8460 30599
rect 8512 30547 8528 30599
rect 8580 30547 9312 30599
rect 9364 30547 9380 30599
rect 9432 30547 9448 30599
rect 9500 30547 10232 30599
rect 10284 30547 10300 30599
rect 10352 30547 10368 30599
rect 10420 30547 11152 30599
rect 11204 30547 11220 30599
rect 11272 30547 11288 30599
rect 11340 30547 11341 30599
rect 6376 30534 11341 30547
rect 4900 30494 5600 30518
rect 4900 30482 5195 30494
rect 4290 30469 5195 30482
rect 3060 30417 3514 30438
rect 4290 30417 4712 30469
rect 4764 30417 4780 30469
rect 4832 30417 4848 30469
rect 4900 30438 5195 30469
rect 5251 30438 5276 30494
rect 5332 30438 5357 30494
rect 5413 30438 5438 30494
rect 5494 30438 5519 30494
rect 5575 30438 5600 30494
rect 6376 30482 6552 30534
rect 6604 30482 6620 30534
rect 6672 30482 6688 30534
rect 6740 30482 7472 30534
rect 7524 30482 7540 30534
rect 7592 30482 7608 30534
rect 7660 30482 8392 30534
rect 8444 30482 8460 30534
rect 8512 30482 8528 30534
rect 8580 30482 9312 30534
rect 9364 30482 9380 30534
rect 9432 30482 9448 30534
rect 9500 30482 10232 30534
rect 10284 30482 10300 30534
rect 10352 30482 10368 30534
rect 10420 30482 11152 30534
rect 11204 30482 11220 30534
rect 11272 30482 11288 30534
rect 11340 30482 11341 30534
rect 6376 30469 11341 30482
rect 4900 30417 5600 30438
rect 6376 30417 6552 30469
rect 6604 30417 6620 30469
rect 6672 30417 6688 30469
rect 6740 30417 7472 30469
rect 7524 30417 7540 30469
rect 7592 30417 7608 30469
rect 7660 30417 8392 30469
rect 8444 30417 8460 30469
rect 8512 30417 8528 30469
rect 8580 30417 9312 30469
rect 9364 30417 9380 30469
rect 9432 30417 9448 30469
rect 9500 30417 10232 30469
rect 10284 30417 10300 30469
rect 10352 30417 10368 30469
rect 10420 30417 11152 30469
rect 11204 30417 11220 30469
rect 11272 30417 11288 30469
rect 11340 30417 11341 30469
rect 187 30414 3514 30417
rect 187 30404 3109 30414
rect 187 30352 2872 30404
rect 2924 30352 2940 30404
rect 2992 30352 3008 30404
rect 3060 30358 3109 30404
rect 3165 30358 3190 30414
rect 3246 30358 3271 30414
rect 3327 30358 3352 30414
rect 3408 30358 3433 30414
rect 3489 30358 3514 30414
rect 4290 30414 5600 30417
rect 4290 30404 5195 30414
rect 3060 30352 3514 30358
rect 4290 30352 4712 30404
rect 4764 30352 4780 30404
rect 4832 30352 4848 30404
rect 4900 30358 5195 30404
rect 5251 30358 5276 30414
rect 5332 30358 5357 30414
rect 5413 30358 5438 30414
rect 5494 30358 5519 30414
rect 5575 30358 5600 30414
rect 6376 30404 11341 30417
rect 4900 30352 5600 30358
rect 6376 30352 6552 30404
rect 6604 30352 6620 30404
rect 6672 30352 6688 30404
rect 6740 30352 7472 30404
rect 7524 30352 7540 30404
rect 7592 30352 7608 30404
rect 7660 30352 8392 30404
rect 8444 30352 8460 30404
rect 8512 30352 8528 30404
rect 8580 30352 9312 30404
rect 9364 30352 9380 30404
rect 9432 30352 9448 30404
rect 9500 30352 10232 30404
rect 10284 30352 10300 30404
rect 10352 30352 10368 30404
rect 10420 30352 11152 30404
rect 11204 30352 11220 30404
rect 11272 30352 11288 30404
rect 11340 30352 11341 30404
rect 187 30339 3514 30352
rect 4290 30339 5600 30352
rect 6376 30339 11341 30352
rect 187 30287 2872 30339
rect 2924 30287 2940 30339
rect 2992 30287 3008 30339
rect 3060 30334 3514 30339
rect 3060 30287 3109 30334
rect 187 30278 3109 30287
rect 3165 30278 3190 30334
rect 3246 30278 3271 30334
rect 3327 30278 3352 30334
rect 3408 30278 3433 30334
rect 3489 30278 3514 30334
rect 4290 30287 4712 30339
rect 4764 30287 4780 30339
rect 4832 30287 4848 30339
rect 4900 30334 5600 30339
rect 4900 30287 5195 30334
rect 187 30274 3514 30278
rect 4290 30278 5195 30287
rect 5251 30278 5276 30334
rect 5332 30278 5357 30334
rect 5413 30278 5438 30334
rect 5494 30278 5519 30334
rect 5575 30278 5600 30334
rect 6376 30287 6552 30339
rect 6604 30287 6620 30339
rect 6672 30287 6688 30339
rect 6740 30287 7472 30339
rect 7524 30287 7540 30339
rect 7592 30287 7608 30339
rect 7660 30287 8392 30339
rect 8444 30287 8460 30339
rect 8512 30287 8528 30339
rect 8580 30287 9312 30339
rect 9364 30287 9380 30339
rect 9432 30287 9448 30339
rect 9500 30287 10232 30339
rect 10284 30287 10300 30339
rect 10352 30287 10368 30339
rect 10420 30287 11152 30339
rect 11204 30287 11220 30339
rect 11272 30287 11288 30339
rect 11340 30287 11341 30339
rect 4290 30274 5600 30278
rect 6376 30274 11341 30287
rect 187 30222 2872 30274
rect 2924 30222 2940 30274
rect 2992 30222 3008 30274
rect 3060 30254 3514 30274
rect 3060 30222 3109 30254
rect 187 30209 3109 30222
rect 187 30157 2872 30209
rect 2924 30157 2940 30209
rect 2992 30157 3008 30209
rect 3060 30198 3109 30209
rect 3165 30198 3190 30254
rect 3246 30198 3271 30254
rect 3327 30198 3352 30254
rect 3408 30198 3433 30254
rect 3489 30198 3514 30254
rect 4290 30222 4712 30274
rect 4764 30222 4780 30274
rect 4832 30222 4848 30274
rect 4900 30254 5600 30274
rect 4900 30222 5195 30254
rect 4290 30209 5195 30222
rect 3060 30174 3514 30198
rect 3060 30157 3109 30174
rect 187 30144 3109 30157
rect 187 30092 2872 30144
rect 2924 30092 2940 30144
rect 2992 30092 3008 30144
rect 3060 30118 3109 30144
rect 3165 30118 3190 30174
rect 3246 30118 3271 30174
rect 3327 30118 3352 30174
rect 3408 30118 3433 30174
rect 3489 30118 3514 30174
rect 4290 30157 4712 30209
rect 4764 30157 4780 30209
rect 4832 30157 4848 30209
rect 4900 30198 5195 30209
rect 5251 30198 5276 30254
rect 5332 30198 5357 30254
rect 5413 30198 5438 30254
rect 5494 30198 5519 30254
rect 5575 30198 5600 30254
rect 6376 30222 6552 30274
rect 6604 30222 6620 30274
rect 6672 30222 6688 30274
rect 6740 30222 7472 30274
rect 7524 30222 7540 30274
rect 7592 30222 7608 30274
rect 7660 30222 8392 30274
rect 8444 30222 8460 30274
rect 8512 30222 8528 30274
rect 8580 30222 9312 30274
rect 9364 30222 9380 30274
rect 9432 30222 9448 30274
rect 9500 30222 10232 30274
rect 10284 30222 10300 30274
rect 10352 30222 10368 30274
rect 10420 30222 11152 30274
rect 11204 30222 11220 30274
rect 11272 30222 11288 30274
rect 11340 30222 11341 30274
rect 6376 30209 11341 30222
rect 4900 30174 5600 30198
rect 4900 30157 5195 30174
rect 4290 30144 5195 30157
rect 3060 30094 3514 30118
rect 3060 30092 3109 30094
rect 187 30079 3109 30092
rect 187 30027 2872 30079
rect 2924 30027 2940 30079
rect 2992 30027 3008 30079
rect 3060 30038 3109 30079
rect 3165 30038 3190 30094
rect 3246 30038 3271 30094
rect 3327 30038 3352 30094
rect 3408 30038 3433 30094
rect 3489 30038 3514 30094
rect 4290 30092 4712 30144
rect 4764 30092 4780 30144
rect 4832 30092 4848 30144
rect 4900 30118 5195 30144
rect 5251 30118 5276 30174
rect 5332 30118 5357 30174
rect 5413 30118 5438 30174
rect 5494 30118 5519 30174
rect 5575 30118 5600 30174
rect 6376 30157 6552 30209
rect 6604 30157 6620 30209
rect 6672 30157 6688 30209
rect 6740 30157 7472 30209
rect 7524 30157 7540 30209
rect 7592 30157 7608 30209
rect 7660 30157 8392 30209
rect 8444 30157 8460 30209
rect 8512 30157 8528 30209
rect 8580 30157 9312 30209
rect 9364 30157 9380 30209
rect 9432 30157 9448 30209
rect 9500 30157 10232 30209
rect 10284 30157 10300 30209
rect 10352 30157 10368 30209
rect 10420 30157 11152 30209
rect 11204 30157 11220 30209
rect 11272 30157 11288 30209
rect 11340 30157 11341 30209
rect 6376 30144 11341 30157
rect 4900 30094 5600 30118
rect 4900 30092 5195 30094
rect 4290 30079 5195 30092
rect 3060 30027 3514 30038
rect 4290 30027 4712 30079
rect 4764 30027 4780 30079
rect 4832 30027 4848 30079
rect 4900 30038 5195 30079
rect 5251 30038 5276 30094
rect 5332 30038 5357 30094
rect 5413 30038 5438 30094
rect 5494 30038 5519 30094
rect 5575 30038 5600 30094
rect 6376 30092 6552 30144
rect 6604 30092 6620 30144
rect 6672 30092 6688 30144
rect 6740 30092 7472 30144
rect 7524 30092 7540 30144
rect 7592 30092 7608 30144
rect 7660 30092 8392 30144
rect 8444 30092 8460 30144
rect 8512 30092 8528 30144
rect 8580 30092 9312 30144
rect 9364 30092 9380 30144
rect 9432 30092 9448 30144
rect 9500 30092 10232 30144
rect 10284 30092 10300 30144
rect 10352 30092 10368 30144
rect 10420 30092 11152 30144
rect 11204 30092 11220 30144
rect 11272 30092 11288 30144
rect 11340 30092 11341 30144
rect 6376 30079 11341 30092
rect 4900 30027 5600 30038
rect 6376 30027 6552 30079
rect 6604 30027 6620 30079
rect 6672 30027 6688 30079
rect 6740 30027 7472 30079
rect 7524 30027 7540 30079
rect 7592 30027 7608 30079
rect 7660 30027 8392 30079
rect 8444 30027 8460 30079
rect 8512 30027 8528 30079
rect 8580 30027 9312 30079
rect 9364 30027 9380 30079
rect 9432 30027 9448 30079
rect 9500 30027 10232 30079
rect 10284 30027 10300 30079
rect 10352 30027 10368 30079
rect 10420 30027 11152 30079
rect 11204 30027 11220 30079
rect 11272 30027 11288 30079
rect 11340 30027 11341 30079
rect 187 30014 3514 30027
rect 4290 30014 5600 30027
rect 6376 30014 11341 30027
rect 187 29962 2872 30014
rect 2924 29962 2940 30014
rect 2992 29962 3008 30014
rect 3060 29962 3109 30014
rect 187 29958 3109 29962
rect 3165 29958 3190 30014
rect 3246 29958 3271 30014
rect 3327 29958 3352 30014
rect 3408 29958 3433 30014
rect 3489 29958 3514 30014
rect 4290 29962 4712 30014
rect 4764 29962 4780 30014
rect 4832 29962 4848 30014
rect 4900 29962 5195 30014
rect 4290 29958 5195 29962
rect 5251 29958 5276 30014
rect 5332 29958 5357 30014
rect 5413 29958 5438 30014
rect 5494 29958 5519 30014
rect 5575 29958 5600 30014
rect 6376 29962 6552 30014
rect 6604 29962 6620 30014
rect 6672 29962 6688 30014
rect 6740 29962 7472 30014
rect 7524 29962 7540 30014
rect 7592 29962 7608 30014
rect 7660 29962 8392 30014
rect 8444 29962 8460 30014
rect 8512 29962 8528 30014
rect 8580 29962 9312 30014
rect 9364 29962 9380 30014
rect 9432 29962 9448 30014
rect 9500 29962 10232 30014
rect 10284 29962 10300 30014
rect 10352 29962 10368 30014
rect 10420 29962 11152 30014
rect 11204 29962 11220 30014
rect 11272 29962 11288 30014
rect 11340 29962 11341 30014
rect 6376 29958 11341 29962
rect 187 29956 11341 29958
rect 187 29775 3356 29956
tri 3356 29775 3537 29956 nw
rect 187 27096 2824 29775
tri 2824 29243 3356 29775 nw
tri 11497 29631 12222 30356 se
rect 12222 29631 14858 32491
tri 3361 29342 3650 29631 se
rect 3650 29629 14858 29631
rect 3650 29625 8580 29629
rect 3650 29573 4281 29625
rect 4333 29573 4359 29625
rect 4411 29573 5201 29625
rect 5253 29573 5279 29625
rect 5331 29573 6121 29625
rect 6173 29573 6199 29625
rect 6251 29573 7041 29625
rect 7093 29573 7119 29625
rect 7171 29573 7961 29625
rect 8013 29573 8039 29625
rect 8091 29573 8580 29625
rect 8636 29573 8661 29629
rect 8717 29573 8742 29629
rect 8798 29573 8823 29629
rect 8879 29625 8904 29629
rect 8960 29625 8985 29629
rect 8879 29573 8881 29625
rect 9041 29573 9066 29629
rect 3650 29561 9066 29573
rect 3650 29509 4281 29561
rect 4333 29509 4359 29561
rect 4411 29509 5201 29561
rect 5253 29509 5279 29561
rect 5331 29509 6121 29561
rect 6173 29509 6199 29561
rect 6251 29509 7041 29561
rect 7093 29509 7119 29561
rect 7171 29509 7961 29561
rect 8013 29509 8039 29561
rect 8091 29549 8881 29561
rect 8933 29549 8959 29561
rect 9011 29549 9066 29561
rect 8091 29509 8580 29549
rect 3650 29497 8580 29509
rect 3650 29445 4281 29497
rect 4333 29445 4359 29497
rect 4411 29445 5201 29497
rect 5253 29445 5279 29497
rect 5331 29445 6121 29497
rect 6173 29445 6199 29497
rect 6251 29445 7041 29497
rect 7093 29445 7119 29497
rect 7171 29445 7961 29497
rect 8013 29445 8039 29497
rect 8091 29493 8580 29497
rect 8636 29493 8661 29549
rect 8717 29493 8742 29549
rect 8798 29493 8823 29549
rect 8879 29509 8881 29549
rect 8879 29497 8904 29509
rect 8960 29497 8985 29509
rect 8879 29493 8881 29497
rect 9041 29493 9066 29549
rect 8091 29469 8881 29493
rect 8933 29469 8959 29493
rect 9011 29469 9066 29493
rect 8091 29445 8580 29469
rect 3650 29433 8580 29445
rect 3650 29381 4281 29433
rect 4333 29381 4359 29433
rect 4411 29381 5201 29433
rect 5253 29381 5279 29433
rect 5331 29381 6121 29433
rect 6173 29381 6199 29433
rect 6251 29381 7041 29433
rect 7093 29381 7119 29433
rect 7171 29381 7961 29433
rect 8013 29381 8039 29433
rect 8091 29413 8580 29433
rect 8636 29413 8661 29469
rect 8717 29413 8742 29469
rect 8798 29413 8823 29469
rect 8879 29445 8881 29469
rect 8879 29433 8904 29445
rect 8960 29433 8985 29445
rect 8879 29413 8881 29433
rect 9041 29413 9066 29469
rect 8091 29389 8881 29413
rect 8933 29389 8959 29413
rect 9011 29389 9066 29413
rect 8091 29381 8580 29389
rect 3650 29369 8580 29381
rect 3650 29342 4281 29369
rect 3361 29336 4281 29342
rect 3413 29284 3439 29336
rect 3491 29317 4281 29336
rect 4333 29317 4359 29369
rect 4411 29317 5201 29369
rect 5253 29317 5279 29369
rect 5331 29317 6121 29369
rect 6173 29317 6199 29369
rect 6251 29317 7041 29369
rect 7093 29317 7119 29369
rect 7171 29317 7961 29369
rect 8013 29317 8039 29369
rect 8091 29333 8580 29369
rect 8636 29333 8661 29389
rect 8717 29333 8742 29389
rect 8798 29333 8823 29389
rect 8879 29381 8881 29389
rect 8879 29369 8904 29381
rect 8960 29369 8985 29381
rect 8879 29333 8881 29369
rect 9041 29333 9066 29389
rect 8091 29317 8881 29333
rect 8933 29317 8959 29333
rect 9011 29317 9066 29333
rect 3491 29309 9066 29317
rect 3491 29305 8580 29309
rect 3491 29284 4281 29305
rect 3361 29270 4281 29284
rect 3413 29218 3439 29270
rect 3491 29253 4281 29270
rect 4333 29253 4359 29305
rect 4411 29253 5201 29305
rect 5253 29253 5279 29305
rect 5331 29253 6121 29305
rect 6173 29253 6199 29305
rect 6251 29253 7041 29305
rect 7093 29253 7119 29305
rect 7171 29253 7961 29305
rect 8013 29253 8039 29305
rect 8091 29253 8580 29305
rect 8636 29253 8661 29309
rect 8717 29253 8742 29309
rect 8798 29253 8823 29309
rect 8879 29305 8904 29309
rect 8960 29305 8985 29309
rect 8879 29253 8881 29305
rect 9041 29253 9066 29309
rect 3491 29241 9066 29253
rect 3491 29218 4281 29241
rect 3361 29204 4281 29218
rect 3413 29152 3439 29204
rect 3491 29189 4281 29204
rect 4333 29189 4359 29241
rect 4411 29189 5201 29241
rect 5253 29189 5279 29241
rect 5331 29189 6121 29241
rect 6173 29189 6199 29241
rect 6251 29189 7041 29241
rect 7093 29189 7119 29241
rect 7171 29189 7961 29241
rect 8013 29189 8039 29241
rect 8091 29229 8881 29241
rect 8933 29229 8959 29241
rect 9011 29229 9066 29241
rect 8091 29189 8580 29229
rect 3491 29177 8580 29189
rect 3491 29152 4281 29177
rect 3361 29138 4281 29152
rect 3413 29086 3439 29138
rect 3491 29125 4281 29138
rect 4333 29125 4359 29177
rect 4411 29125 5201 29177
rect 5253 29125 5279 29177
rect 5331 29125 6121 29177
rect 6173 29125 6199 29177
rect 6251 29125 7041 29177
rect 7093 29125 7119 29177
rect 7171 29125 7961 29177
rect 8013 29125 8039 29177
rect 8091 29173 8580 29177
rect 8636 29173 8661 29229
rect 8717 29173 8742 29229
rect 8798 29173 8823 29229
rect 8879 29189 8881 29229
rect 8879 29177 8904 29189
rect 8960 29177 8985 29189
rect 8879 29173 8881 29177
rect 9041 29173 9066 29229
rect 8091 29149 8881 29173
rect 8933 29149 8959 29173
rect 9011 29149 9066 29173
rect 8091 29125 8580 29149
rect 3491 29113 8580 29125
rect 3491 29086 4281 29113
rect 3361 29072 4281 29086
rect 3413 29020 3439 29072
rect 3491 29061 4281 29072
rect 4333 29061 4359 29113
rect 4411 29061 5201 29113
rect 5253 29061 5279 29113
rect 5331 29061 6121 29113
rect 6173 29061 6199 29113
rect 6251 29061 7041 29113
rect 7093 29061 7119 29113
rect 7171 29061 7961 29113
rect 8013 29061 8039 29113
rect 8091 29093 8580 29113
rect 8636 29093 8661 29149
rect 8717 29093 8742 29149
rect 8798 29093 8823 29149
rect 8879 29125 8881 29149
rect 8879 29113 8904 29125
rect 8960 29113 8985 29125
rect 8879 29093 8881 29113
rect 9041 29093 9066 29149
rect 8091 29069 8881 29093
rect 8933 29069 8959 29093
rect 9011 29069 9066 29093
rect 8091 29061 8580 29069
rect 3491 29049 8580 29061
rect 3491 29020 4281 29049
rect 3361 29006 4281 29020
rect 3413 28954 3439 29006
rect 3491 28997 4281 29006
rect 4333 28997 4359 29049
rect 4411 28997 5201 29049
rect 5253 28997 5279 29049
rect 5331 28997 6121 29049
rect 6173 28997 6199 29049
rect 6251 28997 7041 29049
rect 7093 28997 7119 29049
rect 7171 28997 7961 29049
rect 8013 28997 8039 29049
rect 8091 29013 8580 29049
rect 8636 29013 8661 29069
rect 8717 29013 8742 29069
rect 8798 29013 8823 29069
rect 8879 29061 8881 29069
rect 8879 29049 8904 29061
rect 8960 29049 8985 29061
rect 8879 29013 8881 29049
rect 9041 29013 9066 29069
rect 8091 28997 8881 29013
rect 8933 28997 8959 29013
rect 9011 28997 9066 29013
rect 3491 28989 9066 28997
rect 3491 28985 8580 28989
rect 3491 28954 4281 28985
rect 3361 28940 4281 28954
rect 3413 28888 3439 28940
rect 3491 28933 4281 28940
rect 4333 28933 4359 28985
rect 4411 28933 5201 28985
rect 5253 28933 5279 28985
rect 5331 28933 6121 28985
rect 6173 28933 6199 28985
rect 6251 28933 7041 28985
rect 7093 28933 7119 28985
rect 7171 28933 7961 28985
rect 8013 28933 8039 28985
rect 8091 28933 8580 28985
rect 8636 28933 8661 28989
rect 8717 28933 8742 28989
rect 8798 28933 8823 28989
rect 8879 28985 8904 28989
rect 8960 28985 8985 28989
rect 8879 28933 8881 28985
rect 9041 28933 9066 28989
rect 3491 28921 9066 28933
rect 3491 28888 4281 28921
rect 3361 28874 4281 28888
rect 3413 28822 3439 28874
rect 3491 28869 4281 28874
rect 4333 28869 4359 28921
rect 4411 28869 5201 28921
rect 5253 28869 5279 28921
rect 5331 28869 6121 28921
rect 6173 28869 6199 28921
rect 6251 28869 7041 28921
rect 7093 28869 7119 28921
rect 7171 28869 7961 28921
rect 8013 28869 8039 28921
rect 8091 28909 8881 28921
rect 8933 28909 8959 28921
rect 9011 28909 9066 28921
rect 8091 28869 8580 28909
rect 3491 28857 8580 28869
rect 3491 28822 4281 28857
rect 3361 28808 4281 28822
rect 3413 28756 3439 28808
rect 3491 28805 4281 28808
rect 4333 28805 4359 28857
rect 4411 28805 5201 28857
rect 5253 28805 5279 28857
rect 5331 28805 6121 28857
rect 6173 28805 6199 28857
rect 6251 28805 7041 28857
rect 7093 28805 7119 28857
rect 7171 28805 7961 28857
rect 8013 28805 8039 28857
rect 8091 28853 8580 28857
rect 8636 28853 8661 28909
rect 8717 28853 8742 28909
rect 8798 28853 8823 28909
rect 8879 28869 8881 28909
rect 8879 28857 8904 28869
rect 8960 28857 8985 28869
rect 8879 28853 8881 28857
rect 9041 28853 9066 28909
rect 8091 28829 8881 28853
rect 8933 28829 8959 28853
rect 9011 28829 9066 28853
rect 8091 28805 8580 28829
rect 3491 28793 8580 28805
rect 3491 28756 4281 28793
rect 3361 28742 4281 28756
rect 3413 28690 3439 28742
rect 3491 28741 4281 28742
rect 4333 28741 4359 28793
rect 4411 28741 5201 28793
rect 5253 28741 5279 28793
rect 5331 28741 6121 28793
rect 6173 28741 6199 28793
rect 6251 28741 7041 28793
rect 7093 28741 7119 28793
rect 7171 28741 7961 28793
rect 8013 28741 8039 28793
rect 8091 28773 8580 28793
rect 8636 28773 8661 28829
rect 8717 28773 8742 28829
rect 8798 28773 8823 28829
rect 8879 28805 8881 28829
rect 8879 28793 8904 28805
rect 8960 28793 8985 28805
rect 8879 28773 8881 28793
rect 9041 28773 9066 28829
rect 8091 28749 8881 28773
rect 8933 28749 8959 28773
rect 9011 28749 9066 28773
rect 8091 28741 8580 28749
rect 3491 28729 8580 28741
rect 3491 28690 4281 28729
rect 3361 28677 4281 28690
rect 4333 28677 4359 28729
rect 4411 28677 5201 28729
rect 5253 28677 5279 28729
rect 5331 28677 6121 28729
rect 6173 28677 6199 28729
rect 6251 28677 7041 28729
rect 7093 28677 7119 28729
rect 7171 28677 7961 28729
rect 8013 28677 8039 28729
rect 8091 28693 8580 28729
rect 8636 28693 8661 28749
rect 8717 28693 8742 28749
rect 8798 28693 8823 28749
rect 8879 28741 8881 28749
rect 8879 28729 8904 28741
rect 8960 28729 8985 28741
rect 8879 28693 8881 28729
rect 9041 28693 9066 28749
rect 8091 28677 8881 28693
rect 8933 28677 8959 28693
rect 9011 28677 9066 28693
rect 3361 28676 9066 28677
rect 3413 28624 3439 28676
rect 3491 28669 9066 28676
rect 3491 28664 8580 28669
rect 3491 28624 4281 28664
rect 3361 28612 4281 28624
rect 4333 28612 4359 28664
rect 4411 28612 5201 28664
rect 5253 28612 5279 28664
rect 5331 28612 6121 28664
rect 6173 28612 6199 28664
rect 6251 28612 7041 28664
rect 7093 28612 7119 28664
rect 7171 28612 7961 28664
rect 8013 28612 8039 28664
rect 8091 28613 8580 28664
rect 8636 28613 8661 28669
rect 8717 28613 8742 28669
rect 8798 28613 8823 28669
rect 8879 28664 8904 28669
rect 8960 28664 8985 28669
rect 8879 28613 8881 28664
rect 9041 28613 9066 28669
rect 8091 28612 8881 28613
rect 8933 28612 8959 28613
rect 9011 28612 9066 28613
rect 3361 28610 9066 28612
rect 3413 28558 3439 28610
rect 3491 28599 9066 28610
rect 3491 28558 4281 28599
rect 3361 28547 4281 28558
rect 4333 28547 4359 28599
rect 4411 28547 5201 28599
rect 5253 28547 5279 28599
rect 5331 28547 6121 28599
rect 6173 28547 6199 28599
rect 6251 28547 7041 28599
rect 7093 28547 7119 28599
rect 7171 28547 7961 28599
rect 8013 28547 8039 28599
rect 8091 28589 8881 28599
rect 8933 28589 8959 28599
rect 9011 28589 9066 28599
rect 8091 28547 8580 28589
rect 3361 28544 8580 28547
rect 3413 28492 3439 28544
rect 3491 28534 8580 28544
rect 3491 28492 4281 28534
rect 3361 28482 4281 28492
rect 4333 28482 4359 28534
rect 4411 28482 5201 28534
rect 5253 28482 5279 28534
rect 5331 28482 6121 28534
rect 6173 28482 6199 28534
rect 6251 28482 7041 28534
rect 7093 28482 7119 28534
rect 7171 28482 7961 28534
rect 8013 28482 8039 28534
rect 8091 28533 8580 28534
rect 8636 28533 8661 28589
rect 8717 28533 8742 28589
rect 8798 28533 8823 28589
rect 8879 28547 8881 28589
rect 8879 28534 8904 28547
rect 8960 28534 8985 28547
rect 8879 28533 8881 28534
rect 9041 28533 9066 28589
rect 8091 28509 8881 28533
rect 8933 28509 8959 28533
rect 9011 28509 9066 28533
rect 8091 28482 8580 28509
rect 3361 28478 8580 28482
rect 3413 28426 3439 28478
rect 3491 28469 8580 28478
rect 3491 28426 4281 28469
rect 3361 28417 4281 28426
rect 4333 28417 4359 28469
rect 4411 28417 5201 28469
rect 5253 28417 5279 28469
rect 5331 28417 6121 28469
rect 6173 28417 6199 28469
rect 6251 28417 7041 28469
rect 7093 28417 7119 28469
rect 7171 28417 7961 28469
rect 8013 28417 8039 28469
rect 8091 28453 8580 28469
rect 8636 28453 8661 28509
rect 8717 28453 8742 28509
rect 8798 28453 8823 28509
rect 8879 28482 8881 28509
rect 8879 28469 8904 28482
rect 8960 28469 8985 28482
rect 8879 28453 8881 28469
rect 9041 28453 9066 28509
rect 8091 28429 8881 28453
rect 8933 28429 8959 28453
rect 9011 28429 9066 28453
rect 8091 28417 8580 28429
rect 3361 28412 8580 28417
rect 3413 28360 3439 28412
rect 3491 28404 8580 28412
rect 3491 28360 4281 28404
rect 3361 28352 4281 28360
rect 4333 28352 4359 28404
rect 4411 28352 5201 28404
rect 5253 28352 5279 28404
rect 5331 28352 6121 28404
rect 6173 28352 6199 28404
rect 6251 28352 7041 28404
rect 7093 28352 7119 28404
rect 7171 28352 7961 28404
rect 8013 28352 8039 28404
rect 8091 28373 8580 28404
rect 8636 28373 8661 28429
rect 8717 28373 8742 28429
rect 8798 28373 8823 28429
rect 8879 28417 8881 28429
rect 8879 28404 8904 28417
rect 8960 28404 8985 28417
rect 8879 28373 8881 28404
rect 9041 28373 9066 28429
rect 8091 28352 8881 28373
rect 8933 28352 8959 28373
rect 9011 28352 9066 28373
rect 3361 28349 9066 28352
rect 3361 28346 8580 28349
rect 3413 28294 3439 28346
rect 3491 28339 8580 28346
rect 3491 28294 4281 28339
rect 3361 28287 4281 28294
rect 4333 28287 4359 28339
rect 4411 28287 5201 28339
rect 5253 28287 5279 28339
rect 5331 28287 6121 28339
rect 6173 28287 6199 28339
rect 6251 28287 7041 28339
rect 7093 28287 7119 28339
rect 7171 28287 7961 28339
rect 8013 28287 8039 28339
rect 8091 28293 8580 28339
rect 8636 28293 8661 28349
rect 8717 28293 8742 28349
rect 8798 28293 8823 28349
rect 8879 28339 8904 28349
rect 8960 28339 8985 28349
rect 8879 28293 8881 28339
rect 9041 28293 9066 28349
rect 8091 28287 8881 28293
rect 8933 28287 8959 28293
rect 9011 28287 9066 28293
rect 3361 28280 9066 28287
rect 3413 28228 3439 28280
rect 3491 28274 9066 28280
rect 3491 28228 4281 28274
rect 3361 28222 4281 28228
rect 4333 28222 4359 28274
rect 4411 28222 5201 28274
rect 5253 28222 5279 28274
rect 5331 28222 6121 28274
rect 6173 28222 6199 28274
rect 6251 28222 7041 28274
rect 7093 28222 7119 28274
rect 7171 28222 7961 28274
rect 8013 28222 8039 28274
rect 8091 28269 8881 28274
rect 8933 28269 8959 28274
rect 9011 28269 9066 28274
rect 8091 28222 8580 28269
rect 3361 28214 8580 28222
rect 3413 28162 3439 28214
rect 3491 28213 8580 28214
rect 8636 28213 8661 28269
rect 8717 28213 8742 28269
rect 8798 28213 8823 28269
rect 8879 28222 8881 28269
rect 8879 28213 8904 28222
rect 8960 28213 8985 28222
rect 9041 28213 9066 28269
rect 3491 28209 9066 28213
rect 3491 28162 4281 28209
rect 3361 28157 4281 28162
rect 4333 28157 4359 28209
rect 4411 28157 5201 28209
rect 5253 28157 5279 28209
rect 5331 28157 6121 28209
rect 6173 28157 6199 28209
rect 6251 28157 7041 28209
rect 7093 28157 7119 28209
rect 7171 28157 7961 28209
rect 8013 28157 8039 28209
rect 8091 28189 8881 28209
rect 8933 28189 8959 28209
rect 9011 28189 9066 28209
rect 8091 28157 8580 28189
rect 3361 28148 8580 28157
rect 3413 28096 3439 28148
rect 3491 28144 8580 28148
rect 3491 28096 4281 28144
rect 3361 28092 4281 28096
rect 4333 28092 4359 28144
rect 4411 28092 5201 28144
rect 5253 28092 5279 28144
rect 5331 28092 6121 28144
rect 6173 28092 6199 28144
rect 6251 28092 7041 28144
rect 7093 28092 7119 28144
rect 7171 28092 7961 28144
rect 8013 28092 8039 28144
rect 8091 28133 8580 28144
rect 8636 28133 8661 28189
rect 8717 28133 8742 28189
rect 8798 28133 8823 28189
rect 8879 28157 8881 28189
rect 8879 28144 8904 28157
rect 8960 28144 8985 28157
rect 8879 28133 8881 28144
rect 9041 28133 9066 28189
rect 8091 28109 8881 28133
rect 8933 28109 8959 28133
rect 9011 28109 9066 28133
rect 8091 28092 8580 28109
rect 3361 28082 8580 28092
rect 3413 28030 3439 28082
rect 3491 28079 8580 28082
rect 3491 28030 4281 28079
rect 3361 28027 4281 28030
rect 4333 28027 4359 28079
rect 4411 28027 5201 28079
rect 5253 28027 5279 28079
rect 5331 28027 6121 28079
rect 6173 28027 6199 28079
rect 6251 28027 7041 28079
rect 7093 28027 7119 28079
rect 7171 28027 7961 28079
rect 8013 28027 8039 28079
rect 8091 28053 8580 28079
rect 8636 28053 8661 28109
rect 8717 28053 8742 28109
rect 8798 28053 8823 28109
rect 8879 28092 8881 28109
rect 8879 28079 8904 28092
rect 8960 28079 8985 28092
rect 8879 28053 8881 28079
rect 9041 28053 9066 28109
rect 8091 28029 8881 28053
rect 8933 28029 8959 28053
rect 9011 28029 9066 28053
rect 8091 28027 8580 28029
rect 3361 28016 8580 28027
rect 3413 27964 3439 28016
rect 3491 28014 8580 28016
rect 3491 27964 4281 28014
rect 3361 27962 4281 27964
rect 4333 27962 4359 28014
rect 4411 27962 5201 28014
rect 5253 27962 5279 28014
rect 5331 27962 6121 28014
rect 6173 27962 6199 28014
rect 6251 27962 7041 28014
rect 7093 27962 7119 28014
rect 7171 27962 7961 28014
rect 8013 27962 8039 28014
rect 8091 27973 8580 28014
rect 8636 27973 8661 28029
rect 8717 27973 8742 28029
rect 8798 27973 8823 28029
rect 8879 28027 8881 28029
rect 8879 28014 8904 28027
rect 8960 28014 8985 28027
rect 8879 27973 8881 28014
rect 9041 27973 9066 28029
rect 8091 27962 8881 27973
rect 8933 27962 8959 27973
rect 9011 27962 9066 27973
rect 3361 27949 9066 27962
rect 3413 27897 3439 27949
rect 3491 27897 4281 27949
rect 4333 27897 4359 27949
rect 4411 27897 5201 27949
rect 5253 27897 5279 27949
rect 5331 27897 6121 27949
rect 6173 27897 6199 27949
rect 6251 27897 7041 27949
rect 7093 27897 7119 27949
rect 7171 27897 7961 27949
rect 8013 27897 8039 27949
rect 8091 27897 8580 27949
rect 3361 27893 8580 27897
rect 8636 27893 8661 27949
rect 8717 27893 8742 27949
rect 8798 27893 8823 27949
rect 8879 27897 8881 27949
rect 8879 27893 8904 27897
rect 8960 27893 8985 27897
rect 9041 27893 9066 27949
rect 9762 29625 10666 29629
rect 10722 29625 10747 29629
rect 10803 29625 10828 29629
rect 9762 29573 9801 29625
rect 9853 29573 9879 29625
rect 9931 29573 10666 29625
rect 10884 29573 10909 29629
rect 10965 29573 10990 29629
rect 11046 29573 11071 29629
rect 11127 29573 11152 29629
rect 11848 29625 14858 29629
rect 11848 29573 12561 29625
rect 12613 29573 12639 29625
rect 12691 29573 14858 29625
rect 9762 29561 11152 29573
rect 11848 29561 14858 29573
rect 9762 29509 9801 29561
rect 9853 29509 9879 29561
rect 9931 29549 10721 29561
rect 10773 29549 10799 29561
rect 10851 29549 11152 29561
rect 9931 29509 10666 29549
rect 9762 29497 10666 29509
rect 10722 29497 10747 29509
rect 10803 29497 10828 29509
rect 9762 29445 9801 29497
rect 9853 29445 9879 29497
rect 9931 29493 10666 29497
rect 10884 29493 10909 29549
rect 10965 29493 10990 29549
rect 11046 29493 11071 29549
rect 11127 29493 11152 29549
rect 11848 29509 12561 29561
rect 12613 29509 12639 29561
rect 12691 29509 14858 29561
rect 11848 29497 14858 29509
rect 9931 29469 10721 29493
rect 10773 29469 10799 29493
rect 10851 29469 11152 29493
rect 9931 29445 10666 29469
rect 9762 29433 10666 29445
rect 10722 29433 10747 29445
rect 10803 29433 10828 29445
rect 9762 29381 9801 29433
rect 9853 29381 9879 29433
rect 9931 29413 10666 29433
rect 10884 29413 10909 29469
rect 10965 29413 10990 29469
rect 11046 29413 11071 29469
rect 11127 29413 11152 29469
rect 11848 29445 12561 29497
rect 12613 29445 12639 29497
rect 12691 29445 14858 29497
rect 11848 29433 14858 29445
rect 9931 29389 10721 29413
rect 10773 29389 10799 29413
rect 10851 29389 11152 29413
rect 9931 29381 10666 29389
rect 9762 29369 10666 29381
rect 10722 29369 10747 29381
rect 10803 29369 10828 29381
rect 9762 29317 9801 29369
rect 9853 29317 9879 29369
rect 9931 29333 10666 29369
rect 10884 29333 10909 29389
rect 10965 29333 10990 29389
rect 11046 29333 11071 29389
rect 11127 29333 11152 29389
rect 11848 29381 12561 29433
rect 12613 29381 12639 29433
rect 12691 29381 14858 29433
rect 11848 29369 14858 29381
rect 9931 29317 10721 29333
rect 10773 29317 10799 29333
rect 10851 29317 11152 29333
rect 11848 29317 12561 29369
rect 12613 29317 12639 29369
rect 12691 29317 14858 29369
rect 9762 29309 11152 29317
rect 9762 29305 10666 29309
rect 10722 29305 10747 29309
rect 10803 29305 10828 29309
rect 9762 29253 9801 29305
rect 9853 29253 9879 29305
rect 9931 29253 10666 29305
rect 10884 29253 10909 29309
rect 10965 29253 10990 29309
rect 11046 29253 11071 29309
rect 11127 29253 11152 29309
rect 11848 29305 14858 29317
rect 11848 29253 12561 29305
rect 12613 29253 12639 29305
rect 12691 29253 14858 29305
rect 9762 29241 11152 29253
rect 11848 29241 14858 29253
rect 9762 29189 9801 29241
rect 9853 29189 9879 29241
rect 9931 29229 10721 29241
rect 10773 29229 10799 29241
rect 10851 29229 11152 29241
rect 9931 29189 10666 29229
rect 9762 29177 10666 29189
rect 10722 29177 10747 29189
rect 10803 29177 10828 29189
rect 9762 29125 9801 29177
rect 9853 29125 9879 29177
rect 9931 29173 10666 29177
rect 10884 29173 10909 29229
rect 10965 29173 10990 29229
rect 11046 29173 11071 29229
rect 11127 29173 11152 29229
rect 11848 29189 12561 29241
rect 12613 29189 12639 29241
rect 12691 29189 14858 29241
rect 11848 29177 14858 29189
rect 9931 29149 10721 29173
rect 10773 29149 10799 29173
rect 10851 29149 11152 29173
rect 9931 29125 10666 29149
rect 9762 29113 10666 29125
rect 10722 29113 10747 29125
rect 10803 29113 10828 29125
rect 9762 29061 9801 29113
rect 9853 29061 9879 29113
rect 9931 29093 10666 29113
rect 10884 29093 10909 29149
rect 10965 29093 10990 29149
rect 11046 29093 11071 29149
rect 11127 29093 11152 29149
rect 11848 29125 12561 29177
rect 12613 29125 12639 29177
rect 12691 29125 14858 29177
rect 11848 29113 14858 29125
rect 9931 29069 10721 29093
rect 10773 29069 10799 29093
rect 10851 29069 11152 29093
rect 9931 29061 10666 29069
rect 9762 29049 10666 29061
rect 10722 29049 10747 29061
rect 10803 29049 10828 29061
rect 9762 28997 9801 29049
rect 9853 28997 9879 29049
rect 9931 29013 10666 29049
rect 10884 29013 10909 29069
rect 10965 29013 10990 29069
rect 11046 29013 11071 29069
rect 11127 29013 11152 29069
rect 11848 29061 12561 29113
rect 12613 29061 12639 29113
rect 12691 29061 14858 29113
rect 11848 29049 14858 29061
rect 9931 28997 10721 29013
rect 10773 28997 10799 29013
rect 10851 28997 11152 29013
rect 11848 28997 12561 29049
rect 12613 28997 12639 29049
rect 12691 28997 14858 29049
rect 9762 28989 11152 28997
rect 9762 28985 10666 28989
rect 10722 28985 10747 28989
rect 10803 28985 10828 28989
rect 9762 28933 9801 28985
rect 9853 28933 9879 28985
rect 9931 28933 10666 28985
rect 10884 28933 10909 28989
rect 10965 28933 10990 28989
rect 11046 28933 11071 28989
rect 11127 28933 11152 28989
rect 11848 28985 14858 28997
rect 11848 28933 12561 28985
rect 12613 28933 12639 28985
rect 12691 28933 14858 28985
rect 9762 28921 11152 28933
rect 11848 28921 14858 28933
rect 9762 28869 9801 28921
rect 9853 28869 9879 28921
rect 9931 28909 10721 28921
rect 10773 28909 10799 28921
rect 10851 28909 11152 28921
rect 9931 28869 10666 28909
rect 9762 28857 10666 28869
rect 10722 28857 10747 28869
rect 10803 28857 10828 28869
rect 9762 28805 9801 28857
rect 9853 28805 9879 28857
rect 9931 28853 10666 28857
rect 10884 28853 10909 28909
rect 10965 28853 10990 28909
rect 11046 28853 11071 28909
rect 11127 28853 11152 28909
rect 11848 28869 12561 28921
rect 12613 28869 12639 28921
rect 12691 28869 14858 28921
rect 11848 28857 14858 28869
rect 9931 28829 10721 28853
rect 10773 28829 10799 28853
rect 10851 28829 11152 28853
rect 9931 28805 10666 28829
rect 9762 28793 10666 28805
rect 10722 28793 10747 28805
rect 10803 28793 10828 28805
rect 9762 28741 9801 28793
rect 9853 28741 9879 28793
rect 9931 28773 10666 28793
rect 10884 28773 10909 28829
rect 10965 28773 10990 28829
rect 11046 28773 11071 28829
rect 11127 28773 11152 28829
rect 11848 28805 12561 28857
rect 12613 28805 12639 28857
rect 12691 28805 14858 28857
rect 11848 28793 14858 28805
rect 9931 28749 10721 28773
rect 10773 28749 10799 28773
rect 10851 28749 11152 28773
rect 9931 28741 10666 28749
rect 9762 28729 10666 28741
rect 10722 28729 10747 28741
rect 10803 28729 10828 28741
rect 9762 28677 9801 28729
rect 9853 28677 9879 28729
rect 9931 28693 10666 28729
rect 10884 28693 10909 28749
rect 10965 28693 10990 28749
rect 11046 28693 11071 28749
rect 11127 28693 11152 28749
rect 11848 28741 12561 28793
rect 12613 28741 12639 28793
rect 12691 28741 14858 28793
rect 11848 28729 14858 28741
rect 9931 28677 10721 28693
rect 10773 28677 10799 28693
rect 10851 28677 11152 28693
rect 11848 28677 12561 28729
rect 12613 28677 12639 28729
rect 12691 28677 14858 28729
rect 9762 28669 11152 28677
rect 9762 28664 10666 28669
rect 10722 28664 10747 28669
rect 10803 28664 10828 28669
rect 9762 28612 9801 28664
rect 9853 28612 9879 28664
rect 9931 28613 10666 28664
rect 10884 28613 10909 28669
rect 10965 28613 10990 28669
rect 11046 28613 11071 28669
rect 11127 28613 11152 28669
rect 11848 28664 14858 28677
rect 9931 28612 10721 28613
rect 10773 28612 10799 28613
rect 10851 28612 11152 28613
rect 11848 28612 12561 28664
rect 12613 28612 12639 28664
rect 12691 28612 14858 28664
rect 9762 28599 11152 28612
rect 11848 28599 14858 28612
rect 9762 28547 9801 28599
rect 9853 28547 9879 28599
rect 9931 28589 10721 28599
rect 10773 28589 10799 28599
rect 10851 28589 11152 28599
rect 9931 28547 10666 28589
rect 9762 28534 10666 28547
rect 10722 28534 10747 28547
rect 10803 28534 10828 28547
rect 9762 28482 9801 28534
rect 9853 28482 9879 28534
rect 9931 28533 10666 28534
rect 10884 28533 10909 28589
rect 10965 28533 10990 28589
rect 11046 28533 11071 28589
rect 11127 28533 11152 28589
rect 11848 28547 12561 28599
rect 12613 28547 12639 28599
rect 12691 28547 14858 28599
rect 11848 28534 14858 28547
rect 9931 28509 10721 28533
rect 10773 28509 10799 28533
rect 10851 28509 11152 28533
rect 9931 28482 10666 28509
rect 9762 28469 10666 28482
rect 10722 28469 10747 28482
rect 10803 28469 10828 28482
rect 9762 28417 9801 28469
rect 9853 28417 9879 28469
rect 9931 28453 10666 28469
rect 10884 28453 10909 28509
rect 10965 28453 10990 28509
rect 11046 28453 11071 28509
rect 11127 28453 11152 28509
rect 11848 28482 12561 28534
rect 12613 28482 12639 28534
rect 12691 28482 14858 28534
rect 11848 28469 14858 28482
rect 9931 28429 10721 28453
rect 10773 28429 10799 28453
rect 10851 28429 11152 28453
rect 9931 28417 10666 28429
rect 9762 28404 10666 28417
rect 10722 28404 10747 28417
rect 10803 28404 10828 28417
rect 9762 28352 9801 28404
rect 9853 28352 9879 28404
rect 9931 28373 10666 28404
rect 10884 28373 10909 28429
rect 10965 28373 10990 28429
rect 11046 28373 11071 28429
rect 11127 28373 11152 28429
rect 11848 28417 12561 28469
rect 12613 28417 12639 28469
rect 12691 28417 14858 28469
rect 11848 28404 14858 28417
rect 9931 28352 10721 28373
rect 10773 28352 10799 28373
rect 10851 28352 11152 28373
rect 11848 28352 12561 28404
rect 12613 28352 12639 28404
rect 12691 28352 14858 28404
rect 9762 28349 11152 28352
rect 9762 28339 10666 28349
rect 10722 28339 10747 28349
rect 10803 28339 10828 28349
rect 9762 28287 9801 28339
rect 9853 28287 9879 28339
rect 9931 28293 10666 28339
rect 10884 28293 10909 28349
rect 10965 28293 10990 28349
rect 11046 28293 11071 28349
rect 11127 28293 11152 28349
rect 11848 28339 14858 28352
rect 9931 28287 10721 28293
rect 10773 28287 10799 28293
rect 10851 28287 11152 28293
rect 11848 28287 12561 28339
rect 12613 28287 12639 28339
rect 12691 28287 14858 28339
rect 9762 28274 11152 28287
rect 11848 28274 14858 28287
rect 9762 28222 9801 28274
rect 9853 28222 9879 28274
rect 9931 28269 10721 28274
rect 10773 28269 10799 28274
rect 10851 28269 11152 28274
rect 9931 28222 10666 28269
rect 9762 28213 10666 28222
rect 10722 28213 10747 28222
rect 10803 28213 10828 28222
rect 10884 28213 10909 28269
rect 10965 28213 10990 28269
rect 11046 28213 11071 28269
rect 11127 28213 11152 28269
rect 11848 28222 12561 28274
rect 12613 28222 12639 28274
rect 12691 28222 14858 28274
rect 9762 28209 11152 28213
rect 11848 28209 14858 28222
rect 9762 28157 9801 28209
rect 9853 28157 9879 28209
rect 9931 28189 10721 28209
rect 10773 28189 10799 28209
rect 10851 28189 11152 28209
rect 9931 28157 10666 28189
rect 9762 28144 10666 28157
rect 10722 28144 10747 28157
rect 10803 28144 10828 28157
rect 9762 28092 9801 28144
rect 9853 28092 9879 28144
rect 9931 28133 10666 28144
rect 10884 28133 10909 28189
rect 10965 28133 10990 28189
rect 11046 28133 11071 28189
rect 11127 28133 11152 28189
rect 11848 28157 12561 28209
rect 12613 28157 12639 28209
rect 12691 28157 14858 28209
rect 11848 28144 14858 28157
rect 9931 28109 10721 28133
rect 10773 28109 10799 28133
rect 10851 28109 11152 28133
rect 9931 28092 10666 28109
rect 9762 28079 10666 28092
rect 10722 28079 10747 28092
rect 10803 28079 10828 28092
rect 9762 28027 9801 28079
rect 9853 28027 9879 28079
rect 9931 28053 10666 28079
rect 10884 28053 10909 28109
rect 10965 28053 10990 28109
rect 11046 28053 11071 28109
rect 11127 28053 11152 28109
rect 11848 28092 12561 28144
rect 12613 28092 12639 28144
rect 12691 28092 14858 28144
rect 11848 28079 14858 28092
rect 9931 28029 10721 28053
rect 10773 28029 10799 28053
rect 10851 28029 11152 28053
rect 9931 28027 10666 28029
rect 9762 28014 10666 28027
rect 10722 28014 10747 28027
rect 10803 28014 10828 28027
rect 9762 27962 9801 28014
rect 9853 27962 9879 28014
rect 9931 27973 10666 28014
rect 10884 27973 10909 28029
rect 10965 27973 10990 28029
rect 11046 27973 11071 28029
rect 11127 27973 11152 28029
rect 11848 28027 12561 28079
rect 12613 28027 12639 28079
rect 12691 28027 14858 28079
rect 11848 28014 14858 28027
rect 9931 27962 10721 27973
rect 10773 27962 10799 27973
rect 10851 27962 11152 27973
rect 11848 27962 12561 28014
rect 12613 27962 12639 28014
rect 12691 27962 14858 28014
rect 9762 27949 11152 27962
rect 11848 27949 14858 27962
rect 9762 27897 9801 27949
rect 9853 27897 9879 27949
rect 9931 27897 10666 27949
rect 9762 27893 10666 27897
rect 10722 27893 10747 27897
rect 10803 27893 10828 27897
rect 10884 27893 10909 27949
rect 10965 27893 10990 27949
rect 11046 27893 11071 27949
rect 11127 27893 11152 27949
rect 11848 27897 12561 27949
rect 12613 27897 12639 27949
rect 12691 27897 14858 27949
rect 11848 27893 14858 27897
rect 3361 27891 14858 27893
tri 2824 27096 3562 27834 sw
tri 11502 27171 12222 27891 ne
rect 187 27094 11341 27096
rect 187 27038 3109 27094
rect 3165 27038 3190 27094
rect 3246 27038 3271 27094
rect 3327 27038 3352 27094
rect 3408 27038 3433 27094
rect 3489 27038 3514 27094
rect 187 27014 3514 27038
rect 187 26958 3109 27014
rect 3165 26958 3190 27014
rect 3246 26958 3271 27014
rect 3327 26958 3352 27014
rect 3408 26958 3433 27014
rect 3489 26958 3514 27014
rect 187 26934 3514 26958
rect 187 26878 3109 26934
rect 3165 26878 3190 26934
rect 3246 26878 3271 26934
rect 3327 26878 3352 26934
rect 3408 26878 3433 26934
rect 3489 26878 3514 26934
rect 187 26854 3514 26878
rect 187 26798 3109 26854
rect 3165 26798 3190 26854
rect 3246 26798 3271 26854
rect 3327 26798 3352 26854
rect 3408 26798 3433 26854
rect 3489 26798 3514 26854
rect 187 26774 3514 26798
rect 187 26718 3109 26774
rect 3165 26718 3190 26774
rect 3246 26718 3271 26774
rect 3327 26718 3352 26774
rect 3408 26718 3433 26774
rect 3489 26718 3514 26774
rect 187 26694 3514 26718
rect 187 26638 3109 26694
rect 3165 26638 3190 26694
rect 3246 26638 3271 26694
rect 3327 26638 3352 26694
rect 3408 26638 3433 26694
rect 3489 26638 3514 26694
rect 187 26614 3514 26638
rect 187 26558 3109 26614
rect 3165 26558 3190 26614
rect 3246 26558 3271 26614
rect 3327 26558 3352 26614
rect 3408 26558 3433 26614
rect 3489 26558 3514 26614
rect 187 26534 3514 26558
rect 187 26478 3109 26534
rect 3165 26478 3190 26534
rect 3246 26478 3271 26534
rect 3327 26478 3352 26534
rect 3408 26478 3433 26534
rect 3489 26478 3514 26534
rect 187 26454 3514 26478
rect 187 26398 3109 26454
rect 3165 26398 3190 26454
rect 3246 26398 3271 26454
rect 3327 26398 3352 26454
rect 3408 26398 3433 26454
rect 3489 26398 3514 26454
rect 187 26374 3514 26398
rect 187 26318 3109 26374
rect 3165 26318 3190 26374
rect 3246 26318 3271 26374
rect 3327 26318 3352 26374
rect 3408 26318 3433 26374
rect 3489 26318 3514 26374
rect 187 26294 3514 26318
rect 187 26238 3109 26294
rect 3165 26238 3190 26294
rect 3246 26238 3271 26294
rect 3327 26238 3352 26294
rect 3408 26238 3433 26294
rect 3489 26238 3514 26294
rect 187 26214 3514 26238
rect 187 26158 3109 26214
rect 3165 26158 3190 26214
rect 3246 26158 3271 26214
rect 3327 26158 3352 26214
rect 3408 26158 3433 26214
rect 3489 26158 3514 26214
rect 187 26134 3514 26158
rect 187 26078 3109 26134
rect 3165 26078 3190 26134
rect 3246 26078 3271 26134
rect 3327 26078 3352 26134
rect 3408 26078 3433 26134
rect 3489 26078 3514 26134
rect 187 26054 3514 26078
rect 187 25998 3109 26054
rect 3165 25998 3190 26054
rect 3246 25998 3271 26054
rect 3327 25998 3352 26054
rect 3408 25998 3433 26054
rect 3489 25998 3514 26054
rect 187 25974 3514 25998
rect 187 25918 3109 25974
rect 3165 25918 3190 25974
rect 3246 25918 3271 25974
rect 3327 25918 3352 25974
rect 3408 25918 3433 25974
rect 3489 25918 3514 25974
rect 187 25894 3514 25918
rect 187 25838 3109 25894
rect 3165 25838 3190 25894
rect 3246 25838 3271 25894
rect 3327 25838 3352 25894
rect 3408 25838 3433 25894
rect 3489 25838 3514 25894
rect 187 25814 3514 25838
rect 187 25758 3109 25814
rect 3165 25758 3190 25814
rect 3246 25758 3271 25814
rect 3327 25758 3352 25814
rect 3408 25758 3433 25814
rect 3489 25758 3514 25814
rect 187 25734 3514 25758
rect 187 25678 3109 25734
rect 3165 25678 3190 25734
rect 3246 25678 3271 25734
rect 3327 25678 3352 25734
rect 3408 25678 3433 25734
rect 3489 25678 3514 25734
rect 187 25654 3514 25678
rect 187 25598 3109 25654
rect 3165 25598 3190 25654
rect 3246 25598 3271 25654
rect 3327 25598 3352 25654
rect 3408 25598 3433 25654
rect 3489 25598 3514 25654
rect 187 25574 3514 25598
rect 187 25518 3109 25574
rect 3165 25518 3190 25574
rect 3246 25518 3271 25574
rect 3327 25518 3352 25574
rect 3408 25518 3433 25574
rect 3489 25518 3514 25574
rect 187 25494 3514 25518
rect 187 25438 3109 25494
rect 3165 25438 3190 25494
rect 3246 25438 3271 25494
rect 3327 25438 3352 25494
rect 3408 25438 3433 25494
rect 3489 25438 3514 25494
rect 187 25414 3514 25438
rect 187 25358 3109 25414
rect 3165 25358 3190 25414
rect 3246 25358 3271 25414
rect 3327 25358 3352 25414
rect 3408 25358 3433 25414
rect 3489 25358 3514 25414
rect 4290 27090 5195 27094
rect 4290 27038 4780 27090
rect 4832 27038 4848 27090
rect 4900 27038 5195 27090
rect 5251 27038 5276 27094
rect 5332 27038 5357 27094
rect 5413 27038 5438 27094
rect 5494 27038 5519 27094
rect 5575 27038 5600 27094
rect 6376 27090 11341 27094
rect 6376 27038 6552 27090
rect 6604 27038 6620 27090
rect 6672 27038 6688 27090
rect 6740 27038 7472 27090
rect 7524 27038 7540 27090
rect 7592 27038 7608 27090
rect 7660 27038 8392 27090
rect 8444 27038 8460 27090
rect 8512 27038 8528 27090
rect 8580 27038 9312 27090
rect 9364 27038 9380 27090
rect 9432 27038 9448 27090
rect 9500 27038 10232 27090
rect 10284 27038 10300 27090
rect 10352 27038 10368 27090
rect 10420 27038 11152 27090
rect 11204 27038 11220 27090
rect 11272 27038 11288 27090
rect 11340 27038 11341 27090
rect 4290 27026 5600 27038
rect 6376 27026 11341 27038
rect 4290 26974 4780 27026
rect 4832 26974 4848 27026
rect 4900 27014 5600 27026
rect 4900 26974 5195 27014
rect 4290 26962 5195 26974
rect 4290 26910 4780 26962
rect 4832 26910 4848 26962
rect 4900 26958 5195 26962
rect 5251 26958 5276 27014
rect 5332 26958 5357 27014
rect 5413 26958 5438 27014
rect 5494 26958 5519 27014
rect 5575 26958 5600 27014
rect 6376 26974 6552 27026
rect 6604 26974 6620 27026
rect 6672 26974 6688 27026
rect 6740 26974 7472 27026
rect 7524 26974 7540 27026
rect 7592 26974 7608 27026
rect 7660 26974 8392 27026
rect 8444 26974 8460 27026
rect 8512 26974 8528 27026
rect 8580 26974 9312 27026
rect 9364 26974 9380 27026
rect 9432 26974 9448 27026
rect 9500 26974 10232 27026
rect 10284 26974 10300 27026
rect 10352 26974 10368 27026
rect 10420 26974 11152 27026
rect 11204 26974 11220 27026
rect 11272 26974 11288 27026
rect 11340 26974 11341 27026
rect 6376 26962 11341 26974
rect 4900 26934 5600 26958
rect 4900 26910 5195 26934
rect 4290 26898 5195 26910
rect 4290 26846 4780 26898
rect 4832 26846 4848 26898
rect 4900 26878 5195 26898
rect 5251 26878 5276 26934
rect 5332 26878 5357 26934
rect 5413 26878 5438 26934
rect 5494 26878 5519 26934
rect 5575 26878 5600 26934
rect 6376 26910 6552 26962
rect 6604 26910 6620 26962
rect 6672 26910 6688 26962
rect 6740 26910 7472 26962
rect 7524 26910 7540 26962
rect 7592 26910 7608 26962
rect 7660 26910 8392 26962
rect 8444 26910 8460 26962
rect 8512 26910 8528 26962
rect 8580 26910 9312 26962
rect 9364 26910 9380 26962
rect 9432 26910 9448 26962
rect 9500 26910 10232 26962
rect 10284 26910 10300 26962
rect 10352 26910 10368 26962
rect 10420 26910 11152 26962
rect 11204 26910 11220 26962
rect 11272 26910 11288 26962
rect 11340 26910 11341 26962
rect 6376 26898 11341 26910
rect 4900 26854 5600 26878
rect 4900 26846 5195 26854
rect 4290 26834 5195 26846
rect 4290 26782 4780 26834
rect 4832 26782 4848 26834
rect 4900 26798 5195 26834
rect 5251 26798 5276 26854
rect 5332 26798 5357 26854
rect 5413 26798 5438 26854
rect 5494 26798 5519 26854
rect 5575 26798 5600 26854
rect 6376 26846 6552 26898
rect 6604 26846 6620 26898
rect 6672 26846 6688 26898
rect 6740 26846 7472 26898
rect 7524 26846 7540 26898
rect 7592 26846 7608 26898
rect 7660 26846 8392 26898
rect 8444 26846 8460 26898
rect 8512 26846 8528 26898
rect 8580 26846 9312 26898
rect 9364 26846 9380 26898
rect 9432 26846 9448 26898
rect 9500 26846 10232 26898
rect 10284 26846 10300 26898
rect 10352 26846 10368 26898
rect 10420 26846 11152 26898
rect 11204 26846 11220 26898
rect 11272 26846 11288 26898
rect 11340 26846 11341 26898
rect 6376 26834 11341 26846
rect 4900 26782 5600 26798
rect 6376 26782 6552 26834
rect 6604 26782 6620 26834
rect 6672 26782 6688 26834
rect 6740 26782 7472 26834
rect 7524 26782 7540 26834
rect 7592 26782 7608 26834
rect 7660 26782 8392 26834
rect 8444 26782 8460 26834
rect 8512 26782 8528 26834
rect 8580 26782 9312 26834
rect 9364 26782 9380 26834
rect 9432 26782 9448 26834
rect 9500 26782 10232 26834
rect 10284 26782 10300 26834
rect 10352 26782 10368 26834
rect 10420 26782 11152 26834
rect 11204 26782 11220 26834
rect 11272 26782 11288 26834
rect 11340 26782 11341 26834
rect 4290 26774 5600 26782
rect 4290 26770 5195 26774
rect 4290 26718 4780 26770
rect 4832 26718 4848 26770
rect 4900 26718 5195 26770
rect 5251 26718 5276 26774
rect 5332 26718 5357 26774
rect 5413 26718 5438 26774
rect 5494 26718 5519 26774
rect 5575 26718 5600 26774
rect 6376 26770 11341 26782
rect 6376 26718 6552 26770
rect 6604 26718 6620 26770
rect 6672 26718 6688 26770
rect 6740 26718 7472 26770
rect 7524 26718 7540 26770
rect 7592 26718 7608 26770
rect 7660 26718 8392 26770
rect 8444 26718 8460 26770
rect 8512 26718 8528 26770
rect 8580 26718 9312 26770
rect 9364 26718 9380 26770
rect 9432 26718 9448 26770
rect 9500 26718 10232 26770
rect 10284 26718 10300 26770
rect 10352 26718 10368 26770
rect 10420 26718 11152 26770
rect 11204 26718 11220 26770
rect 11272 26718 11288 26770
rect 11340 26718 11341 26770
rect 4290 26706 5600 26718
rect 6376 26706 11341 26718
rect 4290 26654 4780 26706
rect 4832 26654 4848 26706
rect 4900 26694 5600 26706
rect 4900 26654 5195 26694
rect 4290 26642 5195 26654
rect 4290 26590 4780 26642
rect 4832 26590 4848 26642
rect 4900 26638 5195 26642
rect 5251 26638 5276 26694
rect 5332 26638 5357 26694
rect 5413 26638 5438 26694
rect 5494 26638 5519 26694
rect 5575 26638 5600 26694
rect 6376 26654 6552 26706
rect 6604 26654 6620 26706
rect 6672 26654 6688 26706
rect 6740 26654 7472 26706
rect 7524 26654 7540 26706
rect 7592 26654 7608 26706
rect 7660 26654 8392 26706
rect 8444 26654 8460 26706
rect 8512 26654 8528 26706
rect 8580 26654 9312 26706
rect 9364 26654 9380 26706
rect 9432 26654 9448 26706
rect 9500 26654 10232 26706
rect 10284 26654 10300 26706
rect 10352 26654 10368 26706
rect 10420 26654 11152 26706
rect 11204 26654 11220 26706
rect 11272 26654 11288 26706
rect 11340 26654 11341 26706
rect 6376 26642 11341 26654
rect 4900 26614 5600 26638
rect 4900 26590 5195 26614
rect 4290 26578 5195 26590
rect 4290 26526 4780 26578
rect 4832 26526 4848 26578
rect 4900 26558 5195 26578
rect 5251 26558 5276 26614
rect 5332 26558 5357 26614
rect 5413 26558 5438 26614
rect 5494 26558 5519 26614
rect 5575 26558 5600 26614
rect 6376 26590 6552 26642
rect 6604 26590 6620 26642
rect 6672 26590 6688 26642
rect 6740 26590 7472 26642
rect 7524 26590 7540 26642
rect 7592 26590 7608 26642
rect 7660 26590 8392 26642
rect 8444 26590 8460 26642
rect 8512 26590 8528 26642
rect 8580 26590 9312 26642
rect 9364 26590 9380 26642
rect 9432 26590 9448 26642
rect 9500 26590 10232 26642
rect 10284 26590 10300 26642
rect 10352 26590 10368 26642
rect 10420 26590 11152 26642
rect 11204 26590 11220 26642
rect 11272 26590 11288 26642
rect 11340 26590 11341 26642
rect 6376 26578 11341 26590
rect 4900 26534 5600 26558
rect 4900 26526 5195 26534
rect 4290 26514 5195 26526
rect 4290 26462 4780 26514
rect 4832 26462 4848 26514
rect 4900 26478 5195 26514
rect 5251 26478 5276 26534
rect 5332 26478 5357 26534
rect 5413 26478 5438 26534
rect 5494 26478 5519 26534
rect 5575 26478 5600 26534
rect 6376 26526 6552 26578
rect 6604 26526 6620 26578
rect 6672 26526 6688 26578
rect 6740 26526 7472 26578
rect 7524 26526 7540 26578
rect 7592 26526 7608 26578
rect 7660 26526 8392 26578
rect 8444 26526 8460 26578
rect 8512 26526 8528 26578
rect 8580 26526 9312 26578
rect 9364 26526 9380 26578
rect 9432 26526 9448 26578
rect 9500 26526 10232 26578
rect 10284 26526 10300 26578
rect 10352 26526 10368 26578
rect 10420 26526 11152 26578
rect 11204 26526 11220 26578
rect 11272 26526 11288 26578
rect 11340 26526 11341 26578
rect 6376 26514 11341 26526
rect 4900 26462 5600 26478
rect 6376 26462 6552 26514
rect 6604 26462 6620 26514
rect 6672 26462 6688 26514
rect 6740 26462 7472 26514
rect 7524 26462 7540 26514
rect 7592 26462 7608 26514
rect 7660 26462 8392 26514
rect 8444 26462 8460 26514
rect 8512 26462 8528 26514
rect 8580 26462 9312 26514
rect 9364 26462 9380 26514
rect 9432 26462 9448 26514
rect 9500 26462 10232 26514
rect 10284 26462 10300 26514
rect 10352 26462 10368 26514
rect 10420 26462 11152 26514
rect 11204 26462 11220 26514
rect 11272 26462 11288 26514
rect 11340 26462 11341 26514
rect 4290 26454 5600 26462
rect 4290 26450 5195 26454
rect 4290 26398 4780 26450
rect 4832 26398 4848 26450
rect 4900 26398 5195 26450
rect 5251 26398 5276 26454
rect 5332 26398 5357 26454
rect 5413 26398 5438 26454
rect 5494 26398 5519 26454
rect 5575 26398 5600 26454
rect 6376 26450 11341 26462
rect 6376 26398 6552 26450
rect 6604 26398 6620 26450
rect 6672 26398 6688 26450
rect 6740 26398 7472 26450
rect 7524 26398 7540 26450
rect 7592 26398 7608 26450
rect 7660 26398 8392 26450
rect 8444 26398 8460 26450
rect 8512 26398 8528 26450
rect 8580 26398 9312 26450
rect 9364 26398 9380 26450
rect 9432 26398 9448 26450
rect 9500 26398 10232 26450
rect 10284 26398 10300 26450
rect 10352 26398 10368 26450
rect 10420 26398 11152 26450
rect 11204 26398 11220 26450
rect 11272 26398 11288 26450
rect 11340 26398 11341 26450
rect 4290 26386 5600 26398
rect 6376 26386 11341 26398
rect 4290 26334 4780 26386
rect 4832 26334 4848 26386
rect 4900 26374 5600 26386
rect 4900 26334 5195 26374
rect 4290 26322 5195 26334
rect 4290 26270 4780 26322
rect 4832 26270 4848 26322
rect 4900 26318 5195 26322
rect 5251 26318 5276 26374
rect 5332 26318 5357 26374
rect 5413 26318 5438 26374
rect 5494 26318 5519 26374
rect 5575 26318 5600 26374
rect 6376 26334 6552 26386
rect 6604 26334 6620 26386
rect 6672 26334 6688 26386
rect 6740 26334 7472 26386
rect 7524 26334 7540 26386
rect 7592 26334 7608 26386
rect 7660 26334 8392 26386
rect 8444 26334 8460 26386
rect 8512 26334 8528 26386
rect 8580 26334 9312 26386
rect 9364 26334 9380 26386
rect 9432 26334 9448 26386
rect 9500 26334 10232 26386
rect 10284 26334 10300 26386
rect 10352 26334 10368 26386
rect 10420 26334 11152 26386
rect 11204 26334 11220 26386
rect 11272 26334 11288 26386
rect 11340 26334 11341 26386
rect 6376 26322 11341 26334
rect 4900 26294 5600 26318
rect 4900 26270 5195 26294
rect 4290 26258 5195 26270
rect 4290 26206 4780 26258
rect 4832 26206 4848 26258
rect 4900 26238 5195 26258
rect 5251 26238 5276 26294
rect 5332 26238 5357 26294
rect 5413 26238 5438 26294
rect 5494 26238 5519 26294
rect 5575 26238 5600 26294
rect 6376 26270 6552 26322
rect 6604 26270 6620 26322
rect 6672 26270 6688 26322
rect 6740 26270 7472 26322
rect 7524 26270 7540 26322
rect 7592 26270 7608 26322
rect 7660 26270 8392 26322
rect 8444 26270 8460 26322
rect 8512 26270 8528 26322
rect 8580 26270 9312 26322
rect 9364 26270 9380 26322
rect 9432 26270 9448 26322
rect 9500 26270 10232 26322
rect 10284 26270 10300 26322
rect 10352 26270 10368 26322
rect 10420 26270 11152 26322
rect 11204 26270 11220 26322
rect 11272 26270 11288 26322
rect 11340 26270 11341 26322
rect 6376 26258 11341 26270
rect 4900 26214 5600 26238
rect 4900 26206 5195 26214
rect 4290 26194 5195 26206
rect 4290 26142 4780 26194
rect 4832 26142 4848 26194
rect 4900 26158 5195 26194
rect 5251 26158 5276 26214
rect 5332 26158 5357 26214
rect 5413 26158 5438 26214
rect 5494 26158 5519 26214
rect 5575 26158 5600 26214
rect 6376 26206 6552 26258
rect 6604 26206 6620 26258
rect 6672 26206 6688 26258
rect 6740 26206 7472 26258
rect 7524 26206 7540 26258
rect 7592 26206 7608 26258
rect 7660 26206 8392 26258
rect 8444 26206 8460 26258
rect 8512 26206 8528 26258
rect 8580 26206 9312 26258
rect 9364 26206 9380 26258
rect 9432 26206 9448 26258
rect 9500 26206 10232 26258
rect 10284 26206 10300 26258
rect 10352 26206 10368 26258
rect 10420 26206 11152 26258
rect 11204 26206 11220 26258
rect 11272 26206 11288 26258
rect 11340 26206 11341 26258
rect 6376 26194 11341 26206
rect 4900 26142 5600 26158
rect 6376 26142 6552 26194
rect 6604 26142 6620 26194
rect 6672 26142 6688 26194
rect 6740 26142 7472 26194
rect 7524 26142 7540 26194
rect 7592 26142 7608 26194
rect 7660 26142 8392 26194
rect 8444 26142 8460 26194
rect 8512 26142 8528 26194
rect 8580 26142 9312 26194
rect 9364 26142 9380 26194
rect 9432 26142 9448 26194
rect 9500 26142 10232 26194
rect 10284 26142 10300 26194
rect 10352 26142 10368 26194
rect 10420 26142 11152 26194
rect 11204 26142 11220 26194
rect 11272 26142 11288 26194
rect 11340 26142 11341 26194
rect 4290 26134 5600 26142
rect 4290 26129 5195 26134
rect 4290 26077 4780 26129
rect 4832 26077 4848 26129
rect 4900 26078 5195 26129
rect 5251 26078 5276 26134
rect 5332 26078 5357 26134
rect 5413 26078 5438 26134
rect 5494 26078 5519 26134
rect 5575 26078 5600 26134
rect 6376 26129 11341 26142
rect 4900 26077 5600 26078
rect 6376 26077 6552 26129
rect 6604 26077 6620 26129
rect 6672 26077 6688 26129
rect 6740 26077 7472 26129
rect 7524 26077 7540 26129
rect 7592 26077 7608 26129
rect 7660 26077 8392 26129
rect 8444 26077 8460 26129
rect 8512 26077 8528 26129
rect 8580 26077 9312 26129
rect 9364 26077 9380 26129
rect 9432 26077 9448 26129
rect 9500 26077 10232 26129
rect 10284 26077 10300 26129
rect 10352 26077 10368 26129
rect 10420 26077 11152 26129
rect 11204 26077 11220 26129
rect 11272 26077 11288 26129
rect 11340 26077 11341 26129
rect 4290 26064 5600 26077
rect 6376 26064 11341 26077
rect 4290 26012 4780 26064
rect 4832 26012 4848 26064
rect 4900 26054 5600 26064
rect 4900 26012 5195 26054
rect 4290 25999 5195 26012
rect 4290 25947 4780 25999
rect 4832 25947 4848 25999
rect 4900 25998 5195 25999
rect 5251 25998 5276 26054
rect 5332 25998 5357 26054
rect 5413 25998 5438 26054
rect 5494 25998 5519 26054
rect 5575 25998 5600 26054
rect 6376 26012 6552 26064
rect 6604 26012 6620 26064
rect 6672 26012 6688 26064
rect 6740 26012 7472 26064
rect 7524 26012 7540 26064
rect 7592 26012 7608 26064
rect 7660 26012 8392 26064
rect 8444 26012 8460 26064
rect 8512 26012 8528 26064
rect 8580 26012 9312 26064
rect 9364 26012 9380 26064
rect 9432 26012 9448 26064
rect 9500 26012 10232 26064
rect 10284 26012 10300 26064
rect 10352 26012 10368 26064
rect 10420 26012 11152 26064
rect 11204 26012 11220 26064
rect 11272 26012 11288 26064
rect 11340 26012 11341 26064
rect 6376 25999 11341 26012
rect 4900 25974 5600 25998
rect 4900 25947 5195 25974
rect 4290 25934 5195 25947
rect 4290 25882 4780 25934
rect 4832 25882 4848 25934
rect 4900 25918 5195 25934
rect 5251 25918 5276 25974
rect 5332 25918 5357 25974
rect 5413 25918 5438 25974
rect 5494 25918 5519 25974
rect 5575 25918 5600 25974
rect 6376 25947 6552 25999
rect 6604 25947 6620 25999
rect 6672 25947 6688 25999
rect 6740 25947 7472 25999
rect 7524 25947 7540 25999
rect 7592 25947 7608 25999
rect 7660 25947 8392 25999
rect 8444 25947 8460 25999
rect 8512 25947 8528 25999
rect 8580 25947 9312 25999
rect 9364 25947 9380 25999
rect 9432 25947 9448 25999
rect 9500 25947 10232 25999
rect 10284 25947 10300 25999
rect 10352 25947 10368 25999
rect 10420 25947 11152 25999
rect 11204 25947 11220 25999
rect 11272 25947 11288 25999
rect 11340 25947 11341 25999
rect 6376 25934 11341 25947
rect 4900 25894 5600 25918
rect 4900 25882 5195 25894
rect 4290 25869 5195 25882
rect 4290 25817 4780 25869
rect 4832 25817 4848 25869
rect 4900 25838 5195 25869
rect 5251 25838 5276 25894
rect 5332 25838 5357 25894
rect 5413 25838 5438 25894
rect 5494 25838 5519 25894
rect 5575 25838 5600 25894
rect 6376 25882 6552 25934
rect 6604 25882 6620 25934
rect 6672 25882 6688 25934
rect 6740 25882 7472 25934
rect 7524 25882 7540 25934
rect 7592 25882 7608 25934
rect 7660 25882 8392 25934
rect 8444 25882 8460 25934
rect 8512 25882 8528 25934
rect 8580 25882 9312 25934
rect 9364 25882 9380 25934
rect 9432 25882 9448 25934
rect 9500 25882 10232 25934
rect 10284 25882 10300 25934
rect 10352 25882 10368 25934
rect 10420 25882 11152 25934
rect 11204 25882 11220 25934
rect 11272 25882 11288 25934
rect 11340 25882 11341 25934
rect 6376 25869 11341 25882
rect 4900 25817 5600 25838
rect 6376 25817 6552 25869
rect 6604 25817 6620 25869
rect 6672 25817 6688 25869
rect 6740 25817 7472 25869
rect 7524 25817 7540 25869
rect 7592 25817 7608 25869
rect 7660 25817 8392 25869
rect 8444 25817 8460 25869
rect 8512 25817 8528 25869
rect 8580 25817 9312 25869
rect 9364 25817 9380 25869
rect 9432 25817 9448 25869
rect 9500 25817 10232 25869
rect 10284 25817 10300 25869
rect 10352 25817 10368 25869
rect 10420 25817 11152 25869
rect 11204 25817 11220 25869
rect 11272 25817 11288 25869
rect 11340 25817 11341 25869
rect 4290 25814 5600 25817
rect 4290 25804 5195 25814
rect 4290 25752 4780 25804
rect 4832 25752 4848 25804
rect 4900 25758 5195 25804
rect 5251 25758 5276 25814
rect 5332 25758 5357 25814
rect 5413 25758 5438 25814
rect 5494 25758 5519 25814
rect 5575 25758 5600 25814
rect 6376 25804 11341 25817
rect 4900 25752 5600 25758
rect 6376 25752 6552 25804
rect 6604 25752 6620 25804
rect 6672 25752 6688 25804
rect 6740 25752 7472 25804
rect 7524 25752 7540 25804
rect 7592 25752 7608 25804
rect 7660 25752 8392 25804
rect 8444 25752 8460 25804
rect 8512 25752 8528 25804
rect 8580 25752 9312 25804
rect 9364 25752 9380 25804
rect 9432 25752 9448 25804
rect 9500 25752 10232 25804
rect 10284 25752 10300 25804
rect 10352 25752 10368 25804
rect 10420 25752 11152 25804
rect 11204 25752 11220 25804
rect 11272 25752 11288 25804
rect 11340 25752 11341 25804
rect 4290 25739 5600 25752
rect 6376 25739 11341 25752
rect 4290 25687 4780 25739
rect 4832 25687 4848 25739
rect 4900 25734 5600 25739
rect 4900 25687 5195 25734
rect 4290 25678 5195 25687
rect 5251 25678 5276 25734
rect 5332 25678 5357 25734
rect 5413 25678 5438 25734
rect 5494 25678 5519 25734
rect 5575 25678 5600 25734
rect 6376 25687 6552 25739
rect 6604 25687 6620 25739
rect 6672 25687 6688 25739
rect 6740 25687 7472 25739
rect 7524 25687 7540 25739
rect 7592 25687 7608 25739
rect 7660 25687 8392 25739
rect 8444 25687 8460 25739
rect 8512 25687 8528 25739
rect 8580 25687 9312 25739
rect 9364 25687 9380 25739
rect 9432 25687 9448 25739
rect 9500 25687 10232 25739
rect 10284 25687 10300 25739
rect 10352 25687 10368 25739
rect 10420 25687 11152 25739
rect 11204 25687 11220 25739
rect 11272 25687 11288 25739
rect 11340 25687 11341 25739
rect 4290 25674 5600 25678
rect 6376 25674 11341 25687
rect 4290 25622 4780 25674
rect 4832 25622 4848 25674
rect 4900 25654 5600 25674
rect 4900 25622 5195 25654
rect 4290 25609 5195 25622
rect 4290 25557 4780 25609
rect 4832 25557 4848 25609
rect 4900 25598 5195 25609
rect 5251 25598 5276 25654
rect 5332 25598 5357 25654
rect 5413 25598 5438 25654
rect 5494 25598 5519 25654
rect 5575 25598 5600 25654
rect 6376 25622 6552 25674
rect 6604 25622 6620 25674
rect 6672 25622 6688 25674
rect 6740 25622 7472 25674
rect 7524 25622 7540 25674
rect 7592 25622 7608 25674
rect 7660 25622 8392 25674
rect 8444 25622 8460 25674
rect 8512 25622 8528 25674
rect 8580 25622 9312 25674
rect 9364 25622 9380 25674
rect 9432 25622 9448 25674
rect 9500 25622 10232 25674
rect 10284 25622 10300 25674
rect 10352 25622 10368 25674
rect 10420 25622 11152 25674
rect 11204 25622 11220 25674
rect 11272 25622 11288 25674
rect 11340 25622 11341 25674
rect 6376 25609 11341 25622
rect 4900 25574 5600 25598
rect 4900 25557 5195 25574
rect 4290 25544 5195 25557
rect 4290 25492 4780 25544
rect 4832 25492 4848 25544
rect 4900 25518 5195 25544
rect 5251 25518 5276 25574
rect 5332 25518 5357 25574
rect 5413 25518 5438 25574
rect 5494 25518 5519 25574
rect 5575 25518 5600 25574
rect 6376 25557 6552 25609
rect 6604 25557 6620 25609
rect 6672 25557 6688 25609
rect 6740 25557 7472 25609
rect 7524 25557 7540 25609
rect 7592 25557 7608 25609
rect 7660 25557 8392 25609
rect 8444 25557 8460 25609
rect 8512 25557 8528 25609
rect 8580 25557 9312 25609
rect 9364 25557 9380 25609
rect 9432 25557 9448 25609
rect 9500 25557 10232 25609
rect 10284 25557 10300 25609
rect 10352 25557 10368 25609
rect 10420 25557 11152 25609
rect 11204 25557 11220 25609
rect 11272 25557 11288 25609
rect 11340 25557 11341 25609
rect 6376 25544 11341 25557
rect 4900 25494 5600 25518
rect 4900 25492 5195 25494
rect 4290 25479 5195 25492
rect 4290 25427 4780 25479
rect 4832 25427 4848 25479
rect 4900 25438 5195 25479
rect 5251 25438 5276 25494
rect 5332 25438 5357 25494
rect 5413 25438 5438 25494
rect 5494 25438 5519 25494
rect 5575 25438 5600 25494
rect 6376 25492 6552 25544
rect 6604 25492 6620 25544
rect 6672 25492 6688 25544
rect 6740 25492 7472 25544
rect 7524 25492 7540 25544
rect 7592 25492 7608 25544
rect 7660 25492 8392 25544
rect 8444 25492 8460 25544
rect 8512 25492 8528 25544
rect 8580 25492 9312 25544
rect 9364 25492 9380 25544
rect 9432 25492 9448 25544
rect 9500 25492 10232 25544
rect 10284 25492 10300 25544
rect 10352 25492 10368 25544
rect 10420 25492 11152 25544
rect 11204 25492 11220 25544
rect 11272 25492 11288 25544
rect 11340 25492 11341 25544
rect 6376 25479 11341 25492
rect 4900 25427 5600 25438
rect 6376 25427 6552 25479
rect 6604 25427 6620 25479
rect 6672 25427 6688 25479
rect 6740 25427 7472 25479
rect 7524 25427 7540 25479
rect 7592 25427 7608 25479
rect 7660 25427 8392 25479
rect 8444 25427 8460 25479
rect 8512 25427 8528 25479
rect 8580 25427 9312 25479
rect 9364 25427 9380 25479
rect 9432 25427 9448 25479
rect 9500 25427 10232 25479
rect 10284 25427 10300 25479
rect 10352 25427 10368 25479
rect 10420 25427 11152 25479
rect 11204 25427 11220 25479
rect 11272 25427 11288 25479
rect 11340 25427 11341 25479
rect 4290 25414 5600 25427
rect 6376 25414 11341 25427
rect 4290 25362 4780 25414
rect 4832 25362 4848 25414
rect 4900 25362 5195 25414
rect 4290 25358 5195 25362
rect 5251 25358 5276 25414
rect 5332 25358 5357 25414
rect 5413 25358 5438 25414
rect 5494 25358 5519 25414
rect 5575 25358 5600 25414
rect 6376 25362 6552 25414
rect 6604 25362 6620 25414
rect 6672 25362 6688 25414
rect 6740 25362 7472 25414
rect 7524 25362 7540 25414
rect 7592 25362 7608 25414
rect 7660 25362 8392 25414
rect 8444 25362 8460 25414
rect 8512 25362 8528 25414
rect 8580 25362 9312 25414
rect 9364 25362 9380 25414
rect 9432 25362 9448 25414
rect 9500 25362 10232 25414
rect 10284 25362 10300 25414
rect 10352 25362 10368 25414
rect 10420 25362 11152 25414
rect 11204 25362 11220 25414
rect 11272 25362 11288 25414
rect 11340 25362 11341 25414
rect 6376 25358 11341 25362
rect 187 25356 11341 25358
rect 187 22496 2824 25356
tri 2824 24629 3551 25356 nw
tri 11511 25031 12222 25742 se
rect 12222 25031 14858 27891
rect 4964 25029 14858 25031
rect 4964 25025 8580 25029
rect 4964 24973 5201 25025
rect 5253 24973 5279 25025
rect 5331 24973 6121 25025
rect 6173 24973 6199 25025
rect 6251 24973 7041 25025
rect 7093 24973 7119 25025
rect 7171 24973 7961 25025
rect 8013 24973 8039 25025
rect 8091 24973 8580 25025
rect 8636 24973 8661 25029
rect 8717 24973 8742 25029
rect 8798 24973 8823 25029
rect 8879 25025 8904 25029
rect 8960 25025 8985 25029
rect 8879 24973 8881 25025
rect 9041 24973 9066 25029
rect 4964 24961 9066 24973
rect 4964 24909 5201 24961
rect 5253 24909 5279 24961
rect 5331 24909 6121 24961
rect 6173 24909 6199 24961
rect 6251 24909 7041 24961
rect 7093 24909 7119 24961
rect 7171 24909 7961 24961
rect 8013 24909 8039 24961
rect 8091 24949 8881 24961
rect 8933 24949 8959 24961
rect 9011 24949 9066 24961
rect 8091 24909 8580 24949
rect 4964 24897 8580 24909
rect 4964 24845 5201 24897
rect 5253 24845 5279 24897
rect 5331 24845 6121 24897
rect 6173 24845 6199 24897
rect 6251 24845 7041 24897
rect 7093 24845 7119 24897
rect 7171 24845 7961 24897
rect 8013 24845 8039 24897
rect 8091 24893 8580 24897
rect 8636 24893 8661 24949
rect 8717 24893 8742 24949
rect 8798 24893 8823 24949
rect 8879 24909 8881 24949
rect 8879 24897 8904 24909
rect 8960 24897 8985 24909
rect 8879 24893 8881 24897
rect 9041 24893 9066 24949
rect 8091 24869 8881 24893
rect 8933 24869 8959 24893
rect 9011 24869 9066 24893
rect 8091 24845 8580 24869
rect 4964 24833 8580 24845
rect 4964 24781 5201 24833
rect 5253 24781 5279 24833
rect 5331 24781 6121 24833
rect 6173 24781 6199 24833
rect 6251 24781 7041 24833
rect 7093 24781 7119 24833
rect 7171 24781 7961 24833
rect 8013 24781 8039 24833
rect 8091 24813 8580 24833
rect 8636 24813 8661 24869
rect 8717 24813 8742 24869
rect 8798 24813 8823 24869
rect 8879 24845 8881 24869
rect 8879 24833 8904 24845
rect 8960 24833 8985 24845
rect 8879 24813 8881 24833
rect 9041 24813 9066 24869
rect 8091 24789 8881 24813
rect 8933 24789 8959 24813
rect 9011 24789 9066 24813
rect 8091 24781 8580 24789
rect 4964 24769 8580 24781
rect 4964 24717 5201 24769
rect 5253 24717 5279 24769
rect 5331 24717 6121 24769
rect 6173 24717 6199 24769
rect 6251 24717 7041 24769
rect 7093 24717 7119 24769
rect 7171 24717 7961 24769
rect 8013 24717 8039 24769
rect 8091 24733 8580 24769
rect 8636 24733 8661 24789
rect 8717 24733 8742 24789
rect 8798 24733 8823 24789
rect 8879 24781 8881 24789
rect 8879 24769 8904 24781
rect 8960 24769 8985 24781
rect 8879 24733 8881 24769
rect 9041 24733 9066 24789
rect 8091 24717 8881 24733
rect 8933 24717 8959 24733
rect 9011 24717 9066 24733
rect 4964 24709 9066 24717
rect 4964 24705 8580 24709
rect 4964 24653 5201 24705
rect 5253 24653 5279 24705
rect 5331 24653 6121 24705
rect 6173 24653 6199 24705
rect 6251 24653 7041 24705
rect 7093 24653 7119 24705
rect 7171 24653 7961 24705
rect 8013 24653 8039 24705
rect 8091 24653 8580 24705
rect 8636 24653 8661 24709
rect 8717 24653 8742 24709
rect 8798 24653 8823 24709
rect 8879 24705 8904 24709
rect 8960 24705 8985 24709
rect 8879 24653 8881 24705
rect 9041 24653 9066 24709
rect 4964 24641 9066 24653
rect 4964 24589 5201 24641
rect 5253 24589 5279 24641
rect 5331 24589 6121 24641
rect 6173 24589 6199 24641
rect 6251 24589 7041 24641
rect 7093 24589 7119 24641
rect 7171 24589 7961 24641
rect 8013 24589 8039 24641
rect 8091 24629 8881 24641
rect 8933 24629 8959 24641
rect 9011 24629 9066 24641
rect 8091 24589 8580 24629
rect 4964 24577 8580 24589
rect 4964 24525 5201 24577
rect 5253 24525 5279 24577
rect 5331 24525 6121 24577
rect 6173 24525 6199 24577
rect 6251 24525 7041 24577
rect 7093 24525 7119 24577
rect 7171 24525 7961 24577
rect 8013 24525 8039 24577
rect 8091 24573 8580 24577
rect 8636 24573 8661 24629
rect 8717 24573 8742 24629
rect 8798 24573 8823 24629
rect 8879 24589 8881 24629
rect 8879 24577 8904 24589
rect 8960 24577 8985 24589
rect 8879 24573 8881 24577
rect 9041 24573 9066 24629
rect 8091 24549 8881 24573
rect 8933 24549 8959 24573
rect 9011 24549 9066 24573
rect 8091 24525 8580 24549
rect 4964 24513 8580 24525
rect 4964 24461 5201 24513
rect 5253 24461 5279 24513
rect 5331 24461 6121 24513
rect 6173 24461 6199 24513
rect 6251 24461 7041 24513
rect 7093 24461 7119 24513
rect 7171 24461 7961 24513
rect 8013 24461 8039 24513
rect 8091 24493 8580 24513
rect 8636 24493 8661 24549
rect 8717 24493 8742 24549
rect 8798 24493 8823 24549
rect 8879 24525 8881 24549
rect 8879 24513 8904 24525
rect 8960 24513 8985 24525
rect 8879 24493 8881 24513
rect 9041 24493 9066 24549
rect 8091 24469 8881 24493
rect 8933 24469 8959 24493
rect 9011 24469 9066 24493
rect 8091 24461 8580 24469
rect 4964 24449 8580 24461
rect 4964 24397 5201 24449
rect 5253 24397 5279 24449
rect 5331 24397 6121 24449
rect 6173 24397 6199 24449
rect 6251 24397 7041 24449
rect 7093 24397 7119 24449
rect 7171 24397 7961 24449
rect 8013 24397 8039 24449
rect 8091 24413 8580 24449
rect 8636 24413 8661 24469
rect 8717 24413 8742 24469
rect 8798 24413 8823 24469
rect 8879 24461 8881 24469
rect 8879 24449 8904 24461
rect 8960 24449 8985 24461
rect 8879 24413 8881 24449
rect 9041 24413 9066 24469
rect 8091 24397 8881 24413
rect 8933 24397 8959 24413
rect 9011 24397 9066 24413
rect 4964 24389 9066 24397
rect 4964 24385 8580 24389
rect 4964 24333 5201 24385
rect 5253 24333 5279 24385
rect 5331 24333 6121 24385
rect 6173 24333 6199 24385
rect 6251 24333 7041 24385
rect 7093 24333 7119 24385
rect 7171 24333 7961 24385
rect 8013 24333 8039 24385
rect 8091 24333 8580 24385
rect 8636 24333 8661 24389
rect 8717 24333 8742 24389
rect 8798 24333 8823 24389
rect 8879 24385 8904 24389
rect 8960 24385 8985 24389
rect 8879 24333 8881 24385
rect 9041 24333 9066 24389
rect 4964 24321 9066 24333
rect 4964 24269 5201 24321
rect 5253 24269 5279 24321
rect 5331 24269 6121 24321
rect 6173 24269 6199 24321
rect 6251 24269 7041 24321
rect 7093 24269 7119 24321
rect 7171 24269 7961 24321
rect 8013 24269 8039 24321
rect 8091 24309 8881 24321
rect 8933 24309 8959 24321
rect 9011 24309 9066 24321
rect 8091 24269 8580 24309
rect 4964 24257 8580 24269
rect 4964 24205 5201 24257
rect 5253 24205 5279 24257
rect 5331 24205 6121 24257
rect 6173 24205 6199 24257
rect 6251 24205 7041 24257
rect 7093 24205 7119 24257
rect 7171 24205 7961 24257
rect 8013 24205 8039 24257
rect 8091 24253 8580 24257
rect 8636 24253 8661 24309
rect 8717 24253 8742 24309
rect 8798 24253 8823 24309
rect 8879 24269 8881 24309
rect 8879 24257 8904 24269
rect 8960 24257 8985 24269
rect 8879 24253 8881 24257
rect 9041 24253 9066 24309
rect 8091 24229 8881 24253
rect 8933 24229 8959 24253
rect 9011 24229 9066 24253
rect 8091 24205 8580 24229
rect 4964 24193 8580 24205
rect 4964 24141 5201 24193
rect 5253 24141 5279 24193
rect 5331 24141 6121 24193
rect 6173 24141 6199 24193
rect 6251 24141 7041 24193
rect 7093 24141 7119 24193
rect 7171 24141 7961 24193
rect 8013 24141 8039 24193
rect 8091 24173 8580 24193
rect 8636 24173 8661 24229
rect 8717 24173 8742 24229
rect 8798 24173 8823 24229
rect 8879 24205 8881 24229
rect 8879 24193 8904 24205
rect 8960 24193 8985 24205
rect 8879 24173 8881 24193
rect 9041 24173 9066 24229
rect 8091 24149 8881 24173
rect 8933 24149 8959 24173
rect 9011 24149 9066 24173
rect 8091 24141 8580 24149
rect 4964 24129 8580 24141
rect 4964 24077 5201 24129
rect 5253 24077 5279 24129
rect 5331 24077 6121 24129
rect 6173 24077 6199 24129
rect 6251 24077 7041 24129
rect 7093 24077 7119 24129
rect 7171 24077 7961 24129
rect 8013 24077 8039 24129
rect 8091 24093 8580 24129
rect 8636 24093 8661 24149
rect 8717 24093 8742 24149
rect 8798 24093 8823 24149
rect 8879 24141 8881 24149
rect 8879 24129 8904 24141
rect 8960 24129 8985 24141
rect 8879 24093 8881 24129
rect 9041 24093 9066 24149
rect 8091 24077 8881 24093
rect 8933 24077 8959 24093
rect 9011 24077 9066 24093
rect 4964 24069 9066 24077
rect 4964 24064 8580 24069
rect 4964 24012 5201 24064
rect 5253 24012 5279 24064
rect 5331 24012 6121 24064
rect 6173 24012 6199 24064
rect 6251 24012 7041 24064
rect 7093 24012 7119 24064
rect 7171 24012 7961 24064
rect 8013 24012 8039 24064
rect 8091 24013 8580 24064
rect 8636 24013 8661 24069
rect 8717 24013 8742 24069
rect 8798 24013 8823 24069
rect 8879 24064 8904 24069
rect 8960 24064 8985 24069
rect 8879 24013 8881 24064
rect 9041 24013 9066 24069
rect 8091 24012 8881 24013
rect 8933 24012 8959 24013
rect 9011 24012 9066 24013
rect 4964 23999 9066 24012
rect 4964 23947 5201 23999
rect 5253 23947 5279 23999
rect 5331 23947 6121 23999
rect 6173 23947 6199 23999
rect 6251 23947 7041 23999
rect 7093 23947 7119 23999
rect 7171 23947 7961 23999
rect 8013 23947 8039 23999
rect 8091 23989 8881 23999
rect 8933 23989 8959 23999
rect 9011 23989 9066 23999
rect 8091 23947 8580 23989
rect 4964 23934 8580 23947
rect 4964 23882 5201 23934
rect 5253 23882 5279 23934
rect 5331 23882 6121 23934
rect 6173 23882 6199 23934
rect 6251 23882 7041 23934
rect 7093 23882 7119 23934
rect 7171 23882 7961 23934
rect 8013 23882 8039 23934
rect 8091 23933 8580 23934
rect 8636 23933 8661 23989
rect 8717 23933 8742 23989
rect 8798 23933 8823 23989
rect 8879 23947 8881 23989
rect 8879 23934 8904 23947
rect 8960 23934 8985 23947
rect 8879 23933 8881 23934
rect 9041 23933 9066 23989
rect 8091 23909 8881 23933
rect 8933 23909 8959 23933
rect 9011 23909 9066 23933
rect 8091 23882 8580 23909
rect 4964 23869 8580 23882
rect 4964 23817 5201 23869
rect 5253 23817 5279 23869
rect 5331 23817 6121 23869
rect 6173 23817 6199 23869
rect 6251 23817 7041 23869
rect 7093 23817 7119 23869
rect 7171 23817 7961 23869
rect 8013 23817 8039 23869
rect 8091 23853 8580 23869
rect 8636 23853 8661 23909
rect 8717 23853 8742 23909
rect 8798 23853 8823 23909
rect 8879 23882 8881 23909
rect 8879 23869 8904 23882
rect 8960 23869 8985 23882
rect 8879 23853 8881 23869
rect 9041 23853 9066 23909
rect 8091 23829 8881 23853
rect 8933 23829 8959 23853
rect 9011 23829 9066 23853
rect 8091 23817 8580 23829
rect 4964 23804 8580 23817
rect 4964 23752 5201 23804
rect 5253 23752 5279 23804
rect 5331 23752 6121 23804
rect 6173 23752 6199 23804
rect 6251 23752 7041 23804
rect 7093 23752 7119 23804
rect 7171 23752 7961 23804
rect 8013 23752 8039 23804
rect 8091 23773 8580 23804
rect 8636 23773 8661 23829
rect 8717 23773 8742 23829
rect 8798 23773 8823 23829
rect 8879 23817 8881 23829
rect 8879 23804 8904 23817
rect 8960 23804 8985 23817
rect 8879 23773 8881 23804
rect 9041 23773 9066 23829
rect 8091 23752 8881 23773
rect 8933 23752 8959 23773
rect 9011 23752 9066 23773
rect 4964 23749 9066 23752
rect 4964 23739 8580 23749
rect 4964 23687 5201 23739
rect 5253 23687 5279 23739
rect 5331 23687 6121 23739
rect 6173 23687 6199 23739
rect 6251 23687 7041 23739
rect 7093 23687 7119 23739
rect 7171 23687 7961 23739
rect 8013 23687 8039 23739
rect 8091 23693 8580 23739
rect 8636 23693 8661 23749
rect 8717 23693 8742 23749
rect 8798 23693 8823 23749
rect 8879 23739 8904 23749
rect 8960 23739 8985 23749
rect 8879 23693 8881 23739
rect 9041 23693 9066 23749
rect 8091 23687 8881 23693
rect 8933 23687 8959 23693
rect 9011 23687 9066 23693
rect 4964 23674 9066 23687
rect 4964 23622 5201 23674
rect 5253 23622 5279 23674
rect 5331 23622 6121 23674
rect 6173 23622 6199 23674
rect 6251 23622 7041 23674
rect 7093 23622 7119 23674
rect 7171 23622 7961 23674
rect 8013 23622 8039 23674
rect 8091 23669 8881 23674
rect 8933 23669 8959 23674
rect 9011 23669 9066 23674
rect 8091 23622 8580 23669
rect 4964 23613 8580 23622
rect 8636 23613 8661 23669
rect 8717 23613 8742 23669
rect 8798 23613 8823 23669
rect 8879 23622 8881 23669
rect 8879 23613 8904 23622
rect 8960 23613 8985 23622
rect 9041 23613 9066 23669
rect 4964 23609 9066 23613
rect 4964 23557 5201 23609
rect 5253 23557 5279 23609
rect 5331 23557 6121 23609
rect 6173 23557 6199 23609
rect 6251 23557 7041 23609
rect 7093 23557 7119 23609
rect 7171 23557 7961 23609
rect 8013 23557 8039 23609
rect 8091 23589 8881 23609
rect 8933 23589 8959 23609
rect 9011 23589 9066 23609
rect 8091 23557 8580 23589
rect 4964 23544 8580 23557
rect 4964 23492 5201 23544
rect 5253 23492 5279 23544
rect 5331 23492 6121 23544
rect 6173 23492 6199 23544
rect 6251 23492 7041 23544
rect 7093 23492 7119 23544
rect 7171 23492 7961 23544
rect 8013 23492 8039 23544
rect 8091 23533 8580 23544
rect 8636 23533 8661 23589
rect 8717 23533 8742 23589
rect 8798 23533 8823 23589
rect 8879 23557 8881 23589
rect 8879 23544 8904 23557
rect 8960 23544 8985 23557
rect 8879 23533 8881 23544
rect 9041 23533 9066 23589
rect 8091 23509 8881 23533
rect 8933 23509 8959 23533
rect 9011 23509 9066 23533
rect 8091 23492 8580 23509
rect 4964 23479 8580 23492
rect 3441 23432 3521 23438
rect 3441 23380 3456 23432
rect 3508 23380 3521 23432
rect 3441 23357 3521 23380
rect 3441 23305 3456 23357
rect 3508 23306 3521 23357
rect 4964 23427 5201 23479
rect 5253 23427 5279 23479
rect 5331 23427 6121 23479
rect 6173 23427 6199 23479
rect 6251 23427 7041 23479
rect 7093 23427 7119 23479
rect 7171 23427 7961 23479
rect 8013 23427 8039 23479
rect 8091 23453 8580 23479
rect 8636 23453 8661 23509
rect 8717 23453 8742 23509
rect 8798 23453 8823 23509
rect 8879 23492 8881 23509
rect 8879 23479 8904 23492
rect 8960 23479 8985 23492
rect 8879 23453 8881 23479
rect 9041 23453 9066 23509
rect 8091 23429 8881 23453
rect 8933 23429 8959 23453
rect 9011 23429 9066 23453
rect 8091 23427 8580 23429
rect 4964 23414 8580 23427
rect 4964 23362 5201 23414
rect 5253 23362 5279 23414
rect 5331 23362 6121 23414
rect 6173 23362 6199 23414
rect 6251 23362 7041 23414
rect 7093 23362 7119 23414
rect 7171 23362 7961 23414
rect 8013 23362 8039 23414
rect 8091 23373 8580 23414
rect 8636 23373 8661 23429
rect 8717 23373 8742 23429
rect 8798 23373 8823 23429
rect 8879 23427 8881 23429
rect 8879 23414 8904 23427
rect 8960 23414 8985 23427
rect 8879 23373 8881 23414
rect 9041 23373 9066 23429
rect 8091 23362 8881 23373
rect 8933 23362 8959 23373
rect 9011 23362 9066 23373
rect 4964 23349 9066 23362
tri 3521 23306 3552 23337 sw
rect 3508 23305 3718 23306
rect 3441 23297 3718 23305
tri 3718 23297 3727 23306 sw
rect 4964 23297 5201 23349
rect 5253 23297 5279 23349
rect 5331 23297 6121 23349
rect 6173 23297 6199 23349
rect 6251 23297 7041 23349
rect 7093 23297 7119 23349
rect 7171 23297 7961 23349
rect 8013 23297 8039 23349
rect 8091 23297 8580 23349
rect 3441 23291 3727 23297
tri 3727 23291 3733 23297 sw
rect 4964 23293 8580 23297
rect 8636 23293 8661 23349
rect 8717 23293 8742 23349
rect 8798 23293 8823 23349
rect 8879 23297 8881 23349
rect 8879 23293 8904 23297
rect 8960 23293 8985 23297
rect 9041 23293 9066 23349
rect 9762 25025 10666 25029
rect 10722 25025 10747 25029
rect 10803 25025 10828 25029
rect 9762 24973 9801 25025
rect 9853 24973 9879 25025
rect 9931 24973 10666 25025
rect 10884 24973 10909 25029
rect 10965 24973 10990 25029
rect 11046 24973 11071 25029
rect 11127 24973 11152 25029
rect 11848 25025 14858 25029
rect 11848 24973 12561 25025
rect 12613 24973 12639 25025
rect 12691 24973 14858 25025
rect 9762 24961 11152 24973
rect 11848 24961 14858 24973
rect 9762 24909 9801 24961
rect 9853 24909 9879 24961
rect 9931 24949 10721 24961
rect 10773 24949 10799 24961
rect 10851 24949 11152 24961
rect 9931 24909 10666 24949
rect 9762 24897 10666 24909
rect 10722 24897 10747 24909
rect 10803 24897 10828 24909
rect 9762 24845 9801 24897
rect 9853 24845 9879 24897
rect 9931 24893 10666 24897
rect 10884 24893 10909 24949
rect 10965 24893 10990 24949
rect 11046 24893 11071 24949
rect 11127 24893 11152 24949
rect 11848 24909 12561 24961
rect 12613 24909 12639 24961
rect 12691 24909 14858 24961
rect 11848 24897 14858 24909
rect 9931 24869 10721 24893
rect 10773 24869 10799 24893
rect 10851 24869 11152 24893
rect 9931 24845 10666 24869
rect 9762 24833 10666 24845
rect 10722 24833 10747 24845
rect 10803 24833 10828 24845
rect 9762 24781 9801 24833
rect 9853 24781 9879 24833
rect 9931 24813 10666 24833
rect 10884 24813 10909 24869
rect 10965 24813 10990 24869
rect 11046 24813 11071 24869
rect 11127 24813 11152 24869
rect 11848 24845 12561 24897
rect 12613 24845 12639 24897
rect 12691 24845 14858 24897
rect 11848 24833 14858 24845
rect 9931 24789 10721 24813
rect 10773 24789 10799 24813
rect 10851 24789 11152 24813
rect 9931 24781 10666 24789
rect 9762 24769 10666 24781
rect 10722 24769 10747 24781
rect 10803 24769 10828 24781
rect 9762 24717 9801 24769
rect 9853 24717 9879 24769
rect 9931 24733 10666 24769
rect 10884 24733 10909 24789
rect 10965 24733 10990 24789
rect 11046 24733 11071 24789
rect 11127 24733 11152 24789
rect 11848 24781 12561 24833
rect 12613 24781 12639 24833
rect 12691 24781 14858 24833
rect 11848 24769 14858 24781
rect 9931 24717 10721 24733
rect 10773 24717 10799 24733
rect 10851 24717 11152 24733
rect 11848 24717 12561 24769
rect 12613 24717 12639 24769
rect 12691 24717 14858 24769
rect 9762 24709 11152 24717
rect 9762 24705 10666 24709
rect 10722 24705 10747 24709
rect 10803 24705 10828 24709
rect 9762 24653 9801 24705
rect 9853 24653 9879 24705
rect 9931 24653 10666 24705
rect 10884 24653 10909 24709
rect 10965 24653 10990 24709
rect 11046 24653 11071 24709
rect 11127 24653 11152 24709
rect 11848 24705 14858 24717
rect 11848 24653 12561 24705
rect 12613 24653 12639 24705
rect 12691 24653 14858 24705
rect 9762 24641 11152 24653
rect 11848 24641 14858 24653
rect 9762 24589 9801 24641
rect 9853 24589 9879 24641
rect 9931 24629 10721 24641
rect 10773 24629 10799 24641
rect 10851 24629 11152 24641
rect 9931 24589 10666 24629
rect 9762 24577 10666 24589
rect 10722 24577 10747 24589
rect 10803 24577 10828 24589
rect 9762 24525 9801 24577
rect 9853 24525 9879 24577
rect 9931 24573 10666 24577
rect 10884 24573 10909 24629
rect 10965 24573 10990 24629
rect 11046 24573 11071 24629
rect 11127 24573 11152 24629
rect 11848 24589 12561 24641
rect 12613 24589 12639 24641
rect 12691 24589 14858 24641
rect 11848 24577 14858 24589
rect 9931 24549 10721 24573
rect 10773 24549 10799 24573
rect 10851 24549 11152 24573
rect 9931 24525 10666 24549
rect 9762 24513 10666 24525
rect 10722 24513 10747 24525
rect 10803 24513 10828 24525
rect 9762 24461 9801 24513
rect 9853 24461 9879 24513
rect 9931 24493 10666 24513
rect 10884 24493 10909 24549
rect 10965 24493 10990 24549
rect 11046 24493 11071 24549
rect 11127 24493 11152 24549
rect 11848 24525 12561 24577
rect 12613 24525 12639 24577
rect 12691 24525 14858 24577
rect 11848 24513 14858 24525
rect 9931 24469 10721 24493
rect 10773 24469 10799 24493
rect 10851 24469 11152 24493
rect 9931 24461 10666 24469
rect 9762 24449 10666 24461
rect 10722 24449 10747 24461
rect 10803 24449 10828 24461
rect 9762 24397 9801 24449
rect 9853 24397 9879 24449
rect 9931 24413 10666 24449
rect 10884 24413 10909 24469
rect 10965 24413 10990 24469
rect 11046 24413 11071 24469
rect 11127 24413 11152 24469
rect 11848 24461 12561 24513
rect 12613 24461 12639 24513
rect 12691 24461 14858 24513
rect 11848 24449 14858 24461
rect 9931 24397 10721 24413
rect 10773 24397 10799 24413
rect 10851 24397 11152 24413
rect 11848 24397 12561 24449
rect 12613 24397 12639 24449
rect 12691 24397 14858 24449
rect 9762 24389 11152 24397
rect 9762 24385 10666 24389
rect 10722 24385 10747 24389
rect 10803 24385 10828 24389
rect 9762 24333 9801 24385
rect 9853 24333 9879 24385
rect 9931 24333 10666 24385
rect 10884 24333 10909 24389
rect 10965 24333 10990 24389
rect 11046 24333 11071 24389
rect 11127 24333 11152 24389
rect 11848 24385 14858 24397
rect 11848 24333 12561 24385
rect 12613 24333 12639 24385
rect 12691 24333 14858 24385
rect 9762 24321 11152 24333
rect 11848 24321 14858 24333
rect 9762 24269 9801 24321
rect 9853 24269 9879 24321
rect 9931 24309 10721 24321
rect 10773 24309 10799 24321
rect 10851 24309 11152 24321
rect 9931 24269 10666 24309
rect 9762 24257 10666 24269
rect 10722 24257 10747 24269
rect 10803 24257 10828 24269
rect 9762 24205 9801 24257
rect 9853 24205 9879 24257
rect 9931 24253 10666 24257
rect 10884 24253 10909 24309
rect 10965 24253 10990 24309
rect 11046 24253 11071 24309
rect 11127 24253 11152 24309
rect 11848 24269 12561 24321
rect 12613 24269 12639 24321
rect 12691 24269 14858 24321
rect 11848 24257 14858 24269
rect 9931 24229 10721 24253
rect 10773 24229 10799 24253
rect 10851 24229 11152 24253
rect 9931 24205 10666 24229
rect 9762 24193 10666 24205
rect 10722 24193 10747 24205
rect 10803 24193 10828 24205
rect 9762 24141 9801 24193
rect 9853 24141 9879 24193
rect 9931 24173 10666 24193
rect 10884 24173 10909 24229
rect 10965 24173 10990 24229
rect 11046 24173 11071 24229
rect 11127 24173 11152 24229
rect 11848 24205 12561 24257
rect 12613 24205 12639 24257
rect 12691 24205 14858 24257
rect 11848 24193 14858 24205
rect 9931 24149 10721 24173
rect 10773 24149 10799 24173
rect 10851 24149 11152 24173
rect 9931 24141 10666 24149
rect 9762 24129 10666 24141
rect 10722 24129 10747 24141
rect 10803 24129 10828 24141
rect 9762 24077 9801 24129
rect 9853 24077 9879 24129
rect 9931 24093 10666 24129
rect 10884 24093 10909 24149
rect 10965 24093 10990 24149
rect 11046 24093 11071 24149
rect 11127 24093 11152 24149
rect 11848 24141 12561 24193
rect 12613 24141 12639 24193
rect 12691 24141 14858 24193
rect 11848 24129 14858 24141
rect 9931 24077 10721 24093
rect 10773 24077 10799 24093
rect 10851 24077 11152 24093
rect 11848 24077 12561 24129
rect 12613 24077 12639 24129
rect 12691 24077 14858 24129
rect 9762 24069 11152 24077
rect 9762 24064 10666 24069
rect 10722 24064 10747 24069
rect 10803 24064 10828 24069
rect 9762 24012 9801 24064
rect 9853 24012 9879 24064
rect 9931 24013 10666 24064
rect 10884 24013 10909 24069
rect 10965 24013 10990 24069
rect 11046 24013 11071 24069
rect 11127 24013 11152 24069
rect 11848 24064 14858 24077
rect 9931 24012 10721 24013
rect 10773 24012 10799 24013
rect 10851 24012 11152 24013
rect 11848 24012 12561 24064
rect 12613 24012 12639 24064
rect 12691 24012 14858 24064
rect 9762 23999 11152 24012
rect 11848 23999 14858 24012
rect 9762 23947 9801 23999
rect 9853 23947 9879 23999
rect 9931 23989 10721 23999
rect 10773 23989 10799 23999
rect 10851 23989 11152 23999
rect 9931 23947 10666 23989
rect 9762 23934 10666 23947
rect 10722 23934 10747 23947
rect 10803 23934 10828 23947
rect 9762 23882 9801 23934
rect 9853 23882 9879 23934
rect 9931 23933 10666 23934
rect 10884 23933 10909 23989
rect 10965 23933 10990 23989
rect 11046 23933 11071 23989
rect 11127 23933 11152 23989
rect 11848 23947 12561 23999
rect 12613 23947 12639 23999
rect 12691 23947 14858 23999
rect 11848 23934 14858 23947
rect 9931 23909 10721 23933
rect 10773 23909 10799 23933
rect 10851 23909 11152 23933
rect 9931 23882 10666 23909
rect 9762 23869 10666 23882
rect 10722 23869 10747 23882
rect 10803 23869 10828 23882
rect 9762 23817 9801 23869
rect 9853 23817 9879 23869
rect 9931 23853 10666 23869
rect 10884 23853 10909 23909
rect 10965 23853 10990 23909
rect 11046 23853 11071 23909
rect 11127 23853 11152 23909
rect 11848 23882 12561 23934
rect 12613 23882 12639 23934
rect 12691 23882 14858 23934
rect 11848 23869 14858 23882
rect 9931 23829 10721 23853
rect 10773 23829 10799 23853
rect 10851 23829 11152 23853
rect 9931 23817 10666 23829
rect 9762 23804 10666 23817
rect 10722 23804 10747 23817
rect 10803 23804 10828 23817
rect 9762 23752 9801 23804
rect 9853 23752 9879 23804
rect 9931 23773 10666 23804
rect 10884 23773 10909 23829
rect 10965 23773 10990 23829
rect 11046 23773 11071 23829
rect 11127 23773 11152 23829
rect 11848 23817 12561 23869
rect 12613 23817 12639 23869
rect 12691 23817 14858 23869
rect 11848 23804 14858 23817
rect 9931 23752 10721 23773
rect 10773 23752 10799 23773
rect 10851 23752 11152 23773
rect 11848 23752 12561 23804
rect 12613 23752 12639 23804
rect 12691 23752 14858 23804
rect 9762 23749 11152 23752
rect 9762 23739 10666 23749
rect 10722 23739 10747 23749
rect 10803 23739 10828 23749
rect 9762 23687 9801 23739
rect 9853 23687 9879 23739
rect 9931 23693 10666 23739
rect 10884 23693 10909 23749
rect 10965 23693 10990 23749
rect 11046 23693 11071 23749
rect 11127 23693 11152 23749
rect 11848 23739 14858 23752
rect 9931 23687 10721 23693
rect 10773 23687 10799 23693
rect 10851 23687 11152 23693
rect 11848 23687 12561 23739
rect 12613 23687 12639 23739
rect 12691 23687 14858 23739
rect 9762 23674 11152 23687
rect 11848 23674 14858 23687
rect 9762 23622 9801 23674
rect 9853 23622 9879 23674
rect 9931 23669 10721 23674
rect 10773 23669 10799 23674
rect 10851 23669 11152 23674
rect 9931 23622 10666 23669
rect 9762 23613 10666 23622
rect 10722 23613 10747 23622
rect 10803 23613 10828 23622
rect 10884 23613 10909 23669
rect 10965 23613 10990 23669
rect 11046 23613 11071 23669
rect 11127 23613 11152 23669
rect 11848 23622 12561 23674
rect 12613 23622 12639 23674
rect 12691 23622 14858 23674
rect 9762 23609 11152 23613
rect 11848 23609 14858 23622
rect 9762 23557 9801 23609
rect 9853 23557 9879 23609
rect 9931 23589 10721 23609
rect 10773 23589 10799 23609
rect 10851 23589 11152 23609
rect 9931 23557 10666 23589
rect 9762 23544 10666 23557
rect 10722 23544 10747 23557
rect 10803 23544 10828 23557
rect 9762 23492 9801 23544
rect 9853 23492 9879 23544
rect 9931 23533 10666 23544
rect 10884 23533 10909 23589
rect 10965 23533 10990 23589
rect 11046 23533 11071 23589
rect 11127 23533 11152 23589
rect 11848 23557 12561 23609
rect 12613 23557 12639 23609
rect 12691 23557 14858 23609
rect 11848 23544 14858 23557
rect 9931 23509 10721 23533
rect 10773 23509 10799 23533
rect 10851 23509 11152 23533
rect 9931 23492 10666 23509
rect 9762 23479 10666 23492
rect 10722 23479 10747 23492
rect 10803 23479 10828 23492
rect 9762 23427 9801 23479
rect 9853 23427 9879 23479
rect 9931 23453 10666 23479
rect 10884 23453 10909 23509
rect 10965 23453 10990 23509
rect 11046 23453 11071 23509
rect 11127 23453 11152 23509
rect 11848 23492 12561 23544
rect 12613 23492 12639 23544
rect 12691 23492 14858 23544
rect 11848 23479 14858 23492
rect 9931 23429 10721 23453
rect 10773 23429 10799 23453
rect 10851 23429 11152 23453
rect 9931 23427 10666 23429
rect 9762 23414 10666 23427
rect 10722 23414 10747 23427
rect 10803 23414 10828 23427
rect 9762 23362 9801 23414
rect 9853 23362 9879 23414
rect 9931 23373 10666 23414
rect 10884 23373 10909 23429
rect 10965 23373 10990 23429
rect 11046 23373 11071 23429
rect 11127 23373 11152 23429
rect 11848 23427 12561 23479
rect 12613 23427 12639 23479
rect 12691 23427 14858 23479
rect 11848 23414 14858 23427
rect 9931 23362 10721 23373
rect 10773 23362 10799 23373
rect 10851 23362 11152 23373
rect 11848 23362 12561 23414
rect 12613 23362 12639 23414
rect 12691 23362 14858 23414
rect 9762 23349 11152 23362
rect 11848 23349 14858 23362
rect 9762 23297 9801 23349
rect 9853 23297 9879 23349
rect 9931 23297 10666 23349
rect 9762 23293 10666 23297
rect 10722 23293 10747 23297
rect 10803 23293 10828 23297
rect 10884 23293 10909 23349
rect 10965 23293 10990 23349
rect 11046 23293 11071 23349
rect 11127 23293 11152 23349
rect 11848 23297 12561 23349
rect 12613 23297 12639 23349
rect 12691 23297 14858 23349
rect 11848 23293 14858 23297
rect 4964 23291 14858 23293
rect 3441 23282 3733 23291
rect 3441 23230 3456 23282
rect 3508 23254 3733 23282
rect 3508 23253 3551 23254
tri 3551 23253 3552 23254 nw
tri 3684 23253 3685 23254 ne
rect 3685 23253 3733 23254
tri 3733 23253 3771 23291 sw
rect 3508 23230 3521 23253
rect 3441 23223 3521 23230
tri 3521 23223 3551 23253 nw
tri 3685 23223 3715 23253 ne
rect 3715 23223 3771 23253
tri 3771 23223 3801 23253 sw
tri 3715 23220 3718 23223 ne
rect 3718 23220 3801 23223
tri 3718 23213 3725 23220 ne
rect 3725 23213 3801 23220
tri 3801 23213 3811 23223 sw
tri 2824 22496 3541 23213 sw
tri 3725 23167 3771 23213 ne
rect 3771 23167 3811 23213
tri 3811 23167 3857 23213 sw
tri 3771 23081 3857 23167 ne
tri 3857 23081 3943 23167 sw
tri 3857 22995 3943 23081 ne
tri 3943 22995 4029 23081 sw
tri 3943 22943 3995 22995 ne
rect 3995 22943 4783 22995
rect 4835 22943 4841 22995
tri 4733 22931 4745 22943 ne
rect 4745 22931 4841 22943
tri 4745 22899 4777 22931 ne
rect 4777 22879 4783 22931
rect 4835 22879 4841 22931
tri 11495 22564 12222 23291 ne
rect 187 22494 11341 22496
rect 187 22438 3109 22494
rect 3165 22438 3190 22494
rect 3246 22438 3271 22494
rect 3327 22438 3352 22494
rect 3408 22438 3433 22494
rect 3489 22438 3514 22494
rect 187 22414 3514 22438
rect 187 22358 3109 22414
rect 3165 22358 3190 22414
rect 3246 22358 3271 22414
rect 3327 22358 3352 22414
rect 3408 22358 3433 22414
rect 3489 22358 3514 22414
rect 187 22334 3514 22358
rect 187 22278 3109 22334
rect 3165 22278 3190 22334
rect 3246 22278 3271 22334
rect 3327 22278 3352 22334
rect 3408 22278 3433 22334
rect 3489 22278 3514 22334
rect 187 22254 3514 22278
rect 187 22198 3109 22254
rect 3165 22198 3190 22254
rect 3246 22198 3271 22254
rect 3327 22198 3352 22254
rect 3408 22198 3433 22254
rect 3489 22198 3514 22254
rect 187 22174 3514 22198
rect 187 22118 3109 22174
rect 3165 22118 3190 22174
rect 3246 22118 3271 22174
rect 3327 22118 3352 22174
rect 3408 22118 3433 22174
rect 3489 22118 3514 22174
rect 187 22094 3514 22118
rect 187 22038 3109 22094
rect 3165 22038 3190 22094
rect 3246 22038 3271 22094
rect 3327 22038 3352 22094
rect 3408 22038 3433 22094
rect 3489 22038 3514 22094
rect 187 22014 3514 22038
rect 187 21958 3109 22014
rect 3165 21958 3190 22014
rect 3246 21958 3271 22014
rect 3327 21958 3352 22014
rect 3408 21958 3433 22014
rect 3489 21958 3514 22014
rect 187 21934 3514 21958
rect 187 21878 3109 21934
rect 3165 21878 3190 21934
rect 3246 21878 3271 21934
rect 3327 21878 3352 21934
rect 3408 21878 3433 21934
rect 3489 21878 3514 21934
rect 187 21854 3514 21878
rect 187 21798 3109 21854
rect 3165 21798 3190 21854
rect 3246 21798 3271 21854
rect 3327 21798 3352 21854
rect 3408 21798 3433 21854
rect 3489 21798 3514 21854
rect 187 21774 3514 21798
rect 187 21718 3109 21774
rect 3165 21718 3190 21774
rect 3246 21718 3271 21774
rect 3327 21718 3352 21774
rect 3408 21718 3433 21774
rect 3489 21718 3514 21774
rect 187 21694 3514 21718
rect 187 21638 3109 21694
rect 3165 21638 3190 21694
rect 3246 21638 3271 21694
rect 3327 21638 3352 21694
rect 3408 21638 3433 21694
rect 3489 21638 3514 21694
rect 187 21614 3514 21638
rect 187 21558 3109 21614
rect 3165 21558 3190 21614
rect 3246 21558 3271 21614
rect 3327 21558 3352 21614
rect 3408 21558 3433 21614
rect 3489 21558 3514 21614
rect 187 21534 3514 21558
rect 187 21478 3109 21534
rect 3165 21478 3190 21534
rect 3246 21478 3271 21534
rect 3327 21478 3352 21534
rect 3408 21478 3433 21534
rect 3489 21478 3514 21534
rect 187 21454 3514 21478
rect 187 21398 3109 21454
rect 3165 21398 3190 21454
rect 3246 21398 3271 21454
rect 3327 21398 3352 21454
rect 3408 21398 3433 21454
rect 3489 21398 3514 21454
rect 187 21374 3514 21398
rect 187 21318 3109 21374
rect 3165 21318 3190 21374
rect 3246 21318 3271 21374
rect 3327 21318 3352 21374
rect 3408 21318 3433 21374
rect 3489 21318 3514 21374
rect 187 21294 3514 21318
rect 187 21238 3109 21294
rect 3165 21238 3190 21294
rect 3246 21238 3271 21294
rect 3327 21238 3352 21294
rect 3408 21238 3433 21294
rect 3489 21238 3514 21294
rect 187 21214 3514 21238
rect 187 21158 3109 21214
rect 3165 21158 3190 21214
rect 3246 21158 3271 21214
rect 3327 21158 3352 21214
rect 3408 21158 3433 21214
rect 3489 21158 3514 21214
rect 187 21134 3514 21158
rect 187 21078 3109 21134
rect 3165 21078 3190 21134
rect 3246 21078 3271 21134
rect 3327 21078 3352 21134
rect 3408 21078 3433 21134
rect 3489 21078 3514 21134
rect 187 21054 3514 21078
rect 187 20998 3109 21054
rect 3165 20998 3190 21054
rect 3246 20998 3271 21054
rect 3327 20998 3352 21054
rect 3408 20998 3433 21054
rect 3489 20998 3514 21054
rect 187 20974 3514 20998
rect 187 20918 3109 20974
rect 3165 20918 3190 20974
rect 3246 20918 3271 20974
rect 3327 20918 3352 20974
rect 3408 20918 3433 20974
rect 3489 20918 3514 20974
rect 187 20894 3514 20918
rect 187 20838 3109 20894
rect 3165 20838 3190 20894
rect 3246 20838 3271 20894
rect 3327 20838 3352 20894
rect 3408 20838 3433 20894
rect 3489 20838 3514 20894
rect 187 20814 3514 20838
rect 187 20758 3109 20814
rect 3165 20758 3190 20814
rect 3246 20758 3271 20814
rect 3327 20758 3352 20814
rect 3408 20758 3433 20814
rect 3489 20758 3514 20814
rect 4290 22490 5195 22494
rect 4290 22438 4777 22490
rect 4829 22438 4849 22490
rect 4901 22438 5195 22490
rect 5251 22438 5276 22494
rect 5332 22438 5357 22494
rect 5413 22438 5438 22494
rect 5494 22438 5519 22494
rect 5575 22438 5600 22494
rect 6376 22490 11341 22494
rect 6376 22438 6552 22490
rect 6604 22438 6620 22490
rect 6672 22438 6688 22490
rect 6740 22438 7472 22490
rect 7524 22438 7540 22490
rect 7592 22438 7608 22490
rect 7660 22438 8392 22490
rect 8444 22438 8460 22490
rect 8512 22438 8528 22490
rect 8580 22438 9312 22490
rect 9364 22438 9380 22490
rect 9432 22438 9448 22490
rect 9500 22438 10232 22490
rect 10284 22438 10300 22490
rect 10352 22438 10368 22490
rect 10420 22438 11152 22490
rect 11204 22438 11220 22490
rect 11272 22438 11288 22490
rect 11340 22438 11341 22490
rect 4290 22426 5600 22438
rect 6376 22426 11341 22438
rect 4290 22374 4777 22426
rect 4829 22374 4849 22426
rect 4901 22414 5600 22426
rect 4901 22374 5195 22414
rect 4290 22362 5195 22374
rect 4290 22310 4777 22362
rect 4829 22310 4849 22362
rect 4901 22358 5195 22362
rect 5251 22358 5276 22414
rect 5332 22358 5357 22414
rect 5413 22358 5438 22414
rect 5494 22358 5519 22414
rect 5575 22358 5600 22414
rect 6376 22374 6552 22426
rect 6604 22374 6620 22426
rect 6672 22374 6688 22426
rect 6740 22374 7472 22426
rect 7524 22374 7540 22426
rect 7592 22374 7608 22426
rect 7660 22374 8392 22426
rect 8444 22374 8460 22426
rect 8512 22374 8528 22426
rect 8580 22374 9312 22426
rect 9364 22374 9380 22426
rect 9432 22374 9448 22426
rect 9500 22374 10232 22426
rect 10284 22374 10300 22426
rect 10352 22374 10368 22426
rect 10420 22374 11152 22426
rect 11204 22374 11220 22426
rect 11272 22374 11288 22426
rect 11340 22374 11341 22426
rect 6376 22362 11341 22374
rect 4901 22334 5600 22358
rect 4901 22310 5195 22334
rect 4290 22298 5195 22310
rect 4290 22246 4777 22298
rect 4829 22246 4849 22298
rect 4901 22278 5195 22298
rect 5251 22278 5276 22334
rect 5332 22278 5357 22334
rect 5413 22278 5438 22334
rect 5494 22278 5519 22334
rect 5575 22278 5600 22334
rect 6376 22310 6552 22362
rect 6604 22310 6620 22362
rect 6672 22310 6688 22362
rect 6740 22310 7472 22362
rect 7524 22310 7540 22362
rect 7592 22310 7608 22362
rect 7660 22310 8392 22362
rect 8444 22310 8460 22362
rect 8512 22310 8528 22362
rect 8580 22310 9312 22362
rect 9364 22310 9380 22362
rect 9432 22310 9448 22362
rect 9500 22310 10232 22362
rect 10284 22310 10300 22362
rect 10352 22310 10368 22362
rect 10420 22310 11152 22362
rect 11204 22310 11220 22362
rect 11272 22310 11288 22362
rect 11340 22310 11341 22362
rect 6376 22298 11341 22310
rect 4901 22254 5600 22278
rect 4901 22246 5195 22254
rect 4290 22234 5195 22246
rect 4290 22182 4777 22234
rect 4829 22182 4849 22234
rect 4901 22198 5195 22234
rect 5251 22198 5276 22254
rect 5332 22198 5357 22254
rect 5413 22198 5438 22254
rect 5494 22198 5519 22254
rect 5575 22198 5600 22254
rect 6376 22246 6552 22298
rect 6604 22246 6620 22298
rect 6672 22246 6688 22298
rect 6740 22246 7472 22298
rect 7524 22246 7540 22298
rect 7592 22246 7608 22298
rect 7660 22246 8392 22298
rect 8444 22246 8460 22298
rect 8512 22246 8528 22298
rect 8580 22246 9312 22298
rect 9364 22246 9380 22298
rect 9432 22246 9448 22298
rect 9500 22246 10232 22298
rect 10284 22246 10300 22298
rect 10352 22246 10368 22298
rect 10420 22246 11152 22298
rect 11204 22246 11220 22298
rect 11272 22246 11288 22298
rect 11340 22246 11341 22298
rect 6376 22234 11341 22246
rect 4901 22182 5600 22198
rect 6376 22182 6552 22234
rect 6604 22182 6620 22234
rect 6672 22182 6688 22234
rect 6740 22182 7472 22234
rect 7524 22182 7540 22234
rect 7592 22182 7608 22234
rect 7660 22182 8392 22234
rect 8444 22182 8460 22234
rect 8512 22182 8528 22234
rect 8580 22182 9312 22234
rect 9364 22182 9380 22234
rect 9432 22182 9448 22234
rect 9500 22182 10232 22234
rect 10284 22182 10300 22234
rect 10352 22182 10368 22234
rect 10420 22182 11152 22234
rect 11204 22182 11220 22234
rect 11272 22182 11288 22234
rect 11340 22182 11341 22234
rect 4290 22174 5600 22182
rect 4290 22170 5195 22174
rect 4290 22118 4777 22170
rect 4829 22118 4849 22170
rect 4901 22118 5195 22170
rect 5251 22118 5276 22174
rect 5332 22118 5357 22174
rect 5413 22118 5438 22174
rect 5494 22118 5519 22174
rect 5575 22118 5600 22174
rect 6376 22170 11341 22182
rect 6376 22118 6552 22170
rect 6604 22118 6620 22170
rect 6672 22118 6688 22170
rect 6740 22118 7472 22170
rect 7524 22118 7540 22170
rect 7592 22118 7608 22170
rect 7660 22118 8392 22170
rect 8444 22118 8460 22170
rect 8512 22118 8528 22170
rect 8580 22118 9312 22170
rect 9364 22118 9380 22170
rect 9432 22118 9448 22170
rect 9500 22118 10232 22170
rect 10284 22118 10300 22170
rect 10352 22118 10368 22170
rect 10420 22118 11152 22170
rect 11204 22118 11220 22170
rect 11272 22118 11288 22170
rect 11340 22118 11341 22170
rect 4290 22106 5600 22118
rect 6376 22106 11341 22118
rect 4290 22054 4777 22106
rect 4829 22054 4849 22106
rect 4901 22094 5600 22106
rect 4901 22054 5195 22094
rect 4290 22042 5195 22054
rect 4290 21990 4777 22042
rect 4829 21990 4849 22042
rect 4901 22038 5195 22042
rect 5251 22038 5276 22094
rect 5332 22038 5357 22094
rect 5413 22038 5438 22094
rect 5494 22038 5519 22094
rect 5575 22038 5600 22094
rect 6376 22054 6552 22106
rect 6604 22054 6620 22106
rect 6672 22054 6688 22106
rect 6740 22054 7472 22106
rect 7524 22054 7540 22106
rect 7592 22054 7608 22106
rect 7660 22054 8392 22106
rect 8444 22054 8460 22106
rect 8512 22054 8528 22106
rect 8580 22054 9312 22106
rect 9364 22054 9380 22106
rect 9432 22054 9448 22106
rect 9500 22054 10232 22106
rect 10284 22054 10300 22106
rect 10352 22054 10368 22106
rect 10420 22054 11152 22106
rect 11204 22054 11220 22106
rect 11272 22054 11288 22106
rect 11340 22054 11341 22106
rect 6376 22042 11341 22054
rect 4901 22014 5600 22038
rect 4901 21990 5195 22014
rect 4290 21978 5195 21990
rect 4290 21926 4777 21978
rect 4829 21926 4849 21978
rect 4901 21958 5195 21978
rect 5251 21958 5276 22014
rect 5332 21958 5357 22014
rect 5413 21958 5438 22014
rect 5494 21958 5519 22014
rect 5575 21958 5600 22014
rect 6376 21990 6552 22042
rect 6604 21990 6620 22042
rect 6672 21990 6688 22042
rect 6740 21990 7472 22042
rect 7524 21990 7540 22042
rect 7592 21990 7608 22042
rect 7660 21990 8392 22042
rect 8444 21990 8460 22042
rect 8512 21990 8528 22042
rect 8580 21990 9312 22042
rect 9364 21990 9380 22042
rect 9432 21990 9448 22042
rect 9500 21990 10232 22042
rect 10284 21990 10300 22042
rect 10352 21990 10368 22042
rect 10420 21990 11152 22042
rect 11204 21990 11220 22042
rect 11272 21990 11288 22042
rect 11340 21990 11341 22042
rect 6376 21978 11341 21990
rect 4901 21934 5600 21958
rect 4901 21926 5195 21934
rect 4290 21914 5195 21926
rect 4290 21862 4777 21914
rect 4829 21862 4849 21914
rect 4901 21878 5195 21914
rect 5251 21878 5276 21934
rect 5332 21878 5357 21934
rect 5413 21878 5438 21934
rect 5494 21878 5519 21934
rect 5575 21878 5600 21934
rect 6376 21926 6552 21978
rect 6604 21926 6620 21978
rect 6672 21926 6688 21978
rect 6740 21926 7472 21978
rect 7524 21926 7540 21978
rect 7592 21926 7608 21978
rect 7660 21926 8392 21978
rect 8444 21926 8460 21978
rect 8512 21926 8528 21978
rect 8580 21926 9312 21978
rect 9364 21926 9380 21978
rect 9432 21926 9448 21978
rect 9500 21926 10232 21978
rect 10284 21926 10300 21978
rect 10352 21926 10368 21978
rect 10420 21926 11152 21978
rect 11204 21926 11220 21978
rect 11272 21926 11288 21978
rect 11340 21926 11341 21978
rect 6376 21914 11341 21926
rect 4901 21862 5600 21878
rect 6376 21862 6552 21914
rect 6604 21862 6620 21914
rect 6672 21862 6688 21914
rect 6740 21862 7472 21914
rect 7524 21862 7540 21914
rect 7592 21862 7608 21914
rect 7660 21862 8392 21914
rect 8444 21862 8460 21914
rect 8512 21862 8528 21914
rect 8580 21862 9312 21914
rect 9364 21862 9380 21914
rect 9432 21862 9448 21914
rect 9500 21862 10232 21914
rect 10284 21862 10300 21914
rect 10352 21862 10368 21914
rect 10420 21862 11152 21914
rect 11204 21862 11220 21914
rect 11272 21862 11288 21914
rect 11340 21862 11341 21914
rect 4290 21854 5600 21862
rect 4290 21850 5195 21854
rect 4290 21798 4777 21850
rect 4829 21798 4849 21850
rect 4901 21798 5195 21850
rect 5251 21798 5276 21854
rect 5332 21798 5357 21854
rect 5413 21798 5438 21854
rect 5494 21798 5519 21854
rect 5575 21798 5600 21854
rect 6376 21850 11341 21862
rect 6376 21798 6552 21850
rect 6604 21798 6620 21850
rect 6672 21798 6688 21850
rect 6740 21798 7472 21850
rect 7524 21798 7540 21850
rect 7592 21798 7608 21850
rect 7660 21798 8392 21850
rect 8444 21798 8460 21850
rect 8512 21798 8528 21850
rect 8580 21798 9312 21850
rect 9364 21798 9380 21850
rect 9432 21798 9448 21850
rect 9500 21798 10232 21850
rect 10284 21798 10300 21850
rect 10352 21798 10368 21850
rect 10420 21798 11152 21850
rect 11204 21798 11220 21850
rect 11272 21798 11288 21850
rect 11340 21798 11341 21850
rect 4290 21786 5600 21798
rect 6376 21786 11341 21798
rect 4290 21734 4777 21786
rect 4829 21734 4849 21786
rect 4901 21774 5600 21786
rect 4901 21734 5195 21774
rect 4290 21722 5195 21734
rect 4290 21670 4777 21722
rect 4829 21670 4849 21722
rect 4901 21718 5195 21722
rect 5251 21718 5276 21774
rect 5332 21718 5357 21774
rect 5413 21718 5438 21774
rect 5494 21718 5519 21774
rect 5575 21718 5600 21774
rect 6376 21734 6552 21786
rect 6604 21734 6620 21786
rect 6672 21734 6688 21786
rect 6740 21734 7472 21786
rect 7524 21734 7540 21786
rect 7592 21734 7608 21786
rect 7660 21734 8392 21786
rect 8444 21734 8460 21786
rect 8512 21734 8528 21786
rect 8580 21734 9312 21786
rect 9364 21734 9380 21786
rect 9432 21734 9448 21786
rect 9500 21734 10232 21786
rect 10284 21734 10300 21786
rect 10352 21734 10368 21786
rect 10420 21734 11152 21786
rect 11204 21734 11220 21786
rect 11272 21734 11288 21786
rect 11340 21734 11341 21786
rect 6376 21722 11341 21734
rect 4901 21694 5600 21718
rect 4901 21670 5195 21694
rect 4290 21658 5195 21670
rect 4290 21606 4777 21658
rect 4829 21606 4849 21658
rect 4901 21638 5195 21658
rect 5251 21638 5276 21694
rect 5332 21638 5357 21694
rect 5413 21638 5438 21694
rect 5494 21638 5519 21694
rect 5575 21638 5600 21694
rect 6376 21670 6552 21722
rect 6604 21670 6620 21722
rect 6672 21670 6688 21722
rect 6740 21670 7472 21722
rect 7524 21670 7540 21722
rect 7592 21670 7608 21722
rect 7660 21670 8392 21722
rect 8444 21670 8460 21722
rect 8512 21670 8528 21722
rect 8580 21670 9312 21722
rect 9364 21670 9380 21722
rect 9432 21670 9448 21722
rect 9500 21670 10232 21722
rect 10284 21670 10300 21722
rect 10352 21670 10368 21722
rect 10420 21670 11152 21722
rect 11204 21670 11220 21722
rect 11272 21670 11288 21722
rect 11340 21670 11341 21722
rect 6376 21658 11341 21670
rect 4901 21614 5600 21638
rect 4901 21606 5195 21614
rect 4290 21594 5195 21606
rect 4290 21542 4777 21594
rect 4829 21542 4849 21594
rect 4901 21558 5195 21594
rect 5251 21558 5276 21614
rect 5332 21558 5357 21614
rect 5413 21558 5438 21614
rect 5494 21558 5519 21614
rect 5575 21558 5600 21614
rect 6376 21606 6552 21658
rect 6604 21606 6620 21658
rect 6672 21606 6688 21658
rect 6740 21606 7472 21658
rect 7524 21606 7540 21658
rect 7592 21606 7608 21658
rect 7660 21606 8392 21658
rect 8444 21606 8460 21658
rect 8512 21606 8528 21658
rect 8580 21606 9312 21658
rect 9364 21606 9380 21658
rect 9432 21606 9448 21658
rect 9500 21606 10232 21658
rect 10284 21606 10300 21658
rect 10352 21606 10368 21658
rect 10420 21606 11152 21658
rect 11204 21606 11220 21658
rect 11272 21606 11288 21658
rect 11340 21606 11341 21658
rect 6376 21594 11341 21606
rect 4901 21542 5600 21558
rect 6376 21542 6552 21594
rect 6604 21542 6620 21594
rect 6672 21542 6688 21594
rect 6740 21542 7472 21594
rect 7524 21542 7540 21594
rect 7592 21542 7608 21594
rect 7660 21542 8392 21594
rect 8444 21542 8460 21594
rect 8512 21542 8528 21594
rect 8580 21542 9312 21594
rect 9364 21542 9380 21594
rect 9432 21542 9448 21594
rect 9500 21542 10232 21594
rect 10284 21542 10300 21594
rect 10352 21542 10368 21594
rect 10420 21542 11152 21594
rect 11204 21542 11220 21594
rect 11272 21542 11288 21594
rect 11340 21542 11341 21594
rect 4290 21534 5600 21542
rect 4290 21529 5195 21534
rect 4290 21477 4777 21529
rect 4829 21477 4849 21529
rect 4901 21478 5195 21529
rect 5251 21478 5276 21534
rect 5332 21478 5357 21534
rect 5413 21478 5438 21534
rect 5494 21478 5519 21534
rect 5575 21478 5600 21534
rect 6376 21529 11341 21542
rect 4901 21477 5600 21478
rect 6376 21477 6552 21529
rect 6604 21477 6620 21529
rect 6672 21477 6688 21529
rect 6740 21477 7472 21529
rect 7524 21477 7540 21529
rect 7592 21477 7608 21529
rect 7660 21477 8392 21529
rect 8444 21477 8460 21529
rect 8512 21477 8528 21529
rect 8580 21477 9312 21529
rect 9364 21477 9380 21529
rect 9432 21477 9448 21529
rect 9500 21477 10232 21529
rect 10284 21477 10300 21529
rect 10352 21477 10368 21529
rect 10420 21477 11152 21529
rect 11204 21477 11220 21529
rect 11272 21477 11288 21529
rect 11340 21477 11341 21529
rect 4290 21464 5600 21477
rect 6376 21464 11341 21477
rect 4290 21412 4777 21464
rect 4829 21412 4849 21464
rect 4901 21454 5600 21464
rect 4901 21412 5195 21454
rect 4290 21399 5195 21412
rect 4290 21347 4777 21399
rect 4829 21347 4849 21399
rect 4901 21398 5195 21399
rect 5251 21398 5276 21454
rect 5332 21398 5357 21454
rect 5413 21398 5438 21454
rect 5494 21398 5519 21454
rect 5575 21398 5600 21454
rect 6376 21412 6552 21464
rect 6604 21412 6620 21464
rect 6672 21412 6688 21464
rect 6740 21412 7472 21464
rect 7524 21412 7540 21464
rect 7592 21412 7608 21464
rect 7660 21412 8392 21464
rect 8444 21412 8460 21464
rect 8512 21412 8528 21464
rect 8580 21412 9312 21464
rect 9364 21412 9380 21464
rect 9432 21412 9448 21464
rect 9500 21412 10232 21464
rect 10284 21412 10300 21464
rect 10352 21412 10368 21464
rect 10420 21412 11152 21464
rect 11204 21412 11220 21464
rect 11272 21412 11288 21464
rect 11340 21412 11341 21464
rect 6376 21399 11341 21412
rect 4901 21374 5600 21398
rect 4901 21347 5195 21374
rect 4290 21334 5195 21347
rect 4290 21282 4777 21334
rect 4829 21282 4849 21334
rect 4901 21318 5195 21334
rect 5251 21318 5276 21374
rect 5332 21318 5357 21374
rect 5413 21318 5438 21374
rect 5494 21318 5519 21374
rect 5575 21318 5600 21374
rect 6376 21347 6552 21399
rect 6604 21347 6620 21399
rect 6672 21347 6688 21399
rect 6740 21347 7472 21399
rect 7524 21347 7540 21399
rect 7592 21347 7608 21399
rect 7660 21347 8392 21399
rect 8444 21347 8460 21399
rect 8512 21347 8528 21399
rect 8580 21347 9312 21399
rect 9364 21347 9380 21399
rect 9432 21347 9448 21399
rect 9500 21347 10232 21399
rect 10284 21347 10300 21399
rect 10352 21347 10368 21399
rect 10420 21347 11152 21399
rect 11204 21347 11220 21399
rect 11272 21347 11288 21399
rect 11340 21347 11341 21399
rect 6376 21334 11341 21347
rect 4901 21294 5600 21318
rect 4901 21282 5195 21294
rect 4290 21269 5195 21282
rect 4290 21217 4777 21269
rect 4829 21217 4849 21269
rect 4901 21238 5195 21269
rect 5251 21238 5276 21294
rect 5332 21238 5357 21294
rect 5413 21238 5438 21294
rect 5494 21238 5519 21294
rect 5575 21238 5600 21294
rect 6376 21282 6552 21334
rect 6604 21282 6620 21334
rect 6672 21282 6688 21334
rect 6740 21282 7472 21334
rect 7524 21282 7540 21334
rect 7592 21282 7608 21334
rect 7660 21282 8392 21334
rect 8444 21282 8460 21334
rect 8512 21282 8528 21334
rect 8580 21282 9312 21334
rect 9364 21282 9380 21334
rect 9432 21282 9448 21334
rect 9500 21282 10232 21334
rect 10284 21282 10300 21334
rect 10352 21282 10368 21334
rect 10420 21282 11152 21334
rect 11204 21282 11220 21334
rect 11272 21282 11288 21334
rect 11340 21282 11341 21334
rect 6376 21269 11341 21282
rect 4901 21217 5600 21238
rect 6376 21217 6552 21269
rect 6604 21217 6620 21269
rect 6672 21217 6688 21269
rect 6740 21217 7472 21269
rect 7524 21217 7540 21269
rect 7592 21217 7608 21269
rect 7660 21217 8392 21269
rect 8444 21217 8460 21269
rect 8512 21217 8528 21269
rect 8580 21217 9312 21269
rect 9364 21217 9380 21269
rect 9432 21217 9448 21269
rect 9500 21217 10232 21269
rect 10284 21217 10300 21269
rect 10352 21217 10368 21269
rect 10420 21217 11152 21269
rect 11204 21217 11220 21269
rect 11272 21217 11288 21269
rect 11340 21217 11341 21269
rect 4290 21214 5600 21217
rect 4290 21204 5195 21214
rect 4290 21152 4777 21204
rect 4829 21152 4849 21204
rect 4901 21158 5195 21204
rect 5251 21158 5276 21214
rect 5332 21158 5357 21214
rect 5413 21158 5438 21214
rect 5494 21158 5519 21214
rect 5575 21158 5600 21214
rect 6376 21204 11341 21217
rect 4901 21152 5600 21158
rect 6376 21152 6552 21204
rect 6604 21152 6620 21204
rect 6672 21152 6688 21204
rect 6740 21152 7472 21204
rect 7524 21152 7540 21204
rect 7592 21152 7608 21204
rect 7660 21152 8392 21204
rect 8444 21152 8460 21204
rect 8512 21152 8528 21204
rect 8580 21152 9312 21204
rect 9364 21152 9380 21204
rect 9432 21152 9448 21204
rect 9500 21152 10232 21204
rect 10284 21152 10300 21204
rect 10352 21152 10368 21204
rect 10420 21152 11152 21204
rect 11204 21152 11220 21204
rect 11272 21152 11288 21204
rect 11340 21152 11341 21204
rect 4290 21139 5600 21152
rect 6376 21139 11341 21152
rect 4290 21087 4777 21139
rect 4829 21087 4849 21139
rect 4901 21134 5600 21139
rect 4901 21087 5195 21134
rect 4290 21078 5195 21087
rect 5251 21078 5276 21134
rect 5332 21078 5357 21134
rect 5413 21078 5438 21134
rect 5494 21078 5519 21134
rect 5575 21078 5600 21134
rect 6376 21087 6552 21139
rect 6604 21087 6620 21139
rect 6672 21087 6688 21139
rect 6740 21087 7472 21139
rect 7524 21087 7540 21139
rect 7592 21087 7608 21139
rect 7660 21087 8392 21139
rect 8444 21087 8460 21139
rect 8512 21087 8528 21139
rect 8580 21087 9312 21139
rect 9364 21087 9380 21139
rect 9432 21087 9448 21139
rect 9500 21087 10232 21139
rect 10284 21087 10300 21139
rect 10352 21087 10368 21139
rect 10420 21087 11152 21139
rect 11204 21087 11220 21139
rect 11272 21087 11288 21139
rect 11340 21087 11341 21139
rect 4290 21074 5600 21078
rect 6376 21074 11341 21087
rect 4290 21022 4777 21074
rect 4829 21022 4849 21074
rect 4901 21054 5600 21074
rect 4901 21022 5195 21054
rect 4290 21009 5195 21022
rect 4290 20957 4777 21009
rect 4829 20957 4849 21009
rect 4901 20998 5195 21009
rect 5251 20998 5276 21054
rect 5332 20998 5357 21054
rect 5413 20998 5438 21054
rect 5494 20998 5519 21054
rect 5575 20998 5600 21054
rect 6376 21022 6552 21074
rect 6604 21022 6620 21074
rect 6672 21022 6688 21074
rect 6740 21022 7472 21074
rect 7524 21022 7540 21074
rect 7592 21022 7608 21074
rect 7660 21022 8392 21074
rect 8444 21022 8460 21074
rect 8512 21022 8528 21074
rect 8580 21022 9312 21074
rect 9364 21022 9380 21074
rect 9432 21022 9448 21074
rect 9500 21022 10232 21074
rect 10284 21022 10300 21074
rect 10352 21022 10368 21074
rect 10420 21022 11152 21074
rect 11204 21022 11220 21074
rect 11272 21022 11288 21074
rect 11340 21022 11341 21074
rect 6376 21009 11341 21022
rect 4901 20974 5600 20998
rect 4901 20957 5195 20974
rect 4290 20944 5195 20957
rect 4290 20892 4777 20944
rect 4829 20892 4849 20944
rect 4901 20918 5195 20944
rect 5251 20918 5276 20974
rect 5332 20918 5357 20974
rect 5413 20918 5438 20974
rect 5494 20918 5519 20974
rect 5575 20918 5600 20974
rect 6376 20957 6552 21009
rect 6604 20957 6620 21009
rect 6672 20957 6688 21009
rect 6740 20957 7472 21009
rect 7524 20957 7540 21009
rect 7592 20957 7608 21009
rect 7660 20957 8392 21009
rect 8444 20957 8460 21009
rect 8512 20957 8528 21009
rect 8580 20957 9312 21009
rect 9364 20957 9380 21009
rect 9432 20957 9448 21009
rect 9500 20957 10232 21009
rect 10284 20957 10300 21009
rect 10352 20957 10368 21009
rect 10420 20957 11152 21009
rect 11204 20957 11220 21009
rect 11272 20957 11288 21009
rect 11340 20957 11341 21009
rect 6376 20944 11341 20957
rect 4901 20894 5600 20918
rect 4901 20892 5195 20894
rect 4290 20879 5195 20892
rect 4290 20827 4777 20879
rect 4829 20827 4849 20879
rect 4901 20838 5195 20879
rect 5251 20838 5276 20894
rect 5332 20838 5357 20894
rect 5413 20838 5438 20894
rect 5494 20838 5519 20894
rect 5575 20838 5600 20894
rect 6376 20892 6552 20944
rect 6604 20892 6620 20944
rect 6672 20892 6688 20944
rect 6740 20892 7472 20944
rect 7524 20892 7540 20944
rect 7592 20892 7608 20944
rect 7660 20892 8392 20944
rect 8444 20892 8460 20944
rect 8512 20892 8528 20944
rect 8580 20892 9312 20944
rect 9364 20892 9380 20944
rect 9432 20892 9448 20944
rect 9500 20892 10232 20944
rect 10284 20892 10300 20944
rect 10352 20892 10368 20944
rect 10420 20892 11152 20944
rect 11204 20892 11220 20944
rect 11272 20892 11288 20944
rect 11340 20892 11341 20944
rect 6376 20879 11341 20892
rect 4901 20827 5600 20838
rect 6376 20827 6552 20879
rect 6604 20827 6620 20879
rect 6672 20827 6688 20879
rect 6740 20827 7472 20879
rect 7524 20827 7540 20879
rect 7592 20827 7608 20879
rect 7660 20827 8392 20879
rect 8444 20827 8460 20879
rect 8512 20827 8528 20879
rect 8580 20827 9312 20879
rect 9364 20827 9380 20879
rect 9432 20827 9448 20879
rect 9500 20827 10232 20879
rect 10284 20827 10300 20879
rect 10352 20827 10368 20879
rect 10420 20827 11152 20879
rect 11204 20827 11220 20879
rect 11272 20827 11288 20879
rect 11340 20827 11341 20879
rect 4290 20814 5600 20827
rect 6376 20814 11341 20827
rect 4290 20762 4777 20814
rect 4829 20762 4849 20814
rect 4901 20762 5195 20814
rect 4290 20758 5195 20762
rect 5251 20758 5276 20814
rect 5332 20758 5357 20814
rect 5413 20758 5438 20814
rect 5494 20758 5519 20814
rect 5575 20758 5600 20814
rect 6376 20762 6552 20814
rect 6604 20762 6620 20814
rect 6672 20762 6688 20814
rect 6740 20762 7472 20814
rect 7524 20762 7540 20814
rect 7592 20762 7608 20814
rect 7660 20762 8392 20814
rect 8444 20762 8460 20814
rect 8512 20762 8528 20814
rect 8580 20762 9312 20814
rect 9364 20762 9380 20814
rect 9432 20762 9448 20814
rect 9500 20762 10232 20814
rect 10284 20762 10300 20814
rect 10352 20762 10368 20814
rect 10420 20762 11152 20814
rect 11204 20762 11220 20814
rect 11272 20762 11288 20814
rect 11340 20762 11341 20814
rect 6376 20758 11341 20762
rect 187 20756 11341 20758
rect 187 17896 2824 20756
tri 2824 20048 3532 20756 nw
tri 11511 20431 12222 21142 se
rect 12222 20431 14858 23291
rect 4964 20429 14858 20431
rect 4964 20425 7640 20429
rect 4964 20373 5201 20425
rect 5253 20373 5279 20425
rect 5331 20373 6121 20425
rect 6173 20373 6199 20425
rect 6251 20373 7041 20425
rect 7093 20373 7119 20425
rect 7171 20373 7640 20425
rect 7696 20373 7726 20429
rect 7782 20373 7812 20429
rect 7868 20373 7898 20429
rect 7954 20425 7984 20429
rect 8040 20425 8070 20429
rect 7954 20373 7961 20425
rect 8126 20373 8156 20429
rect 8212 20373 8242 20429
rect 8298 20373 8327 20429
rect 8383 20373 8412 20429
rect 8468 20373 8497 20429
rect 8553 20425 9079 20429
rect 8553 20373 8881 20425
rect 8933 20373 8959 20425
rect 9011 20373 9079 20425
rect 9135 20373 9170 20429
rect 9226 20373 9260 20429
rect 9316 20373 9350 20429
rect 9406 20373 9440 20429
rect 9496 20373 9530 20429
rect 9586 20373 9620 20429
rect 9676 20373 9710 20429
rect 9766 20425 14858 20429
rect 9766 20373 9801 20425
rect 9853 20373 9879 20425
rect 9931 20373 10721 20425
rect 10773 20373 10799 20425
rect 10851 20373 11641 20425
rect 11693 20373 11719 20425
rect 11771 20373 12561 20425
rect 12613 20373 12639 20425
rect 12691 20373 14858 20425
rect 4964 20361 14858 20373
rect 4964 20309 5201 20361
rect 5253 20309 5279 20361
rect 5331 20309 6121 20361
rect 6173 20309 6199 20361
rect 6251 20309 7041 20361
rect 7093 20309 7119 20361
rect 7171 20349 7961 20361
rect 8013 20349 8039 20361
rect 8091 20349 8881 20361
rect 7171 20309 7640 20349
rect 4964 20297 7640 20309
rect 4964 20245 5201 20297
rect 5253 20245 5279 20297
rect 5331 20245 6121 20297
rect 6173 20245 6199 20297
rect 6251 20245 7041 20297
rect 7093 20245 7119 20297
rect 7171 20293 7640 20297
rect 7696 20293 7726 20349
rect 7782 20293 7812 20349
rect 7868 20293 7898 20349
rect 7954 20309 7961 20349
rect 7954 20297 7984 20309
rect 8040 20297 8070 20309
rect 7954 20293 7961 20297
rect 8126 20293 8156 20349
rect 8212 20293 8242 20349
rect 8298 20293 8327 20349
rect 8383 20293 8412 20349
rect 8468 20293 8497 20349
rect 8553 20309 8881 20349
rect 8933 20309 8959 20361
rect 9011 20349 9801 20361
rect 9011 20309 9079 20349
rect 8553 20297 9079 20309
rect 8553 20293 8881 20297
rect 7171 20269 7961 20293
rect 8013 20269 8039 20293
rect 8091 20269 8881 20293
rect 7171 20245 7640 20269
rect 4964 20233 7640 20245
rect 4964 20181 5201 20233
rect 5253 20181 5279 20233
rect 5331 20181 6121 20233
rect 6173 20181 6199 20233
rect 6251 20181 7041 20233
rect 7093 20181 7119 20233
rect 7171 20213 7640 20233
rect 7696 20213 7726 20269
rect 7782 20213 7812 20269
rect 7868 20213 7898 20269
rect 7954 20245 7961 20269
rect 7954 20233 7984 20245
rect 8040 20233 8070 20245
rect 7954 20213 7961 20233
rect 8126 20213 8156 20269
rect 8212 20213 8242 20269
rect 8298 20213 8327 20269
rect 8383 20213 8412 20269
rect 8468 20213 8497 20269
rect 8553 20245 8881 20269
rect 8933 20245 8959 20297
rect 9011 20293 9079 20297
rect 9135 20293 9170 20349
rect 9226 20293 9260 20349
rect 9316 20293 9350 20349
rect 9406 20293 9440 20349
rect 9496 20293 9530 20349
rect 9586 20293 9620 20349
rect 9676 20293 9710 20349
rect 9766 20309 9801 20349
rect 9853 20309 9879 20361
rect 9931 20309 10721 20361
rect 10773 20309 10799 20361
rect 10851 20309 11641 20361
rect 11693 20309 11719 20361
rect 11771 20309 12561 20361
rect 12613 20309 12639 20361
rect 12691 20309 14858 20361
rect 9766 20297 14858 20309
rect 9766 20293 9801 20297
rect 9011 20269 9801 20293
rect 9011 20245 9079 20269
rect 8553 20233 9079 20245
rect 8553 20213 8881 20233
rect 7171 20189 7961 20213
rect 8013 20189 8039 20213
rect 8091 20189 8881 20213
rect 7171 20181 7640 20189
rect 4964 20169 7640 20181
rect 4964 20117 5201 20169
rect 5253 20117 5279 20169
rect 5331 20117 6121 20169
rect 6173 20117 6199 20169
rect 6251 20117 7041 20169
rect 7093 20117 7119 20169
rect 7171 20133 7640 20169
rect 7696 20133 7726 20189
rect 7782 20133 7812 20189
rect 7868 20133 7898 20189
rect 7954 20181 7961 20189
rect 7954 20169 7984 20181
rect 8040 20169 8070 20181
rect 7954 20133 7961 20169
rect 8126 20133 8156 20189
rect 8212 20133 8242 20189
rect 8298 20133 8327 20189
rect 8383 20133 8412 20189
rect 8468 20133 8497 20189
rect 8553 20181 8881 20189
rect 8933 20181 8959 20233
rect 9011 20213 9079 20233
rect 9135 20213 9170 20269
rect 9226 20213 9260 20269
rect 9316 20213 9350 20269
rect 9406 20213 9440 20269
rect 9496 20213 9530 20269
rect 9586 20213 9620 20269
rect 9676 20213 9710 20269
rect 9766 20245 9801 20269
rect 9853 20245 9879 20297
rect 9931 20245 10721 20297
rect 10773 20245 10799 20297
rect 10851 20245 11641 20297
rect 11693 20245 11719 20297
rect 11771 20245 12561 20297
rect 12613 20245 12639 20297
rect 12691 20245 14858 20297
rect 9766 20233 14858 20245
rect 9766 20213 9801 20233
rect 9011 20189 9801 20213
rect 9011 20181 9079 20189
rect 8553 20169 9079 20181
rect 8553 20133 8881 20169
rect 7171 20117 7961 20133
rect 8013 20117 8039 20133
rect 8091 20117 8881 20133
rect 8933 20117 8959 20169
rect 9011 20133 9079 20169
rect 9135 20133 9170 20189
rect 9226 20133 9260 20189
rect 9316 20133 9350 20189
rect 9406 20133 9440 20189
rect 9496 20133 9530 20189
rect 9586 20133 9620 20189
rect 9676 20133 9710 20189
rect 9766 20181 9801 20189
rect 9853 20181 9879 20233
rect 9931 20181 10721 20233
rect 10773 20181 10799 20233
rect 10851 20181 11641 20233
rect 11693 20181 11719 20233
rect 11771 20181 12561 20233
rect 12613 20181 12639 20233
rect 12691 20181 14858 20233
rect 9766 20169 14858 20181
rect 9766 20133 9801 20169
rect 9011 20117 9801 20133
rect 9853 20117 9879 20169
rect 9931 20117 10721 20169
rect 10773 20117 10799 20169
rect 10851 20117 11641 20169
rect 11693 20117 11719 20169
rect 11771 20117 12561 20169
rect 12613 20117 12639 20169
rect 12691 20117 14858 20169
rect 4964 20109 14858 20117
rect 4964 20105 7640 20109
rect 4964 20053 5201 20105
rect 5253 20053 5279 20105
rect 5331 20053 6121 20105
rect 6173 20053 6199 20105
rect 6251 20053 7041 20105
rect 7093 20053 7119 20105
rect 7171 20053 7640 20105
rect 7696 20053 7726 20109
rect 7782 20053 7812 20109
rect 7868 20053 7898 20109
rect 7954 20105 7984 20109
rect 8040 20105 8070 20109
rect 7954 20053 7961 20105
rect 8126 20053 8156 20109
rect 8212 20053 8242 20109
rect 8298 20053 8327 20109
rect 8383 20053 8412 20109
rect 8468 20053 8497 20109
rect 8553 20105 9079 20109
rect 8553 20053 8881 20105
rect 8933 20053 8959 20105
rect 9011 20053 9079 20105
rect 9135 20053 9170 20109
rect 9226 20053 9260 20109
rect 9316 20053 9350 20109
rect 9406 20053 9440 20109
rect 9496 20053 9530 20109
rect 9586 20053 9620 20109
rect 9676 20053 9710 20109
rect 9766 20105 14858 20109
rect 9766 20053 9801 20105
rect 9853 20053 9879 20105
rect 9931 20053 10721 20105
rect 10773 20053 10799 20105
rect 10851 20053 11641 20105
rect 11693 20053 11719 20105
rect 11771 20053 12561 20105
rect 12613 20053 12639 20105
rect 12691 20053 14858 20105
rect 4964 20041 14858 20053
rect 4964 19989 5201 20041
rect 5253 19989 5279 20041
rect 5331 19989 6121 20041
rect 6173 19989 6199 20041
rect 6251 19989 7041 20041
rect 7093 19989 7119 20041
rect 7171 20029 7961 20041
rect 8013 20029 8039 20041
rect 8091 20029 8881 20041
rect 7171 19989 7640 20029
rect 4964 19977 7640 19989
rect 4964 19925 5201 19977
rect 5253 19925 5279 19977
rect 5331 19925 6121 19977
rect 6173 19925 6199 19977
rect 6251 19925 7041 19977
rect 7093 19925 7119 19977
rect 7171 19973 7640 19977
rect 7696 19973 7726 20029
rect 7782 19973 7812 20029
rect 7868 19973 7898 20029
rect 7954 19989 7961 20029
rect 7954 19977 7984 19989
rect 8040 19977 8070 19989
rect 7954 19973 7961 19977
rect 8126 19973 8156 20029
rect 8212 19973 8242 20029
rect 8298 19973 8327 20029
rect 8383 19973 8412 20029
rect 8468 19973 8497 20029
rect 8553 19989 8881 20029
rect 8933 19989 8959 20041
rect 9011 20029 9801 20041
rect 9011 19989 9079 20029
rect 8553 19977 9079 19989
rect 8553 19973 8881 19977
rect 7171 19949 7961 19973
rect 8013 19949 8039 19973
rect 8091 19949 8881 19973
rect 7171 19925 7640 19949
rect 4964 19913 7640 19925
rect 4964 19861 5201 19913
rect 5253 19861 5279 19913
rect 5331 19861 6121 19913
rect 6173 19861 6199 19913
rect 6251 19861 7041 19913
rect 7093 19861 7119 19913
rect 7171 19893 7640 19913
rect 7696 19893 7726 19949
rect 7782 19893 7812 19949
rect 7868 19893 7898 19949
rect 7954 19925 7961 19949
rect 7954 19913 7984 19925
rect 8040 19913 8070 19925
rect 7954 19893 7961 19913
rect 8126 19893 8156 19949
rect 8212 19893 8242 19949
rect 8298 19893 8327 19949
rect 8383 19893 8412 19949
rect 8468 19893 8497 19949
rect 8553 19925 8881 19949
rect 8933 19925 8959 19977
rect 9011 19973 9079 19977
rect 9135 19973 9170 20029
rect 9226 19973 9260 20029
rect 9316 19973 9350 20029
rect 9406 19973 9440 20029
rect 9496 19973 9530 20029
rect 9586 19973 9620 20029
rect 9676 19973 9710 20029
rect 9766 19989 9801 20029
rect 9853 19989 9879 20041
rect 9931 19989 10721 20041
rect 10773 19989 10799 20041
rect 10851 19989 11641 20041
rect 11693 19989 11719 20041
rect 11771 19989 12561 20041
rect 12613 19989 12639 20041
rect 12691 19989 14858 20041
rect 9766 19977 14858 19989
rect 9766 19973 9801 19977
rect 9011 19949 9801 19973
rect 9011 19925 9079 19949
rect 8553 19913 9079 19925
rect 8553 19893 8881 19913
rect 7171 19869 7961 19893
rect 8013 19869 8039 19893
rect 8091 19869 8881 19893
rect 7171 19861 7640 19869
rect 4964 19849 7640 19861
rect 4964 19797 5201 19849
rect 5253 19797 5279 19849
rect 5331 19797 6121 19849
rect 6173 19797 6199 19849
rect 6251 19797 7041 19849
rect 7093 19797 7119 19849
rect 7171 19813 7640 19849
rect 7696 19813 7726 19869
rect 7782 19813 7812 19869
rect 7868 19813 7898 19869
rect 7954 19861 7961 19869
rect 7954 19849 7984 19861
rect 8040 19849 8070 19861
rect 7954 19813 7961 19849
rect 8126 19813 8156 19869
rect 8212 19813 8242 19869
rect 8298 19813 8327 19869
rect 8383 19813 8412 19869
rect 8468 19813 8497 19869
rect 8553 19861 8881 19869
rect 8933 19861 8959 19913
rect 9011 19893 9079 19913
rect 9135 19893 9170 19949
rect 9226 19893 9260 19949
rect 9316 19893 9350 19949
rect 9406 19893 9440 19949
rect 9496 19893 9530 19949
rect 9586 19893 9620 19949
rect 9676 19893 9710 19949
rect 9766 19925 9801 19949
rect 9853 19925 9879 19977
rect 9931 19925 10721 19977
rect 10773 19925 10799 19977
rect 10851 19925 11641 19977
rect 11693 19925 11719 19977
rect 11771 19925 12561 19977
rect 12613 19925 12639 19977
rect 12691 19925 14858 19977
rect 9766 19913 14858 19925
rect 9766 19893 9801 19913
rect 9011 19869 9801 19893
rect 9011 19861 9079 19869
rect 8553 19849 9079 19861
rect 8553 19813 8881 19849
rect 7171 19797 7961 19813
rect 8013 19797 8039 19813
rect 8091 19797 8881 19813
rect 8933 19797 8959 19849
rect 9011 19813 9079 19849
rect 9135 19813 9170 19869
rect 9226 19813 9260 19869
rect 9316 19813 9350 19869
rect 9406 19813 9440 19869
rect 9496 19813 9530 19869
rect 9586 19813 9620 19869
rect 9676 19813 9710 19869
rect 9766 19861 9801 19869
rect 9853 19861 9879 19913
rect 9931 19861 10721 19913
rect 10773 19861 10799 19913
rect 10851 19861 11641 19913
rect 11693 19861 11719 19913
rect 11771 19861 12561 19913
rect 12613 19861 12639 19913
rect 12691 19861 14858 19913
rect 9766 19849 14858 19861
rect 9766 19813 9801 19849
rect 9011 19797 9801 19813
rect 9853 19797 9879 19849
rect 9931 19797 10721 19849
rect 10773 19797 10799 19849
rect 10851 19797 11641 19849
rect 11693 19797 11719 19849
rect 11771 19797 12561 19849
rect 12613 19797 12639 19849
rect 12691 19797 14858 19849
rect 4964 19789 14858 19797
rect 4964 19785 7640 19789
rect 4964 19733 5201 19785
rect 5253 19733 5279 19785
rect 5331 19733 6121 19785
rect 6173 19733 6199 19785
rect 6251 19733 7041 19785
rect 7093 19733 7119 19785
rect 7171 19733 7640 19785
rect 7696 19733 7726 19789
rect 7782 19733 7812 19789
rect 7868 19733 7898 19789
rect 7954 19785 7984 19789
rect 8040 19785 8070 19789
rect 7954 19733 7961 19785
rect 8126 19733 8156 19789
rect 8212 19733 8242 19789
rect 8298 19733 8327 19789
rect 8383 19733 8412 19789
rect 8468 19733 8497 19789
rect 8553 19785 9079 19789
rect 8553 19733 8881 19785
rect 8933 19733 8959 19785
rect 9011 19733 9079 19785
rect 9135 19733 9170 19789
rect 9226 19733 9260 19789
rect 9316 19733 9350 19789
rect 9406 19733 9440 19789
rect 9496 19733 9530 19789
rect 9586 19733 9620 19789
rect 9676 19733 9710 19789
rect 9766 19785 14858 19789
rect 9766 19733 9801 19785
rect 9853 19733 9879 19785
rect 9931 19733 10721 19785
rect 10773 19733 10799 19785
rect 10851 19733 11641 19785
rect 11693 19733 11719 19785
rect 11771 19733 12561 19785
rect 12613 19733 12639 19785
rect 12691 19733 14858 19785
rect 4964 19721 14858 19733
rect 4964 19669 5201 19721
rect 5253 19669 5279 19721
rect 5331 19669 6121 19721
rect 6173 19669 6199 19721
rect 6251 19669 7041 19721
rect 7093 19669 7119 19721
rect 7171 19709 7961 19721
rect 8013 19709 8039 19721
rect 8091 19709 8881 19721
rect 7171 19669 7640 19709
rect 4964 19657 7640 19669
rect 4964 19605 5201 19657
rect 5253 19605 5279 19657
rect 5331 19605 6121 19657
rect 6173 19605 6199 19657
rect 6251 19605 7041 19657
rect 7093 19605 7119 19657
rect 7171 19653 7640 19657
rect 7696 19653 7726 19709
rect 7782 19653 7812 19709
rect 7868 19653 7898 19709
rect 7954 19669 7961 19709
rect 7954 19657 7984 19669
rect 8040 19657 8070 19669
rect 7954 19653 7961 19657
rect 8126 19653 8156 19709
rect 8212 19653 8242 19709
rect 8298 19653 8327 19709
rect 8383 19653 8412 19709
rect 8468 19653 8497 19709
rect 8553 19669 8881 19709
rect 8933 19669 8959 19721
rect 9011 19709 9801 19721
rect 9011 19669 9079 19709
rect 8553 19657 9079 19669
rect 8553 19653 8881 19657
rect 7171 19629 7961 19653
rect 8013 19629 8039 19653
rect 8091 19629 8881 19653
rect 7171 19605 7640 19629
rect 4964 19593 7640 19605
rect 4964 19541 5201 19593
rect 5253 19541 5279 19593
rect 5331 19541 6121 19593
rect 6173 19541 6199 19593
rect 6251 19541 7041 19593
rect 7093 19541 7119 19593
rect 7171 19573 7640 19593
rect 7696 19573 7726 19629
rect 7782 19573 7812 19629
rect 7868 19573 7898 19629
rect 7954 19605 7961 19629
rect 7954 19593 7984 19605
rect 8040 19593 8070 19605
rect 7954 19573 7961 19593
rect 8126 19573 8156 19629
rect 8212 19573 8242 19629
rect 8298 19573 8327 19629
rect 8383 19573 8412 19629
rect 8468 19573 8497 19629
rect 8553 19605 8881 19629
rect 8933 19605 8959 19657
rect 9011 19653 9079 19657
rect 9135 19653 9170 19709
rect 9226 19653 9260 19709
rect 9316 19653 9350 19709
rect 9406 19653 9440 19709
rect 9496 19653 9530 19709
rect 9586 19653 9620 19709
rect 9676 19653 9710 19709
rect 9766 19669 9801 19709
rect 9853 19669 9879 19721
rect 9931 19669 10721 19721
rect 10773 19669 10799 19721
rect 10851 19669 11641 19721
rect 11693 19669 11719 19721
rect 11771 19669 12561 19721
rect 12613 19669 12639 19721
rect 12691 19669 14858 19721
rect 9766 19657 14858 19669
rect 9766 19653 9801 19657
rect 9011 19629 9801 19653
rect 9011 19605 9079 19629
rect 8553 19593 9079 19605
rect 8553 19573 8881 19593
rect 7171 19549 7961 19573
rect 8013 19549 8039 19573
rect 8091 19549 8881 19573
rect 7171 19541 7640 19549
rect 4964 19529 7640 19541
rect 4964 19477 5201 19529
rect 5253 19477 5279 19529
rect 5331 19477 6121 19529
rect 6173 19477 6199 19529
rect 6251 19477 7041 19529
rect 7093 19477 7119 19529
rect 7171 19493 7640 19529
rect 7696 19493 7726 19549
rect 7782 19493 7812 19549
rect 7868 19493 7898 19549
rect 7954 19541 7961 19549
rect 7954 19529 7984 19541
rect 8040 19529 8070 19541
rect 7954 19493 7961 19529
rect 8126 19493 8156 19549
rect 8212 19493 8242 19549
rect 8298 19493 8327 19549
rect 8383 19493 8412 19549
rect 8468 19493 8497 19549
rect 8553 19541 8881 19549
rect 8933 19541 8959 19593
rect 9011 19573 9079 19593
rect 9135 19573 9170 19629
rect 9226 19573 9260 19629
rect 9316 19573 9350 19629
rect 9406 19573 9440 19629
rect 9496 19573 9530 19629
rect 9586 19573 9620 19629
rect 9676 19573 9710 19629
rect 9766 19605 9801 19629
rect 9853 19605 9879 19657
rect 9931 19605 10721 19657
rect 10773 19605 10799 19657
rect 10851 19605 11641 19657
rect 11693 19605 11719 19657
rect 11771 19605 12561 19657
rect 12613 19605 12639 19657
rect 12691 19605 14858 19657
rect 9766 19593 14858 19605
rect 9766 19573 9801 19593
rect 9011 19549 9801 19573
rect 9011 19541 9079 19549
rect 8553 19529 9079 19541
rect 8553 19493 8881 19529
rect 7171 19477 7961 19493
rect 8013 19477 8039 19493
rect 8091 19477 8881 19493
rect 8933 19477 8959 19529
rect 9011 19493 9079 19529
rect 9135 19493 9170 19549
rect 9226 19493 9260 19549
rect 9316 19493 9350 19549
rect 9406 19493 9440 19549
rect 9496 19493 9530 19549
rect 9586 19493 9620 19549
rect 9676 19493 9710 19549
rect 9766 19541 9801 19549
rect 9853 19541 9879 19593
rect 9931 19541 10721 19593
rect 10773 19541 10799 19593
rect 10851 19541 11641 19593
rect 11693 19541 11719 19593
rect 11771 19541 12561 19593
rect 12613 19541 12639 19593
rect 12691 19541 14858 19593
rect 9766 19529 14858 19541
rect 9766 19493 9801 19529
rect 9011 19477 9801 19493
rect 9853 19477 9879 19529
rect 9931 19477 10721 19529
rect 10773 19477 10799 19529
rect 10851 19477 11641 19529
rect 11693 19477 11719 19529
rect 11771 19477 12561 19529
rect 12613 19477 12639 19529
rect 12691 19477 14858 19529
rect 4964 19469 14858 19477
rect 4964 19464 7640 19469
rect 4964 19412 5201 19464
rect 5253 19412 5279 19464
rect 5331 19412 6121 19464
rect 6173 19412 6199 19464
rect 6251 19412 7041 19464
rect 7093 19412 7119 19464
rect 7171 19413 7640 19464
rect 7696 19413 7726 19469
rect 7782 19413 7812 19469
rect 7868 19413 7898 19469
rect 7954 19464 7984 19469
rect 8040 19464 8070 19469
rect 7954 19413 7961 19464
rect 8126 19413 8156 19469
rect 8212 19413 8242 19469
rect 8298 19413 8327 19469
rect 8383 19413 8412 19469
rect 8468 19413 8497 19469
rect 8553 19464 9079 19469
rect 8553 19413 8881 19464
rect 7171 19412 7961 19413
rect 8013 19412 8039 19413
rect 8091 19412 8881 19413
rect 8933 19412 8959 19464
rect 9011 19413 9079 19464
rect 9135 19413 9170 19469
rect 9226 19413 9260 19469
rect 9316 19413 9350 19469
rect 9406 19413 9440 19469
rect 9496 19413 9530 19469
rect 9586 19413 9620 19469
rect 9676 19413 9710 19469
rect 9766 19464 14858 19469
rect 9766 19413 9801 19464
rect 9011 19412 9801 19413
rect 9853 19412 9879 19464
rect 9931 19412 10721 19464
rect 10773 19412 10799 19464
rect 10851 19412 11641 19464
rect 11693 19412 11719 19464
rect 11771 19412 12561 19464
rect 12613 19412 12639 19464
rect 12691 19412 14858 19464
rect 4964 19399 14858 19412
rect 4964 19347 5201 19399
rect 5253 19347 5279 19399
rect 5331 19347 6121 19399
rect 6173 19347 6199 19399
rect 6251 19347 7041 19399
rect 7093 19347 7119 19399
rect 7171 19389 7961 19399
rect 8013 19389 8039 19399
rect 8091 19389 8881 19399
rect 7171 19347 7640 19389
rect 4964 19334 7640 19347
rect 4964 19282 5201 19334
rect 5253 19282 5279 19334
rect 5331 19282 6121 19334
rect 6173 19282 6199 19334
rect 6251 19282 7041 19334
rect 7093 19282 7119 19334
rect 7171 19333 7640 19334
rect 7696 19333 7726 19389
rect 7782 19333 7812 19389
rect 7868 19333 7898 19389
rect 7954 19347 7961 19389
rect 7954 19334 7984 19347
rect 8040 19334 8070 19347
rect 7954 19333 7961 19334
rect 8126 19333 8156 19389
rect 8212 19333 8242 19389
rect 8298 19333 8327 19389
rect 8383 19333 8412 19389
rect 8468 19333 8497 19389
rect 8553 19347 8881 19389
rect 8933 19347 8959 19399
rect 9011 19389 9801 19399
rect 9011 19347 9079 19389
rect 8553 19334 9079 19347
rect 8553 19333 8881 19334
rect 7171 19309 7961 19333
rect 8013 19309 8039 19333
rect 8091 19309 8881 19333
rect 7171 19282 7640 19309
rect 4964 19269 7640 19282
rect 4964 19217 5201 19269
rect 5253 19217 5279 19269
rect 5331 19217 6121 19269
rect 6173 19217 6199 19269
rect 6251 19217 7041 19269
rect 7093 19217 7119 19269
rect 7171 19253 7640 19269
rect 7696 19253 7726 19309
rect 7782 19253 7812 19309
rect 7868 19253 7898 19309
rect 7954 19282 7961 19309
rect 7954 19269 7984 19282
rect 8040 19269 8070 19282
rect 7954 19253 7961 19269
rect 8126 19253 8156 19309
rect 8212 19253 8242 19309
rect 8298 19253 8327 19309
rect 8383 19253 8412 19309
rect 8468 19253 8497 19309
rect 8553 19282 8881 19309
rect 8933 19282 8959 19334
rect 9011 19333 9079 19334
rect 9135 19333 9170 19389
rect 9226 19333 9260 19389
rect 9316 19333 9350 19389
rect 9406 19333 9440 19389
rect 9496 19333 9530 19389
rect 9586 19333 9620 19389
rect 9676 19333 9710 19389
rect 9766 19347 9801 19389
rect 9853 19347 9879 19399
rect 9931 19347 10721 19399
rect 10773 19347 10799 19399
rect 10851 19347 11641 19399
rect 11693 19347 11719 19399
rect 11771 19347 12561 19399
rect 12613 19347 12639 19399
rect 12691 19347 14858 19399
rect 9766 19334 14858 19347
rect 9766 19333 9801 19334
rect 9011 19309 9801 19333
rect 9011 19282 9079 19309
rect 8553 19269 9079 19282
rect 8553 19253 8881 19269
rect 7171 19229 7961 19253
rect 8013 19229 8039 19253
rect 8091 19229 8881 19253
rect 7171 19217 7640 19229
rect 4964 19204 7640 19217
rect 4964 19152 5201 19204
rect 5253 19152 5279 19204
rect 5331 19152 6121 19204
rect 6173 19152 6199 19204
rect 6251 19152 7041 19204
rect 7093 19152 7119 19204
rect 7171 19173 7640 19204
rect 7696 19173 7726 19229
rect 7782 19173 7812 19229
rect 7868 19173 7898 19229
rect 7954 19217 7961 19229
rect 7954 19204 7984 19217
rect 8040 19204 8070 19217
rect 7954 19173 7961 19204
rect 8126 19173 8156 19229
rect 8212 19173 8242 19229
rect 8298 19173 8327 19229
rect 8383 19173 8412 19229
rect 8468 19173 8497 19229
rect 8553 19217 8881 19229
rect 8933 19217 8959 19269
rect 9011 19253 9079 19269
rect 9135 19253 9170 19309
rect 9226 19253 9260 19309
rect 9316 19253 9350 19309
rect 9406 19253 9440 19309
rect 9496 19253 9530 19309
rect 9586 19253 9620 19309
rect 9676 19253 9710 19309
rect 9766 19282 9801 19309
rect 9853 19282 9879 19334
rect 9931 19282 10721 19334
rect 10773 19282 10799 19334
rect 10851 19282 11641 19334
rect 11693 19282 11719 19334
rect 11771 19282 12561 19334
rect 12613 19282 12639 19334
rect 12691 19282 14858 19334
rect 9766 19269 14858 19282
rect 9766 19253 9801 19269
rect 9011 19229 9801 19253
rect 9011 19217 9079 19229
rect 8553 19204 9079 19217
rect 8553 19173 8881 19204
rect 7171 19152 7961 19173
rect 8013 19152 8039 19173
rect 8091 19152 8881 19173
rect 8933 19152 8959 19204
rect 9011 19173 9079 19204
rect 9135 19173 9170 19229
rect 9226 19173 9260 19229
rect 9316 19173 9350 19229
rect 9406 19173 9440 19229
rect 9496 19173 9530 19229
rect 9586 19173 9620 19229
rect 9676 19173 9710 19229
rect 9766 19217 9801 19229
rect 9853 19217 9879 19269
rect 9931 19217 10721 19269
rect 10773 19217 10799 19269
rect 10851 19217 11641 19269
rect 11693 19217 11719 19269
rect 11771 19217 12561 19269
rect 12613 19217 12639 19269
rect 12691 19217 14858 19269
rect 9766 19204 14858 19217
rect 9766 19173 9801 19204
rect 9011 19152 9801 19173
rect 9853 19152 9879 19204
rect 9931 19152 10721 19204
rect 10773 19152 10799 19204
rect 10851 19152 11641 19204
rect 11693 19152 11719 19204
rect 11771 19152 12561 19204
rect 12613 19152 12639 19204
rect 12691 19152 14858 19204
rect 4964 19149 14858 19152
rect 4964 19139 7640 19149
rect 4964 19087 5201 19139
rect 5253 19087 5279 19139
rect 5331 19087 6121 19139
rect 6173 19087 6199 19139
rect 6251 19087 7041 19139
rect 7093 19087 7119 19139
rect 7171 19093 7640 19139
rect 7696 19093 7726 19149
rect 7782 19093 7812 19149
rect 7868 19093 7898 19149
rect 7954 19139 7984 19149
rect 8040 19139 8070 19149
rect 7954 19093 7961 19139
rect 8126 19093 8156 19149
rect 8212 19093 8242 19149
rect 8298 19093 8327 19149
rect 8383 19093 8412 19149
rect 8468 19093 8497 19149
rect 8553 19139 9079 19149
rect 8553 19093 8881 19139
rect 7171 19087 7961 19093
rect 8013 19087 8039 19093
rect 8091 19087 8881 19093
rect 8933 19087 8959 19139
rect 9011 19093 9079 19139
rect 9135 19093 9170 19149
rect 9226 19093 9260 19149
rect 9316 19093 9350 19149
rect 9406 19093 9440 19149
rect 9496 19093 9530 19149
rect 9586 19093 9620 19149
rect 9676 19093 9710 19149
rect 9766 19139 14858 19149
rect 9766 19093 9801 19139
rect 9011 19087 9801 19093
rect 9853 19087 9879 19139
rect 9931 19087 10721 19139
rect 10773 19087 10799 19139
rect 10851 19087 11641 19139
rect 11693 19087 11719 19139
rect 11771 19087 12561 19139
rect 12613 19087 12639 19139
rect 12691 19087 14858 19139
rect 4964 19074 14858 19087
rect 4964 19022 5201 19074
rect 5253 19022 5279 19074
rect 5331 19022 6121 19074
rect 6173 19022 6199 19074
rect 6251 19022 7041 19074
rect 7093 19022 7119 19074
rect 7171 19069 7961 19074
rect 8013 19069 8039 19074
rect 8091 19069 8881 19074
rect 7171 19022 7640 19069
rect 4964 19013 7640 19022
rect 7696 19013 7726 19069
rect 7782 19013 7812 19069
rect 7868 19013 7898 19069
rect 7954 19022 7961 19069
rect 7954 19013 7984 19022
rect 8040 19013 8070 19022
rect 8126 19013 8156 19069
rect 8212 19013 8242 19069
rect 8298 19013 8327 19069
rect 8383 19013 8412 19069
rect 8468 19013 8497 19069
rect 8553 19022 8881 19069
rect 8933 19022 8959 19074
rect 9011 19069 9801 19074
rect 9011 19022 9079 19069
rect 8553 19013 9079 19022
rect 9135 19013 9170 19069
rect 9226 19013 9260 19069
rect 9316 19013 9350 19069
rect 9406 19013 9440 19069
rect 9496 19013 9530 19069
rect 9586 19013 9620 19069
rect 9676 19013 9710 19069
rect 9766 19022 9801 19069
rect 9853 19022 9879 19074
rect 9931 19022 10721 19074
rect 10773 19022 10799 19074
rect 10851 19022 11641 19074
rect 11693 19022 11719 19074
rect 11771 19022 12561 19074
rect 12613 19022 12639 19074
rect 12691 19022 14858 19074
rect 9766 19013 14858 19022
rect 4964 19009 14858 19013
rect 4964 18957 5201 19009
rect 5253 18957 5279 19009
rect 5331 18957 6121 19009
rect 6173 18957 6199 19009
rect 6251 18957 7041 19009
rect 7093 18957 7119 19009
rect 7171 18989 7961 19009
rect 8013 18989 8039 19009
rect 8091 18989 8881 19009
rect 7171 18957 7640 18989
rect 4964 18944 7640 18957
rect 4964 18892 5201 18944
rect 5253 18892 5279 18944
rect 5331 18892 6121 18944
rect 6173 18892 6199 18944
rect 6251 18892 7041 18944
rect 7093 18892 7119 18944
rect 7171 18933 7640 18944
rect 7696 18933 7726 18989
rect 7782 18933 7812 18989
rect 7868 18933 7898 18989
rect 7954 18957 7961 18989
rect 7954 18944 7984 18957
rect 8040 18944 8070 18957
rect 7954 18933 7961 18944
rect 8126 18933 8156 18989
rect 8212 18933 8242 18989
rect 8298 18933 8327 18989
rect 8383 18933 8412 18989
rect 8468 18933 8497 18989
rect 8553 18957 8881 18989
rect 8933 18957 8959 19009
rect 9011 18989 9801 19009
rect 9011 18957 9079 18989
rect 8553 18944 9079 18957
rect 8553 18933 8881 18944
rect 7171 18909 7961 18933
rect 8013 18909 8039 18933
rect 8091 18909 8881 18933
rect 7171 18892 7640 18909
rect 4964 18879 7640 18892
rect 4964 18827 5201 18879
rect 5253 18827 5279 18879
rect 5331 18827 6121 18879
rect 6173 18827 6199 18879
rect 6251 18827 7041 18879
rect 7093 18827 7119 18879
rect 7171 18853 7640 18879
rect 7696 18853 7726 18909
rect 7782 18853 7812 18909
rect 7868 18853 7898 18909
rect 7954 18892 7961 18909
rect 7954 18879 7984 18892
rect 8040 18879 8070 18892
rect 7954 18853 7961 18879
rect 8126 18853 8156 18909
rect 8212 18853 8242 18909
rect 8298 18853 8327 18909
rect 8383 18853 8412 18909
rect 8468 18853 8497 18909
rect 8553 18892 8881 18909
rect 8933 18892 8959 18944
rect 9011 18933 9079 18944
rect 9135 18933 9170 18989
rect 9226 18933 9260 18989
rect 9316 18933 9350 18989
rect 9406 18933 9440 18989
rect 9496 18933 9530 18989
rect 9586 18933 9620 18989
rect 9676 18933 9710 18989
rect 9766 18957 9801 18989
rect 9853 18957 9879 19009
rect 9931 18957 10721 19009
rect 10773 18957 10799 19009
rect 10851 18957 11641 19009
rect 11693 18957 11719 19009
rect 11771 18957 12561 19009
rect 12613 18957 12639 19009
rect 12691 18957 14858 19009
rect 9766 18944 14858 18957
rect 9766 18933 9801 18944
rect 9011 18909 9801 18933
rect 9011 18892 9079 18909
rect 8553 18879 9079 18892
rect 8553 18853 8881 18879
rect 7171 18829 7961 18853
rect 8013 18829 8039 18853
rect 8091 18829 8881 18853
rect 7171 18827 7640 18829
rect 4964 18814 7640 18827
rect 4964 18762 5201 18814
rect 5253 18762 5279 18814
rect 5331 18762 6121 18814
rect 6173 18762 6199 18814
rect 6251 18762 7041 18814
rect 7093 18762 7119 18814
rect 7171 18773 7640 18814
rect 7696 18773 7726 18829
rect 7782 18773 7812 18829
rect 7868 18773 7898 18829
rect 7954 18827 7961 18829
rect 7954 18814 7984 18827
rect 8040 18814 8070 18827
rect 7954 18773 7961 18814
rect 8126 18773 8156 18829
rect 8212 18773 8242 18829
rect 8298 18773 8327 18829
rect 8383 18773 8412 18829
rect 8468 18773 8497 18829
rect 8553 18827 8881 18829
rect 8933 18827 8959 18879
rect 9011 18853 9079 18879
rect 9135 18853 9170 18909
rect 9226 18853 9260 18909
rect 9316 18853 9350 18909
rect 9406 18853 9440 18909
rect 9496 18853 9530 18909
rect 9586 18853 9620 18909
rect 9676 18853 9710 18909
rect 9766 18892 9801 18909
rect 9853 18892 9879 18944
rect 9931 18892 10721 18944
rect 10773 18892 10799 18944
rect 10851 18892 11641 18944
rect 11693 18892 11719 18944
rect 11771 18892 12561 18944
rect 12613 18892 12639 18944
rect 12691 18892 14858 18944
rect 9766 18879 14858 18892
rect 9766 18853 9801 18879
rect 9011 18829 9801 18853
rect 9011 18827 9079 18829
rect 8553 18814 9079 18827
rect 8553 18773 8881 18814
rect 7171 18762 7961 18773
rect 8013 18762 8039 18773
rect 8091 18762 8881 18773
rect 8933 18762 8959 18814
rect 9011 18773 9079 18814
rect 9135 18773 9170 18829
rect 9226 18773 9260 18829
rect 9316 18773 9350 18829
rect 9406 18773 9440 18829
rect 9496 18773 9530 18829
rect 9586 18773 9620 18829
rect 9676 18773 9710 18829
rect 9766 18827 9801 18829
rect 9853 18827 9879 18879
rect 9931 18827 10721 18879
rect 10773 18827 10799 18879
rect 10851 18827 11641 18879
rect 11693 18827 11719 18879
rect 11771 18827 12561 18879
rect 12613 18827 12639 18879
rect 12691 18827 14858 18879
rect 9766 18814 14858 18827
rect 9766 18773 9801 18814
rect 9011 18762 9801 18773
rect 9853 18762 9879 18814
rect 9931 18762 10721 18814
rect 10773 18762 10799 18814
rect 10851 18762 11641 18814
rect 11693 18762 11719 18814
rect 11771 18762 12561 18814
rect 12613 18762 12639 18814
rect 12691 18762 14858 18814
rect 4964 18749 14858 18762
rect 4964 18697 5201 18749
rect 5253 18697 5279 18749
rect 5331 18697 6121 18749
rect 6173 18697 6199 18749
rect 6251 18697 7041 18749
rect 7093 18697 7119 18749
rect 7171 18697 7640 18749
rect 4964 18693 7640 18697
rect 7696 18693 7726 18749
rect 7782 18693 7812 18749
rect 7868 18693 7898 18749
rect 7954 18697 7961 18749
rect 7954 18693 7984 18697
rect 8040 18693 8070 18697
rect 8126 18693 8156 18749
rect 8212 18693 8242 18749
rect 8298 18693 8327 18749
rect 8383 18693 8412 18749
rect 8468 18693 8497 18749
rect 8553 18697 8881 18749
rect 8933 18697 8959 18749
rect 9011 18697 9079 18749
rect 8553 18693 9079 18697
rect 9135 18693 9170 18749
rect 9226 18693 9260 18749
rect 9316 18693 9350 18749
rect 9406 18693 9440 18749
rect 9496 18693 9530 18749
rect 9586 18693 9620 18749
rect 9676 18693 9710 18749
rect 9766 18697 9801 18749
rect 9853 18697 9879 18749
rect 9931 18697 10721 18749
rect 10773 18697 10799 18749
rect 10851 18697 11641 18749
rect 11693 18697 11719 18749
rect 11771 18697 12561 18749
rect 12613 18697 12639 18749
rect 12691 18697 14858 18749
rect 9766 18693 14858 18697
rect 4964 18691 14858 18693
tri 2824 17896 3533 18605 sw
tri 11513 17982 12222 18691 ne
rect 187 17894 11341 17896
rect 187 17890 5188 17894
rect 187 17838 4712 17890
rect 4764 17838 4780 17890
rect 4832 17838 4848 17890
rect 4900 17838 5188 17890
rect 5244 17838 5270 17894
rect 5326 17838 5352 17894
rect 5408 17838 5434 17894
rect 5490 17838 5516 17894
rect 5572 17838 5598 17894
rect 5654 17890 5680 17894
rect 5736 17890 5762 17894
rect 5818 17890 5844 17894
rect 5752 17838 5762 17890
rect 5820 17838 5844 17890
rect 5900 17838 5926 17894
rect 5982 17838 6008 17894
rect 6064 17838 6090 17894
rect 6146 17838 6172 17894
rect 6228 17838 6254 17894
rect 6310 17838 6336 17894
rect 6392 17838 6418 17894
rect 6474 17838 6500 17894
rect 6556 17890 6582 17894
rect 6638 17890 6664 17894
rect 6720 17890 6746 17894
rect 6740 17838 6746 17890
rect 6802 17838 6828 17894
rect 6884 17838 6909 17894
rect 6965 17838 6990 17894
rect 7046 17838 7071 17894
rect 7127 17838 7152 17894
rect 7208 17838 7233 17894
rect 7289 17838 7314 17894
rect 7370 17890 11341 17894
rect 7370 17838 7472 17890
rect 7524 17838 7540 17890
rect 7592 17838 7608 17890
rect 7660 17838 8392 17890
rect 8444 17838 8460 17890
rect 8512 17838 8528 17890
rect 8580 17838 9312 17890
rect 9364 17838 9380 17890
rect 9432 17838 9448 17890
rect 9500 17838 10232 17890
rect 10284 17838 10300 17890
rect 10352 17838 10368 17890
rect 10420 17838 11152 17890
rect 11204 17838 11220 17890
rect 11272 17838 11288 17890
rect 11340 17838 11341 17890
rect 187 17826 11341 17838
rect 187 17774 4712 17826
rect 4764 17774 4780 17826
rect 4832 17774 4848 17826
rect 4900 17814 5632 17826
rect 5684 17814 5700 17826
rect 5752 17814 5768 17826
rect 5820 17814 6552 17826
rect 6604 17814 6620 17826
rect 6672 17814 6688 17826
rect 6740 17814 7472 17826
rect 4900 17774 5188 17814
rect 187 17762 5188 17774
rect 187 17710 4712 17762
rect 4764 17710 4780 17762
rect 4832 17710 4848 17762
rect 4900 17758 5188 17762
rect 5244 17758 5270 17814
rect 5326 17758 5352 17814
rect 5408 17758 5434 17814
rect 5490 17758 5516 17814
rect 5572 17758 5598 17814
rect 5752 17774 5762 17814
rect 5820 17774 5844 17814
rect 5654 17762 5680 17774
rect 5736 17762 5762 17774
rect 5818 17762 5844 17774
rect 5752 17758 5762 17762
rect 5820 17758 5844 17762
rect 5900 17758 5926 17814
rect 5982 17758 6008 17814
rect 6064 17758 6090 17814
rect 6146 17758 6172 17814
rect 6228 17758 6254 17814
rect 6310 17758 6336 17814
rect 6392 17758 6418 17814
rect 6474 17758 6500 17814
rect 6740 17774 6746 17814
rect 6556 17762 6582 17774
rect 6638 17762 6664 17774
rect 6720 17762 6746 17774
rect 6740 17758 6746 17762
rect 6802 17758 6828 17814
rect 6884 17758 6909 17814
rect 6965 17758 6990 17814
rect 7046 17758 7071 17814
rect 7127 17758 7152 17814
rect 7208 17758 7233 17814
rect 7289 17758 7314 17814
rect 7370 17774 7472 17814
rect 7524 17774 7540 17826
rect 7592 17774 7608 17826
rect 7660 17774 8392 17826
rect 8444 17774 8460 17826
rect 8512 17774 8528 17826
rect 8580 17774 9312 17826
rect 9364 17774 9380 17826
rect 9432 17774 9448 17826
rect 9500 17774 10232 17826
rect 10284 17774 10300 17826
rect 10352 17774 10368 17826
rect 10420 17774 11152 17826
rect 11204 17774 11220 17826
rect 11272 17774 11288 17826
rect 11340 17774 11341 17826
rect 7370 17762 11341 17774
rect 7370 17758 7472 17762
rect 4900 17734 5632 17758
rect 5684 17734 5700 17758
rect 5752 17734 5768 17758
rect 5820 17734 6552 17758
rect 6604 17734 6620 17758
rect 6672 17734 6688 17758
rect 6740 17734 7472 17758
rect 4900 17710 5188 17734
rect 187 17698 5188 17710
rect 187 17646 4712 17698
rect 4764 17646 4780 17698
rect 4832 17646 4848 17698
rect 4900 17678 5188 17698
rect 5244 17678 5270 17734
rect 5326 17678 5352 17734
rect 5408 17678 5434 17734
rect 5490 17678 5516 17734
rect 5572 17678 5598 17734
rect 5752 17710 5762 17734
rect 5820 17710 5844 17734
rect 5654 17698 5680 17710
rect 5736 17698 5762 17710
rect 5818 17698 5844 17710
rect 5752 17678 5762 17698
rect 5820 17678 5844 17698
rect 5900 17678 5926 17734
rect 5982 17678 6008 17734
rect 6064 17678 6090 17734
rect 6146 17678 6172 17734
rect 6228 17678 6254 17734
rect 6310 17678 6336 17734
rect 6392 17678 6418 17734
rect 6474 17678 6500 17734
rect 6740 17710 6746 17734
rect 6556 17698 6582 17710
rect 6638 17698 6664 17710
rect 6720 17698 6746 17710
rect 6740 17678 6746 17698
rect 6802 17678 6828 17734
rect 6884 17678 6909 17734
rect 6965 17678 6990 17734
rect 7046 17678 7071 17734
rect 7127 17678 7152 17734
rect 7208 17678 7233 17734
rect 7289 17678 7314 17734
rect 7370 17710 7472 17734
rect 7524 17710 7540 17762
rect 7592 17710 7608 17762
rect 7660 17710 8392 17762
rect 8444 17710 8460 17762
rect 8512 17710 8528 17762
rect 8580 17710 9312 17762
rect 9364 17710 9380 17762
rect 9432 17710 9448 17762
rect 9500 17710 10232 17762
rect 10284 17710 10300 17762
rect 10352 17710 10368 17762
rect 10420 17710 11152 17762
rect 11204 17710 11220 17762
rect 11272 17710 11288 17762
rect 11340 17710 11341 17762
rect 7370 17698 11341 17710
rect 7370 17678 7472 17698
rect 4900 17654 5632 17678
rect 5684 17654 5700 17678
rect 5752 17654 5768 17678
rect 5820 17654 6552 17678
rect 6604 17654 6620 17678
rect 6672 17654 6688 17678
rect 6740 17654 7472 17678
rect 4900 17646 5188 17654
rect 187 17634 5188 17646
rect 187 17582 4712 17634
rect 4764 17582 4780 17634
rect 4832 17582 4848 17634
rect 4900 17598 5188 17634
rect 5244 17598 5270 17654
rect 5326 17598 5352 17654
rect 5408 17598 5434 17654
rect 5490 17598 5516 17654
rect 5572 17598 5598 17654
rect 5752 17646 5762 17654
rect 5820 17646 5844 17654
rect 5654 17634 5680 17646
rect 5736 17634 5762 17646
rect 5818 17634 5844 17646
rect 5752 17598 5762 17634
rect 5820 17598 5844 17634
rect 5900 17598 5926 17654
rect 5982 17598 6008 17654
rect 6064 17598 6090 17654
rect 6146 17598 6172 17654
rect 6228 17598 6254 17654
rect 6310 17598 6336 17654
rect 6392 17598 6418 17654
rect 6474 17598 6500 17654
rect 6740 17646 6746 17654
rect 6556 17634 6582 17646
rect 6638 17634 6664 17646
rect 6720 17634 6746 17646
rect 6740 17598 6746 17634
rect 6802 17598 6828 17654
rect 6884 17598 6909 17654
rect 6965 17598 6990 17654
rect 7046 17598 7071 17654
rect 7127 17598 7152 17654
rect 7208 17598 7233 17654
rect 7289 17598 7314 17654
rect 7370 17646 7472 17654
rect 7524 17646 7540 17698
rect 7592 17646 7608 17698
rect 7660 17646 8392 17698
rect 8444 17646 8460 17698
rect 8512 17646 8528 17698
rect 8580 17646 9312 17698
rect 9364 17646 9380 17698
rect 9432 17646 9448 17698
rect 9500 17646 10232 17698
rect 10284 17646 10300 17698
rect 10352 17646 10368 17698
rect 10420 17646 11152 17698
rect 11204 17646 11220 17698
rect 11272 17646 11288 17698
rect 11340 17646 11341 17698
rect 7370 17634 11341 17646
rect 7370 17598 7472 17634
rect 4900 17582 5632 17598
rect 5684 17582 5700 17598
rect 5752 17582 5768 17598
rect 5820 17582 6552 17598
rect 6604 17582 6620 17598
rect 6672 17582 6688 17598
rect 6740 17582 7472 17598
rect 7524 17582 7540 17634
rect 7592 17582 7608 17634
rect 7660 17582 8392 17634
rect 8444 17582 8460 17634
rect 8512 17582 8528 17634
rect 8580 17582 9312 17634
rect 9364 17582 9380 17634
rect 9432 17582 9448 17634
rect 9500 17582 10232 17634
rect 10284 17582 10300 17634
rect 10352 17582 10368 17634
rect 10420 17582 11152 17634
rect 11204 17582 11220 17634
rect 11272 17582 11288 17634
rect 11340 17582 11341 17634
rect 187 17574 11341 17582
rect 187 17570 5188 17574
rect 187 17518 4712 17570
rect 4764 17518 4780 17570
rect 4832 17518 4848 17570
rect 4900 17518 5188 17570
rect 5244 17518 5270 17574
rect 5326 17518 5352 17574
rect 5408 17518 5434 17574
rect 5490 17518 5516 17574
rect 5572 17518 5598 17574
rect 5654 17570 5680 17574
rect 5736 17570 5762 17574
rect 5818 17570 5844 17574
rect 5752 17518 5762 17570
rect 5820 17518 5844 17570
rect 5900 17518 5926 17574
rect 5982 17518 6008 17574
rect 6064 17518 6090 17574
rect 6146 17518 6172 17574
rect 6228 17518 6254 17574
rect 6310 17518 6336 17574
rect 6392 17518 6418 17574
rect 6474 17518 6500 17574
rect 6556 17570 6582 17574
rect 6638 17570 6664 17574
rect 6720 17570 6746 17574
rect 6740 17518 6746 17570
rect 6802 17518 6828 17574
rect 6884 17518 6909 17574
rect 6965 17518 6990 17574
rect 7046 17518 7071 17574
rect 7127 17518 7152 17574
rect 7208 17518 7233 17574
rect 7289 17518 7314 17574
rect 7370 17570 11341 17574
rect 7370 17518 7472 17570
rect 7524 17518 7540 17570
rect 7592 17518 7608 17570
rect 7660 17518 8392 17570
rect 8444 17518 8460 17570
rect 8512 17518 8528 17570
rect 8580 17518 9312 17570
rect 9364 17518 9380 17570
rect 9432 17518 9448 17570
rect 9500 17518 10232 17570
rect 10284 17518 10300 17570
rect 10352 17518 10368 17570
rect 10420 17518 11152 17570
rect 11204 17518 11220 17570
rect 11272 17518 11288 17570
rect 11340 17518 11341 17570
rect 187 17506 11341 17518
rect 187 17454 4712 17506
rect 4764 17454 4780 17506
rect 4832 17454 4848 17506
rect 4900 17494 5632 17506
rect 5684 17494 5700 17506
rect 5752 17494 5768 17506
rect 5820 17494 6552 17506
rect 6604 17494 6620 17506
rect 6672 17494 6688 17506
rect 6740 17494 7472 17506
rect 4900 17454 5188 17494
rect 187 17442 5188 17454
rect 187 17390 4712 17442
rect 4764 17390 4780 17442
rect 4832 17390 4848 17442
rect 4900 17438 5188 17442
rect 5244 17438 5270 17494
rect 5326 17438 5352 17494
rect 5408 17438 5434 17494
rect 5490 17438 5516 17494
rect 5572 17438 5598 17494
rect 5752 17454 5762 17494
rect 5820 17454 5844 17494
rect 5654 17442 5680 17454
rect 5736 17442 5762 17454
rect 5818 17442 5844 17454
rect 5752 17438 5762 17442
rect 5820 17438 5844 17442
rect 5900 17438 5926 17494
rect 5982 17438 6008 17494
rect 6064 17438 6090 17494
rect 6146 17438 6172 17494
rect 6228 17438 6254 17494
rect 6310 17438 6336 17494
rect 6392 17438 6418 17494
rect 6474 17438 6500 17494
rect 6740 17454 6746 17494
rect 6556 17442 6582 17454
rect 6638 17442 6664 17454
rect 6720 17442 6746 17454
rect 6740 17438 6746 17442
rect 6802 17438 6828 17494
rect 6884 17438 6909 17494
rect 6965 17438 6990 17494
rect 7046 17438 7071 17494
rect 7127 17438 7152 17494
rect 7208 17438 7233 17494
rect 7289 17438 7314 17494
rect 7370 17454 7472 17494
rect 7524 17454 7540 17506
rect 7592 17454 7608 17506
rect 7660 17454 8392 17506
rect 8444 17454 8460 17506
rect 8512 17454 8528 17506
rect 8580 17454 9312 17506
rect 9364 17454 9380 17506
rect 9432 17454 9448 17506
rect 9500 17454 10232 17506
rect 10284 17454 10300 17506
rect 10352 17454 10368 17506
rect 10420 17454 11152 17506
rect 11204 17454 11220 17506
rect 11272 17454 11288 17506
rect 11340 17454 11341 17506
rect 7370 17442 11341 17454
rect 7370 17438 7472 17442
rect 4900 17414 5632 17438
rect 5684 17414 5700 17438
rect 5752 17414 5768 17438
rect 5820 17414 6552 17438
rect 6604 17414 6620 17438
rect 6672 17414 6688 17438
rect 6740 17414 7472 17438
rect 4900 17390 5188 17414
rect 187 17378 5188 17390
rect 187 17326 4712 17378
rect 4764 17326 4780 17378
rect 4832 17326 4848 17378
rect 4900 17358 5188 17378
rect 5244 17358 5270 17414
rect 5326 17358 5352 17414
rect 5408 17358 5434 17414
rect 5490 17358 5516 17414
rect 5572 17358 5598 17414
rect 5752 17390 5762 17414
rect 5820 17390 5844 17414
rect 5654 17378 5680 17390
rect 5736 17378 5762 17390
rect 5818 17378 5844 17390
rect 5752 17358 5762 17378
rect 5820 17358 5844 17378
rect 5900 17358 5926 17414
rect 5982 17358 6008 17414
rect 6064 17358 6090 17414
rect 6146 17358 6172 17414
rect 6228 17358 6254 17414
rect 6310 17358 6336 17414
rect 6392 17358 6418 17414
rect 6474 17358 6500 17414
rect 6740 17390 6746 17414
rect 6556 17378 6582 17390
rect 6638 17378 6664 17390
rect 6720 17378 6746 17390
rect 6740 17358 6746 17378
rect 6802 17358 6828 17414
rect 6884 17358 6909 17414
rect 6965 17358 6990 17414
rect 7046 17358 7071 17414
rect 7127 17358 7152 17414
rect 7208 17358 7233 17414
rect 7289 17358 7314 17414
rect 7370 17390 7472 17414
rect 7524 17390 7540 17442
rect 7592 17390 7608 17442
rect 7660 17390 8392 17442
rect 8444 17390 8460 17442
rect 8512 17390 8528 17442
rect 8580 17390 9312 17442
rect 9364 17390 9380 17442
rect 9432 17390 9448 17442
rect 9500 17390 10232 17442
rect 10284 17390 10300 17442
rect 10352 17390 10368 17442
rect 10420 17390 11152 17442
rect 11204 17390 11220 17442
rect 11272 17390 11288 17442
rect 11340 17390 11341 17442
rect 7370 17378 11341 17390
rect 7370 17358 7472 17378
rect 4900 17334 5632 17358
rect 5684 17334 5700 17358
rect 5752 17334 5768 17358
rect 5820 17334 6552 17358
rect 6604 17334 6620 17358
rect 6672 17334 6688 17358
rect 6740 17334 7472 17358
rect 4900 17326 5188 17334
rect 187 17314 5188 17326
rect 187 17262 4712 17314
rect 4764 17262 4780 17314
rect 4832 17262 4848 17314
rect 4900 17278 5188 17314
rect 5244 17278 5270 17334
rect 5326 17278 5352 17334
rect 5408 17278 5434 17334
rect 5490 17278 5516 17334
rect 5572 17278 5598 17334
rect 5752 17326 5762 17334
rect 5820 17326 5844 17334
rect 5654 17314 5680 17326
rect 5736 17314 5762 17326
rect 5818 17314 5844 17326
rect 5752 17278 5762 17314
rect 5820 17278 5844 17314
rect 5900 17278 5926 17334
rect 5982 17278 6008 17334
rect 6064 17278 6090 17334
rect 6146 17278 6172 17334
rect 6228 17278 6254 17334
rect 6310 17278 6336 17334
rect 6392 17278 6418 17334
rect 6474 17278 6500 17334
rect 6740 17326 6746 17334
rect 6556 17314 6582 17326
rect 6638 17314 6664 17326
rect 6720 17314 6746 17326
rect 6740 17278 6746 17314
rect 6802 17278 6828 17334
rect 6884 17278 6909 17334
rect 6965 17278 6990 17334
rect 7046 17278 7071 17334
rect 7127 17278 7152 17334
rect 7208 17278 7233 17334
rect 7289 17278 7314 17334
rect 7370 17326 7472 17334
rect 7524 17326 7540 17378
rect 7592 17326 7608 17378
rect 7660 17326 8392 17378
rect 8444 17326 8460 17378
rect 8512 17326 8528 17378
rect 8580 17326 9312 17378
rect 9364 17326 9380 17378
rect 9432 17326 9448 17378
rect 9500 17326 10232 17378
rect 10284 17326 10300 17378
rect 10352 17326 10368 17378
rect 10420 17326 11152 17378
rect 11204 17326 11220 17378
rect 11272 17326 11288 17378
rect 11340 17326 11341 17378
rect 7370 17314 11341 17326
rect 7370 17278 7472 17314
rect 4900 17262 5632 17278
rect 5684 17262 5700 17278
rect 5752 17262 5768 17278
rect 5820 17262 6552 17278
rect 6604 17262 6620 17278
rect 6672 17262 6688 17278
rect 6740 17262 7472 17278
rect 7524 17262 7540 17314
rect 7592 17262 7608 17314
rect 7660 17262 8392 17314
rect 8444 17262 8460 17314
rect 8512 17262 8528 17314
rect 8580 17262 9312 17314
rect 9364 17262 9380 17314
rect 9432 17262 9448 17314
rect 9500 17262 10232 17314
rect 10284 17262 10300 17314
rect 10352 17262 10368 17314
rect 10420 17262 11152 17314
rect 11204 17262 11220 17314
rect 11272 17262 11288 17314
rect 11340 17262 11341 17314
rect 187 17254 11341 17262
rect 187 17250 5188 17254
rect 187 17198 4712 17250
rect 4764 17198 4780 17250
rect 4832 17198 4848 17250
rect 4900 17198 5188 17250
rect 5244 17198 5270 17254
rect 5326 17198 5352 17254
rect 5408 17198 5434 17254
rect 5490 17198 5516 17254
rect 5572 17198 5598 17254
rect 5654 17250 5680 17254
rect 5736 17250 5762 17254
rect 5818 17250 5844 17254
rect 5752 17198 5762 17250
rect 5820 17198 5844 17250
rect 5900 17198 5926 17254
rect 5982 17198 6008 17254
rect 6064 17198 6090 17254
rect 6146 17198 6172 17254
rect 6228 17198 6254 17254
rect 6310 17198 6336 17254
rect 6392 17198 6418 17254
rect 6474 17198 6500 17254
rect 6556 17250 6582 17254
rect 6638 17250 6664 17254
rect 6720 17250 6746 17254
rect 6740 17198 6746 17250
rect 6802 17198 6828 17254
rect 6884 17198 6909 17254
rect 6965 17198 6990 17254
rect 7046 17198 7071 17254
rect 7127 17198 7152 17254
rect 7208 17198 7233 17254
rect 7289 17198 7314 17254
rect 7370 17250 11341 17254
rect 7370 17198 7472 17250
rect 7524 17198 7540 17250
rect 7592 17198 7608 17250
rect 7660 17198 8392 17250
rect 8444 17198 8460 17250
rect 8512 17198 8528 17250
rect 8580 17198 9312 17250
rect 9364 17198 9380 17250
rect 9432 17198 9448 17250
rect 9500 17198 10232 17250
rect 10284 17198 10300 17250
rect 10352 17198 10368 17250
rect 10420 17198 11152 17250
rect 11204 17198 11220 17250
rect 11272 17198 11288 17250
rect 11340 17198 11341 17250
rect 187 17186 11341 17198
rect 187 17134 4712 17186
rect 4764 17134 4780 17186
rect 4832 17134 4848 17186
rect 4900 17174 5632 17186
rect 5684 17174 5700 17186
rect 5752 17174 5768 17186
rect 5820 17174 6552 17186
rect 6604 17174 6620 17186
rect 6672 17174 6688 17186
rect 6740 17174 7472 17186
rect 4900 17134 5188 17174
rect 187 17122 5188 17134
rect 187 17070 4712 17122
rect 4764 17070 4780 17122
rect 4832 17070 4848 17122
rect 4900 17118 5188 17122
rect 5244 17118 5270 17174
rect 5326 17118 5352 17174
rect 5408 17118 5434 17174
rect 5490 17118 5516 17174
rect 5572 17118 5598 17174
rect 5752 17134 5762 17174
rect 5820 17134 5844 17174
rect 5654 17122 5680 17134
rect 5736 17122 5762 17134
rect 5818 17122 5844 17134
rect 5752 17118 5762 17122
rect 5820 17118 5844 17122
rect 5900 17118 5926 17174
rect 5982 17118 6008 17174
rect 6064 17118 6090 17174
rect 6146 17118 6172 17174
rect 6228 17118 6254 17174
rect 6310 17118 6336 17174
rect 6392 17118 6418 17174
rect 6474 17118 6500 17174
rect 6740 17134 6746 17174
rect 6556 17122 6582 17134
rect 6638 17122 6664 17134
rect 6720 17122 6746 17134
rect 6740 17118 6746 17122
rect 6802 17118 6828 17174
rect 6884 17118 6909 17174
rect 6965 17118 6990 17174
rect 7046 17118 7071 17174
rect 7127 17118 7152 17174
rect 7208 17118 7233 17174
rect 7289 17118 7314 17174
rect 7370 17134 7472 17174
rect 7524 17134 7540 17186
rect 7592 17134 7608 17186
rect 7660 17134 8392 17186
rect 8444 17134 8460 17186
rect 8512 17134 8528 17186
rect 8580 17134 9312 17186
rect 9364 17134 9380 17186
rect 9432 17134 9448 17186
rect 9500 17134 10232 17186
rect 10284 17134 10300 17186
rect 10352 17134 10368 17186
rect 10420 17134 11152 17186
rect 11204 17134 11220 17186
rect 11272 17134 11288 17186
rect 11340 17134 11341 17186
rect 7370 17122 11341 17134
rect 7370 17118 7472 17122
rect 4900 17094 5632 17118
rect 5684 17094 5700 17118
rect 5752 17094 5768 17118
rect 5820 17094 6552 17118
rect 6604 17094 6620 17118
rect 6672 17094 6688 17118
rect 6740 17094 7472 17118
rect 4900 17070 5188 17094
rect 187 17058 5188 17070
rect 187 17006 4712 17058
rect 4764 17006 4780 17058
rect 4832 17006 4848 17058
rect 4900 17038 5188 17058
rect 5244 17038 5270 17094
rect 5326 17038 5352 17094
rect 5408 17038 5434 17094
rect 5490 17038 5516 17094
rect 5572 17038 5598 17094
rect 5752 17070 5762 17094
rect 5820 17070 5844 17094
rect 5654 17058 5680 17070
rect 5736 17058 5762 17070
rect 5818 17058 5844 17070
rect 5752 17038 5762 17058
rect 5820 17038 5844 17058
rect 5900 17038 5926 17094
rect 5982 17038 6008 17094
rect 6064 17038 6090 17094
rect 6146 17038 6172 17094
rect 6228 17038 6254 17094
rect 6310 17038 6336 17094
rect 6392 17038 6418 17094
rect 6474 17038 6500 17094
rect 6740 17070 6746 17094
rect 6556 17058 6582 17070
rect 6638 17058 6664 17070
rect 6720 17058 6746 17070
rect 6740 17038 6746 17058
rect 6802 17038 6828 17094
rect 6884 17038 6909 17094
rect 6965 17038 6990 17094
rect 7046 17038 7071 17094
rect 7127 17038 7152 17094
rect 7208 17038 7233 17094
rect 7289 17038 7314 17094
rect 7370 17070 7472 17094
rect 7524 17070 7540 17122
rect 7592 17070 7608 17122
rect 7660 17070 8392 17122
rect 8444 17070 8460 17122
rect 8512 17070 8528 17122
rect 8580 17070 9312 17122
rect 9364 17070 9380 17122
rect 9432 17070 9448 17122
rect 9500 17070 10232 17122
rect 10284 17070 10300 17122
rect 10352 17070 10368 17122
rect 10420 17070 11152 17122
rect 11204 17070 11220 17122
rect 11272 17070 11288 17122
rect 11340 17070 11341 17122
rect 7370 17058 11341 17070
rect 7370 17038 7472 17058
rect 4900 17014 5632 17038
rect 5684 17014 5700 17038
rect 5752 17014 5768 17038
rect 5820 17014 6552 17038
rect 6604 17014 6620 17038
rect 6672 17014 6688 17038
rect 6740 17014 7472 17038
rect 4900 17006 5188 17014
rect 187 16994 5188 17006
rect 187 16942 4712 16994
rect 4764 16942 4780 16994
rect 4832 16942 4848 16994
rect 4900 16958 5188 16994
rect 5244 16958 5270 17014
rect 5326 16958 5352 17014
rect 5408 16958 5434 17014
rect 5490 16958 5516 17014
rect 5572 16958 5598 17014
rect 5752 17006 5762 17014
rect 5820 17006 5844 17014
rect 5654 16994 5680 17006
rect 5736 16994 5762 17006
rect 5818 16994 5844 17006
rect 5752 16958 5762 16994
rect 5820 16958 5844 16994
rect 5900 16958 5926 17014
rect 5982 16958 6008 17014
rect 6064 16958 6090 17014
rect 6146 16958 6172 17014
rect 6228 16958 6254 17014
rect 6310 16958 6336 17014
rect 6392 16958 6418 17014
rect 6474 16958 6500 17014
rect 6740 17006 6746 17014
rect 6556 16994 6582 17006
rect 6638 16994 6664 17006
rect 6720 16994 6746 17006
rect 6740 16958 6746 16994
rect 6802 16958 6828 17014
rect 6884 16958 6909 17014
rect 6965 16958 6990 17014
rect 7046 16958 7071 17014
rect 7127 16958 7152 17014
rect 7208 16958 7233 17014
rect 7289 16958 7314 17014
rect 7370 17006 7472 17014
rect 7524 17006 7540 17058
rect 7592 17006 7608 17058
rect 7660 17006 8392 17058
rect 8444 17006 8460 17058
rect 8512 17006 8528 17058
rect 8580 17006 9312 17058
rect 9364 17006 9380 17058
rect 9432 17006 9448 17058
rect 9500 17006 10232 17058
rect 10284 17006 10300 17058
rect 10352 17006 10368 17058
rect 10420 17006 11152 17058
rect 11204 17006 11220 17058
rect 11272 17006 11288 17058
rect 11340 17006 11341 17058
rect 7370 16994 11341 17006
rect 7370 16958 7472 16994
rect 4900 16942 5632 16958
rect 5684 16942 5700 16958
rect 5752 16942 5768 16958
rect 5820 16942 6552 16958
rect 6604 16942 6620 16958
rect 6672 16942 6688 16958
rect 6740 16942 7472 16958
rect 7524 16942 7540 16994
rect 7592 16942 7608 16994
rect 7660 16942 8392 16994
rect 8444 16942 8460 16994
rect 8512 16942 8528 16994
rect 8580 16942 9312 16994
rect 9364 16942 9380 16994
rect 9432 16942 9448 16994
rect 9500 16942 10232 16994
rect 10284 16942 10300 16994
rect 10352 16942 10368 16994
rect 10420 16942 11152 16994
rect 11204 16942 11220 16994
rect 11272 16942 11288 16994
rect 11340 16942 11341 16994
rect 187 16934 11341 16942
rect 187 16929 5188 16934
rect 187 16877 4712 16929
rect 4764 16877 4780 16929
rect 4832 16877 4848 16929
rect 4900 16878 5188 16929
rect 5244 16878 5270 16934
rect 5326 16878 5352 16934
rect 5408 16878 5434 16934
rect 5490 16878 5516 16934
rect 5572 16878 5598 16934
rect 5654 16929 5680 16934
rect 5736 16929 5762 16934
rect 5818 16929 5844 16934
rect 5752 16878 5762 16929
rect 5820 16878 5844 16929
rect 5900 16878 5926 16934
rect 5982 16878 6008 16934
rect 6064 16878 6090 16934
rect 6146 16878 6172 16934
rect 6228 16878 6254 16934
rect 6310 16878 6336 16934
rect 6392 16878 6418 16934
rect 6474 16878 6500 16934
rect 6556 16929 6582 16934
rect 6638 16929 6664 16934
rect 6720 16929 6746 16934
rect 6740 16878 6746 16929
rect 6802 16878 6828 16934
rect 6884 16878 6909 16934
rect 6965 16878 6990 16934
rect 7046 16878 7071 16934
rect 7127 16878 7152 16934
rect 7208 16878 7233 16934
rect 7289 16878 7314 16934
rect 7370 16929 11341 16934
rect 7370 16878 7472 16929
rect 4900 16877 5632 16878
rect 5684 16877 5700 16878
rect 5752 16877 5768 16878
rect 5820 16877 6552 16878
rect 6604 16877 6620 16878
rect 6672 16877 6688 16878
rect 6740 16877 7472 16878
rect 7524 16877 7540 16929
rect 7592 16877 7608 16929
rect 7660 16877 8392 16929
rect 8444 16877 8460 16929
rect 8512 16877 8528 16929
rect 8580 16877 9312 16929
rect 9364 16877 9380 16929
rect 9432 16877 9448 16929
rect 9500 16877 10232 16929
rect 10284 16877 10300 16929
rect 10352 16877 10368 16929
rect 10420 16877 11152 16929
rect 11204 16877 11220 16929
rect 11272 16877 11288 16929
rect 11340 16877 11341 16929
rect 187 16864 11341 16877
rect 187 16812 4712 16864
rect 4764 16812 4780 16864
rect 4832 16812 4848 16864
rect 4900 16854 5632 16864
rect 5684 16854 5700 16864
rect 5752 16854 5768 16864
rect 5820 16854 6552 16864
rect 6604 16854 6620 16864
rect 6672 16854 6688 16864
rect 6740 16854 7472 16864
rect 4900 16812 5188 16854
rect 187 16799 5188 16812
rect 187 16747 4712 16799
rect 4764 16747 4780 16799
rect 4832 16747 4848 16799
rect 4900 16798 5188 16799
rect 5244 16798 5270 16854
rect 5326 16798 5352 16854
rect 5408 16798 5434 16854
rect 5490 16798 5516 16854
rect 5572 16798 5598 16854
rect 5752 16812 5762 16854
rect 5820 16812 5844 16854
rect 5654 16799 5680 16812
rect 5736 16799 5762 16812
rect 5818 16799 5844 16812
rect 5752 16798 5762 16799
rect 5820 16798 5844 16799
rect 5900 16798 5926 16854
rect 5982 16798 6008 16854
rect 6064 16798 6090 16854
rect 6146 16798 6172 16854
rect 6228 16798 6254 16854
rect 6310 16798 6336 16854
rect 6392 16798 6418 16854
rect 6474 16798 6500 16854
rect 6740 16812 6746 16854
rect 6556 16799 6582 16812
rect 6638 16799 6664 16812
rect 6720 16799 6746 16812
rect 6740 16798 6746 16799
rect 6802 16798 6828 16854
rect 6884 16798 6909 16854
rect 6965 16798 6990 16854
rect 7046 16798 7071 16854
rect 7127 16798 7152 16854
rect 7208 16798 7233 16854
rect 7289 16798 7314 16854
rect 7370 16812 7472 16854
rect 7524 16812 7540 16864
rect 7592 16812 7608 16864
rect 7660 16812 8392 16864
rect 8444 16812 8460 16864
rect 8512 16812 8528 16864
rect 8580 16812 9312 16864
rect 9364 16812 9380 16864
rect 9432 16812 9448 16864
rect 9500 16812 10232 16864
rect 10284 16812 10300 16864
rect 10352 16812 10368 16864
rect 10420 16812 11152 16864
rect 11204 16812 11220 16864
rect 11272 16812 11288 16864
rect 11340 16812 11341 16864
rect 7370 16799 11341 16812
rect 7370 16798 7472 16799
rect 4900 16774 5632 16798
rect 5684 16774 5700 16798
rect 5752 16774 5768 16798
rect 5820 16774 6552 16798
rect 6604 16774 6620 16798
rect 6672 16774 6688 16798
rect 6740 16774 7472 16798
rect 4900 16747 5188 16774
rect 187 16734 5188 16747
rect 187 16682 4712 16734
rect 4764 16682 4780 16734
rect 4832 16682 4848 16734
rect 4900 16718 5188 16734
rect 5244 16718 5270 16774
rect 5326 16718 5352 16774
rect 5408 16718 5434 16774
rect 5490 16718 5516 16774
rect 5572 16718 5598 16774
rect 5752 16747 5762 16774
rect 5820 16747 5844 16774
rect 5654 16734 5680 16747
rect 5736 16734 5762 16747
rect 5818 16734 5844 16747
rect 5752 16718 5762 16734
rect 5820 16718 5844 16734
rect 5900 16718 5926 16774
rect 5982 16718 6008 16774
rect 6064 16718 6090 16774
rect 6146 16718 6172 16774
rect 6228 16718 6254 16774
rect 6310 16718 6336 16774
rect 6392 16718 6418 16774
rect 6474 16718 6500 16774
rect 6740 16747 6746 16774
rect 6556 16734 6582 16747
rect 6638 16734 6664 16747
rect 6720 16734 6746 16747
rect 6740 16718 6746 16734
rect 6802 16718 6828 16774
rect 6884 16718 6909 16774
rect 6965 16718 6990 16774
rect 7046 16718 7071 16774
rect 7127 16718 7152 16774
rect 7208 16718 7233 16774
rect 7289 16718 7314 16774
rect 7370 16747 7472 16774
rect 7524 16747 7540 16799
rect 7592 16747 7608 16799
rect 7660 16747 8392 16799
rect 8444 16747 8460 16799
rect 8512 16747 8528 16799
rect 8580 16747 9312 16799
rect 9364 16747 9380 16799
rect 9432 16747 9448 16799
rect 9500 16747 10232 16799
rect 10284 16747 10300 16799
rect 10352 16747 10368 16799
rect 10420 16747 11152 16799
rect 11204 16747 11220 16799
rect 11272 16747 11288 16799
rect 11340 16747 11341 16799
rect 7370 16734 11341 16747
rect 7370 16718 7472 16734
rect 4900 16694 5632 16718
rect 5684 16694 5700 16718
rect 5752 16694 5768 16718
rect 5820 16694 6552 16718
rect 6604 16694 6620 16718
rect 6672 16694 6688 16718
rect 6740 16694 7472 16718
rect 4900 16682 5188 16694
rect 187 16669 5188 16682
rect 187 16617 4712 16669
rect 4764 16617 4780 16669
rect 4832 16617 4848 16669
rect 4900 16638 5188 16669
rect 5244 16638 5270 16694
rect 5326 16638 5352 16694
rect 5408 16638 5434 16694
rect 5490 16638 5516 16694
rect 5572 16638 5598 16694
rect 5752 16682 5762 16694
rect 5820 16682 5844 16694
rect 5654 16669 5680 16682
rect 5736 16669 5762 16682
rect 5818 16669 5844 16682
rect 5752 16638 5762 16669
rect 5820 16638 5844 16669
rect 5900 16638 5926 16694
rect 5982 16638 6008 16694
rect 6064 16638 6090 16694
rect 6146 16638 6172 16694
rect 6228 16638 6254 16694
rect 6310 16638 6336 16694
rect 6392 16638 6418 16694
rect 6474 16638 6500 16694
rect 6740 16682 6746 16694
rect 6556 16669 6582 16682
rect 6638 16669 6664 16682
rect 6720 16669 6746 16682
rect 6740 16638 6746 16669
rect 6802 16638 6828 16694
rect 6884 16638 6909 16694
rect 6965 16638 6990 16694
rect 7046 16638 7071 16694
rect 7127 16638 7152 16694
rect 7208 16638 7233 16694
rect 7289 16638 7314 16694
rect 7370 16682 7472 16694
rect 7524 16682 7540 16734
rect 7592 16682 7608 16734
rect 7660 16682 8392 16734
rect 8444 16682 8460 16734
rect 8512 16682 8528 16734
rect 8580 16682 9312 16734
rect 9364 16682 9380 16734
rect 9432 16682 9448 16734
rect 9500 16682 10232 16734
rect 10284 16682 10300 16734
rect 10352 16682 10368 16734
rect 10420 16682 11152 16734
rect 11204 16682 11220 16734
rect 11272 16682 11288 16734
rect 11340 16682 11341 16734
rect 7370 16669 11341 16682
rect 7370 16638 7472 16669
rect 4900 16617 5632 16638
rect 5684 16617 5700 16638
rect 5752 16617 5768 16638
rect 5820 16617 6552 16638
rect 6604 16617 6620 16638
rect 6672 16617 6688 16638
rect 6740 16617 7472 16638
rect 7524 16617 7540 16669
rect 7592 16617 7608 16669
rect 7660 16617 8392 16669
rect 8444 16617 8460 16669
rect 8512 16617 8528 16669
rect 8580 16617 9312 16669
rect 9364 16617 9380 16669
rect 9432 16617 9448 16669
rect 9500 16617 10232 16669
rect 10284 16617 10300 16669
rect 10352 16617 10368 16669
rect 10420 16617 11152 16669
rect 11204 16617 11220 16669
rect 11272 16617 11288 16669
rect 11340 16617 11341 16669
rect 187 16614 11341 16617
rect 187 16604 5188 16614
rect 187 16552 4712 16604
rect 4764 16552 4780 16604
rect 4832 16552 4848 16604
rect 4900 16558 5188 16604
rect 5244 16558 5270 16614
rect 5326 16558 5352 16614
rect 5408 16558 5434 16614
rect 5490 16558 5516 16614
rect 5572 16558 5598 16614
rect 5654 16604 5680 16614
rect 5736 16604 5762 16614
rect 5818 16604 5844 16614
rect 5752 16558 5762 16604
rect 5820 16558 5844 16604
rect 5900 16558 5926 16614
rect 5982 16558 6008 16614
rect 6064 16558 6090 16614
rect 6146 16558 6172 16614
rect 6228 16558 6254 16614
rect 6310 16558 6336 16614
rect 6392 16558 6418 16614
rect 6474 16558 6500 16614
rect 6556 16604 6582 16614
rect 6638 16604 6664 16614
rect 6720 16604 6746 16614
rect 6740 16558 6746 16604
rect 6802 16558 6828 16614
rect 6884 16558 6909 16614
rect 6965 16558 6990 16614
rect 7046 16558 7071 16614
rect 7127 16558 7152 16614
rect 7208 16558 7233 16614
rect 7289 16558 7314 16614
rect 7370 16604 11341 16614
rect 7370 16558 7472 16604
rect 4900 16552 5632 16558
rect 5684 16552 5700 16558
rect 5752 16552 5768 16558
rect 5820 16552 6552 16558
rect 6604 16552 6620 16558
rect 6672 16552 6688 16558
rect 6740 16552 7472 16558
rect 7524 16552 7540 16604
rect 7592 16552 7608 16604
rect 7660 16552 8392 16604
rect 8444 16552 8460 16604
rect 8512 16552 8528 16604
rect 8580 16552 9312 16604
rect 9364 16552 9380 16604
rect 9432 16552 9448 16604
rect 9500 16552 10232 16604
rect 10284 16552 10300 16604
rect 10352 16552 10368 16604
rect 10420 16552 11152 16604
rect 11204 16552 11220 16604
rect 11272 16552 11288 16604
rect 11340 16552 11341 16604
rect 187 16539 11341 16552
rect 187 16487 4712 16539
rect 4764 16487 4780 16539
rect 4832 16487 4848 16539
rect 4900 16534 5632 16539
rect 5684 16534 5700 16539
rect 5752 16534 5768 16539
rect 5820 16534 6552 16539
rect 6604 16534 6620 16539
rect 6672 16534 6688 16539
rect 6740 16534 7472 16539
rect 4900 16487 5188 16534
rect 187 16478 5188 16487
rect 5244 16478 5270 16534
rect 5326 16478 5352 16534
rect 5408 16478 5434 16534
rect 5490 16478 5516 16534
rect 5572 16478 5598 16534
rect 5752 16487 5762 16534
rect 5820 16487 5844 16534
rect 5654 16478 5680 16487
rect 5736 16478 5762 16487
rect 5818 16478 5844 16487
rect 5900 16478 5926 16534
rect 5982 16478 6008 16534
rect 6064 16478 6090 16534
rect 6146 16478 6172 16534
rect 6228 16478 6254 16534
rect 6310 16478 6336 16534
rect 6392 16478 6418 16534
rect 6474 16478 6500 16534
rect 6740 16487 6746 16534
rect 6556 16478 6582 16487
rect 6638 16478 6664 16487
rect 6720 16478 6746 16487
rect 6802 16478 6828 16534
rect 6884 16478 6909 16534
rect 6965 16478 6990 16534
rect 7046 16478 7071 16534
rect 7127 16478 7152 16534
rect 7208 16478 7233 16534
rect 7289 16478 7314 16534
rect 7370 16487 7472 16534
rect 7524 16487 7540 16539
rect 7592 16487 7608 16539
rect 7660 16487 8392 16539
rect 8444 16487 8460 16539
rect 8512 16487 8528 16539
rect 8580 16487 9312 16539
rect 9364 16487 9380 16539
rect 9432 16487 9448 16539
rect 9500 16487 10232 16539
rect 10284 16487 10300 16539
rect 10352 16487 10368 16539
rect 10420 16487 11152 16539
rect 11204 16487 11220 16539
rect 11272 16487 11288 16539
rect 11340 16487 11341 16539
rect 7370 16478 11341 16487
rect 187 16474 11341 16478
rect 187 16422 4712 16474
rect 4764 16422 4780 16474
rect 4832 16422 4848 16474
rect 4900 16454 5632 16474
rect 5684 16454 5700 16474
rect 5752 16454 5768 16474
rect 5820 16454 6552 16474
rect 6604 16454 6620 16474
rect 6672 16454 6688 16474
rect 6740 16454 7472 16474
rect 4900 16422 5188 16454
rect 187 16409 5188 16422
rect 187 16357 4712 16409
rect 4764 16357 4780 16409
rect 4832 16357 4848 16409
rect 4900 16398 5188 16409
rect 5244 16398 5270 16454
rect 5326 16398 5352 16454
rect 5408 16398 5434 16454
rect 5490 16398 5516 16454
rect 5572 16398 5598 16454
rect 5752 16422 5762 16454
rect 5820 16422 5844 16454
rect 5654 16409 5680 16422
rect 5736 16409 5762 16422
rect 5818 16409 5844 16422
rect 5752 16398 5762 16409
rect 5820 16398 5844 16409
rect 5900 16398 5926 16454
rect 5982 16398 6008 16454
rect 6064 16398 6090 16454
rect 6146 16398 6172 16454
rect 6228 16398 6254 16454
rect 6310 16398 6336 16454
rect 6392 16398 6418 16454
rect 6474 16398 6500 16454
rect 6740 16422 6746 16454
rect 6556 16409 6582 16422
rect 6638 16409 6664 16422
rect 6720 16409 6746 16422
rect 6740 16398 6746 16409
rect 6802 16398 6828 16454
rect 6884 16398 6909 16454
rect 6965 16398 6990 16454
rect 7046 16398 7071 16454
rect 7127 16398 7152 16454
rect 7208 16398 7233 16454
rect 7289 16398 7314 16454
rect 7370 16422 7472 16454
rect 7524 16422 7540 16474
rect 7592 16422 7608 16474
rect 7660 16422 8392 16474
rect 8444 16422 8460 16474
rect 8512 16422 8528 16474
rect 8580 16422 9312 16474
rect 9364 16422 9380 16474
rect 9432 16422 9448 16474
rect 9500 16422 10232 16474
rect 10284 16422 10300 16474
rect 10352 16422 10368 16474
rect 10420 16422 11152 16474
rect 11204 16422 11220 16474
rect 11272 16422 11288 16474
rect 11340 16422 11341 16474
rect 7370 16409 11341 16422
rect 7370 16398 7472 16409
rect 4900 16374 5632 16398
rect 5684 16374 5700 16398
rect 5752 16374 5768 16398
rect 5820 16374 6552 16398
rect 6604 16374 6620 16398
rect 6672 16374 6688 16398
rect 6740 16374 7472 16398
rect 4900 16357 5188 16374
rect 187 16344 5188 16357
rect 187 16292 4712 16344
rect 4764 16292 4780 16344
rect 4832 16292 4848 16344
rect 4900 16318 5188 16344
rect 5244 16318 5270 16374
rect 5326 16318 5352 16374
rect 5408 16318 5434 16374
rect 5490 16318 5516 16374
rect 5572 16318 5598 16374
rect 5752 16357 5762 16374
rect 5820 16357 5844 16374
rect 5654 16344 5680 16357
rect 5736 16344 5762 16357
rect 5818 16344 5844 16357
rect 5752 16318 5762 16344
rect 5820 16318 5844 16344
rect 5900 16318 5926 16374
rect 5982 16318 6008 16374
rect 6064 16318 6090 16374
rect 6146 16318 6172 16374
rect 6228 16318 6254 16374
rect 6310 16318 6336 16374
rect 6392 16318 6418 16374
rect 6474 16318 6500 16374
rect 6740 16357 6746 16374
rect 6556 16344 6582 16357
rect 6638 16344 6664 16357
rect 6720 16344 6746 16357
rect 6740 16318 6746 16344
rect 6802 16318 6828 16374
rect 6884 16318 6909 16374
rect 6965 16318 6990 16374
rect 7046 16318 7071 16374
rect 7127 16318 7152 16374
rect 7208 16318 7233 16374
rect 7289 16318 7314 16374
rect 7370 16357 7472 16374
rect 7524 16357 7540 16409
rect 7592 16357 7608 16409
rect 7660 16357 8392 16409
rect 8444 16357 8460 16409
rect 8512 16357 8528 16409
rect 8580 16357 9312 16409
rect 9364 16357 9380 16409
rect 9432 16357 9448 16409
rect 9500 16357 10232 16409
rect 10284 16357 10300 16409
rect 10352 16357 10368 16409
rect 10420 16357 11152 16409
rect 11204 16357 11220 16409
rect 11272 16357 11288 16409
rect 11340 16357 11341 16409
rect 7370 16344 11341 16357
rect 7370 16318 7472 16344
rect 4900 16294 5632 16318
rect 5684 16294 5700 16318
rect 5752 16294 5768 16318
rect 5820 16294 6552 16318
rect 6604 16294 6620 16318
rect 6672 16294 6688 16318
rect 6740 16294 7472 16318
rect 4900 16292 5188 16294
rect 187 16279 5188 16292
rect 187 16227 4712 16279
rect 4764 16227 4780 16279
rect 4832 16227 4848 16279
rect 4900 16238 5188 16279
rect 5244 16238 5270 16294
rect 5326 16238 5352 16294
rect 5408 16238 5434 16294
rect 5490 16238 5516 16294
rect 5572 16238 5598 16294
rect 5752 16292 5762 16294
rect 5820 16292 5844 16294
rect 5654 16279 5680 16292
rect 5736 16279 5762 16292
rect 5818 16279 5844 16292
rect 5752 16238 5762 16279
rect 5820 16238 5844 16279
rect 5900 16238 5926 16294
rect 5982 16238 6008 16294
rect 6064 16238 6090 16294
rect 6146 16238 6172 16294
rect 6228 16238 6254 16294
rect 6310 16238 6336 16294
rect 6392 16238 6418 16294
rect 6474 16238 6500 16294
rect 6740 16292 6746 16294
rect 6556 16279 6582 16292
rect 6638 16279 6664 16292
rect 6720 16279 6746 16292
rect 6740 16238 6746 16279
rect 6802 16238 6828 16294
rect 6884 16238 6909 16294
rect 6965 16238 6990 16294
rect 7046 16238 7071 16294
rect 7127 16238 7152 16294
rect 7208 16238 7233 16294
rect 7289 16238 7314 16294
rect 7370 16292 7472 16294
rect 7524 16292 7540 16344
rect 7592 16292 7608 16344
rect 7660 16292 8392 16344
rect 8444 16292 8460 16344
rect 8512 16292 8528 16344
rect 8580 16292 9312 16344
rect 9364 16292 9380 16344
rect 9432 16292 9448 16344
rect 9500 16292 10232 16344
rect 10284 16292 10300 16344
rect 10352 16292 10368 16344
rect 10420 16292 11152 16344
rect 11204 16292 11220 16344
rect 11272 16292 11288 16344
rect 11340 16292 11341 16344
rect 7370 16279 11341 16292
rect 7370 16238 7472 16279
rect 4900 16227 5632 16238
rect 5684 16227 5700 16238
rect 5752 16227 5768 16238
rect 5820 16227 6552 16238
rect 6604 16227 6620 16238
rect 6672 16227 6688 16238
rect 6740 16227 7472 16238
rect 7524 16227 7540 16279
rect 7592 16227 7608 16279
rect 7660 16227 8392 16279
rect 8444 16227 8460 16279
rect 8512 16227 8528 16279
rect 8580 16227 9312 16279
rect 9364 16227 9380 16279
rect 9432 16227 9448 16279
rect 9500 16227 10232 16279
rect 10284 16227 10300 16279
rect 10352 16227 10368 16279
rect 10420 16227 11152 16279
rect 11204 16227 11220 16279
rect 11272 16227 11288 16279
rect 11340 16227 11341 16279
rect 187 16214 11341 16227
rect 187 16162 4712 16214
rect 4764 16162 4780 16214
rect 4832 16162 4848 16214
rect 4900 16162 5188 16214
rect 187 16158 5188 16162
rect 5244 16158 5270 16214
rect 5326 16158 5352 16214
rect 5408 16158 5434 16214
rect 5490 16158 5516 16214
rect 5572 16158 5598 16214
rect 5752 16162 5762 16214
rect 5820 16162 5844 16214
rect 5654 16158 5680 16162
rect 5736 16158 5762 16162
rect 5818 16158 5844 16162
rect 5900 16158 5926 16214
rect 5982 16158 6008 16214
rect 6064 16158 6090 16214
rect 6146 16158 6172 16214
rect 6228 16158 6254 16214
rect 6310 16158 6336 16214
rect 6392 16158 6418 16214
rect 6474 16158 6500 16214
rect 6740 16162 6746 16214
rect 6556 16158 6582 16162
rect 6638 16158 6664 16162
rect 6720 16158 6746 16162
rect 6802 16158 6828 16214
rect 6884 16158 6909 16214
rect 6965 16158 6990 16214
rect 7046 16158 7071 16214
rect 7127 16158 7152 16214
rect 7208 16158 7233 16214
rect 7289 16158 7314 16214
rect 7370 16162 7472 16214
rect 7524 16162 7540 16214
rect 7592 16162 7608 16214
rect 7660 16162 8392 16214
rect 8444 16162 8460 16214
rect 8512 16162 8528 16214
rect 8580 16162 9312 16214
rect 9364 16162 9380 16214
rect 9432 16162 9448 16214
rect 9500 16162 10232 16214
rect 10284 16162 10300 16214
rect 10352 16162 10368 16214
rect 10420 16162 11152 16214
rect 11204 16162 11220 16214
rect 11272 16162 11288 16214
rect 11340 16162 11341 16214
rect 7370 16158 11341 16162
rect 187 16156 11341 16158
rect 187 13599 2824 16156
tri 2824 15448 3532 16156 nw
tri 11511 15831 12222 16542 se
rect 12222 15831 14858 18691
rect 4964 15829 14858 15831
rect 4964 15825 7587 15829
rect 4964 15773 5201 15825
rect 5253 15773 5279 15825
rect 5331 15773 6121 15825
rect 6173 15773 6199 15825
rect 6251 15773 7041 15825
rect 7093 15773 7119 15825
rect 7171 15773 7587 15825
rect 7643 15773 7669 15829
rect 7725 15773 7751 15829
rect 7807 15773 7833 15829
rect 7889 15773 7915 15829
rect 7971 15825 7997 15829
rect 8053 15825 8079 15829
rect 8135 15773 8161 15829
rect 8217 15773 8243 15829
rect 8299 15773 8325 15829
rect 8381 15773 8407 15829
rect 8463 15773 8489 15829
rect 8545 15773 8571 15829
rect 8627 15773 8653 15829
rect 8709 15773 8735 15829
rect 8791 15773 8817 15829
rect 8873 15825 8899 15829
rect 8955 15825 8981 15829
rect 8873 15773 8881 15825
rect 8955 15773 8959 15825
rect 9037 15773 9063 15829
rect 9119 15773 9145 15829
rect 9201 15773 9227 15829
rect 9283 15773 9308 15829
rect 9364 15773 9389 15829
rect 9445 15773 9470 15829
rect 9526 15773 9551 15829
rect 9607 15773 9632 15829
rect 9688 15773 9713 15829
rect 9769 15825 14858 15829
rect 9769 15773 9801 15825
rect 9853 15773 9879 15825
rect 9931 15773 10721 15825
rect 10773 15773 10799 15825
rect 10851 15773 11641 15825
rect 11693 15773 11719 15825
rect 11771 15773 12561 15825
rect 12613 15773 12639 15825
rect 12691 15773 14858 15825
rect 4964 15761 14858 15773
rect 4964 15709 5201 15761
rect 5253 15709 5279 15761
rect 5331 15709 6121 15761
rect 6173 15709 6199 15761
rect 6251 15709 7041 15761
rect 7093 15709 7119 15761
rect 7171 15749 7961 15761
rect 8013 15749 8039 15761
rect 8091 15749 8881 15761
rect 8933 15749 8959 15761
rect 9011 15749 9801 15761
rect 7171 15709 7587 15749
rect 4964 15697 7587 15709
rect 4964 15645 5201 15697
rect 5253 15645 5279 15697
rect 5331 15645 6121 15697
rect 6173 15645 6199 15697
rect 6251 15645 7041 15697
rect 7093 15645 7119 15697
rect 7171 15693 7587 15697
rect 7643 15693 7669 15749
rect 7725 15693 7751 15749
rect 7807 15693 7833 15749
rect 7889 15693 7915 15749
rect 7971 15697 7997 15709
rect 8053 15697 8079 15709
rect 8135 15693 8161 15749
rect 8217 15693 8243 15749
rect 8299 15693 8325 15749
rect 8381 15693 8407 15749
rect 8463 15693 8489 15749
rect 8545 15693 8571 15749
rect 8627 15693 8653 15749
rect 8709 15693 8735 15749
rect 8791 15693 8817 15749
rect 8873 15709 8881 15749
rect 8955 15709 8959 15749
rect 8873 15697 8899 15709
rect 8955 15697 8981 15709
rect 8873 15693 8881 15697
rect 8955 15693 8959 15697
rect 9037 15693 9063 15749
rect 9119 15693 9145 15749
rect 9201 15693 9227 15749
rect 9283 15693 9308 15749
rect 9364 15693 9389 15749
rect 9445 15693 9470 15749
rect 9526 15693 9551 15749
rect 9607 15693 9632 15749
rect 9688 15693 9713 15749
rect 9769 15709 9801 15749
rect 9853 15709 9879 15761
rect 9931 15709 10721 15761
rect 10773 15709 10799 15761
rect 10851 15709 11641 15761
rect 11693 15709 11719 15761
rect 11771 15709 12561 15761
rect 12613 15709 12639 15761
rect 12691 15709 14858 15761
rect 9769 15697 14858 15709
rect 9769 15693 9801 15697
rect 7171 15669 7961 15693
rect 8013 15669 8039 15693
rect 8091 15669 8881 15693
rect 8933 15669 8959 15693
rect 9011 15669 9801 15693
rect 7171 15645 7587 15669
rect 4964 15633 7587 15645
rect 4964 15581 5201 15633
rect 5253 15581 5279 15633
rect 5331 15581 6121 15633
rect 6173 15581 6199 15633
rect 6251 15581 7041 15633
rect 7093 15581 7119 15633
rect 7171 15613 7587 15633
rect 7643 15613 7669 15669
rect 7725 15613 7751 15669
rect 7807 15613 7833 15669
rect 7889 15613 7915 15669
rect 7971 15633 7997 15645
rect 8053 15633 8079 15645
rect 8135 15613 8161 15669
rect 8217 15613 8243 15669
rect 8299 15613 8325 15669
rect 8381 15613 8407 15669
rect 8463 15613 8489 15669
rect 8545 15613 8571 15669
rect 8627 15613 8653 15669
rect 8709 15613 8735 15669
rect 8791 15613 8817 15669
rect 8873 15645 8881 15669
rect 8955 15645 8959 15669
rect 8873 15633 8899 15645
rect 8955 15633 8981 15645
rect 8873 15613 8881 15633
rect 8955 15613 8959 15633
rect 9037 15613 9063 15669
rect 9119 15613 9145 15669
rect 9201 15613 9227 15669
rect 9283 15613 9308 15669
rect 9364 15613 9389 15669
rect 9445 15613 9470 15669
rect 9526 15613 9551 15669
rect 9607 15613 9632 15669
rect 9688 15613 9713 15669
rect 9769 15645 9801 15669
rect 9853 15645 9879 15697
rect 9931 15645 10721 15697
rect 10773 15645 10799 15697
rect 10851 15645 11641 15697
rect 11693 15645 11719 15697
rect 11771 15645 12561 15697
rect 12613 15645 12639 15697
rect 12691 15645 14858 15697
rect 9769 15633 14858 15645
rect 9769 15613 9801 15633
rect 7171 15589 7961 15613
rect 8013 15589 8039 15613
rect 8091 15589 8881 15613
rect 8933 15589 8959 15613
rect 9011 15589 9801 15613
rect 7171 15581 7587 15589
rect 4964 15569 7587 15581
rect 4964 15517 5201 15569
rect 5253 15517 5279 15569
rect 5331 15517 6121 15569
rect 6173 15517 6199 15569
rect 6251 15517 7041 15569
rect 7093 15517 7119 15569
rect 7171 15533 7587 15569
rect 7643 15533 7669 15589
rect 7725 15533 7751 15589
rect 7807 15533 7833 15589
rect 7889 15533 7915 15589
rect 7971 15569 7997 15581
rect 8053 15569 8079 15581
rect 8135 15533 8161 15589
rect 8217 15533 8243 15589
rect 8299 15533 8325 15589
rect 8381 15533 8407 15589
rect 8463 15533 8489 15589
rect 8545 15533 8571 15589
rect 8627 15533 8653 15589
rect 8709 15533 8735 15589
rect 8791 15533 8817 15589
rect 8873 15581 8881 15589
rect 8955 15581 8959 15589
rect 8873 15569 8899 15581
rect 8955 15569 8981 15581
rect 8873 15533 8881 15569
rect 8955 15533 8959 15569
rect 9037 15533 9063 15589
rect 9119 15533 9145 15589
rect 9201 15533 9227 15589
rect 9283 15533 9308 15589
rect 9364 15533 9389 15589
rect 9445 15533 9470 15589
rect 9526 15533 9551 15589
rect 9607 15533 9632 15589
rect 9688 15533 9713 15589
rect 9769 15581 9801 15589
rect 9853 15581 9879 15633
rect 9931 15581 10721 15633
rect 10773 15581 10799 15633
rect 10851 15581 11641 15633
rect 11693 15581 11719 15633
rect 11771 15581 12561 15633
rect 12613 15581 12639 15633
rect 12691 15581 14858 15633
rect 9769 15569 14858 15581
rect 9769 15533 9801 15569
rect 7171 15517 7961 15533
rect 8013 15517 8039 15533
rect 8091 15517 8881 15533
rect 8933 15517 8959 15533
rect 9011 15517 9801 15533
rect 9853 15517 9879 15569
rect 9931 15517 10721 15569
rect 10773 15517 10799 15569
rect 10851 15517 11641 15569
rect 11693 15517 11719 15569
rect 11771 15517 12561 15569
rect 12613 15517 12639 15569
rect 12691 15517 14858 15569
rect 4964 15509 14858 15517
rect 4964 15505 7587 15509
rect 4964 15453 5201 15505
rect 5253 15453 5279 15505
rect 5331 15453 6121 15505
rect 6173 15453 6199 15505
rect 6251 15453 7041 15505
rect 7093 15453 7119 15505
rect 7171 15453 7587 15505
rect 7643 15453 7669 15509
rect 7725 15453 7751 15509
rect 7807 15453 7833 15509
rect 7889 15453 7915 15509
rect 7971 15505 7997 15509
rect 8053 15505 8079 15509
rect 8135 15453 8161 15509
rect 8217 15453 8243 15509
rect 8299 15453 8325 15509
rect 8381 15453 8407 15509
rect 8463 15453 8489 15509
rect 8545 15453 8571 15509
rect 8627 15453 8653 15509
rect 8709 15453 8735 15509
rect 8791 15453 8817 15509
rect 8873 15505 8899 15509
rect 8955 15505 8981 15509
rect 8873 15453 8881 15505
rect 8955 15453 8959 15505
rect 9037 15453 9063 15509
rect 9119 15453 9145 15509
rect 9201 15453 9227 15509
rect 9283 15453 9308 15509
rect 9364 15453 9389 15509
rect 9445 15453 9470 15509
rect 9526 15453 9551 15509
rect 9607 15453 9632 15509
rect 9688 15453 9713 15509
rect 9769 15505 14858 15509
rect 9769 15453 9801 15505
rect 9853 15453 9879 15505
rect 9931 15453 10721 15505
rect 10773 15453 10799 15505
rect 10851 15453 11641 15505
rect 11693 15453 11719 15505
rect 11771 15453 12561 15505
rect 12613 15453 12639 15505
rect 12691 15453 14858 15505
rect 4964 15441 14858 15453
rect 4964 15389 5201 15441
rect 5253 15389 5279 15441
rect 5331 15389 6121 15441
rect 6173 15389 6199 15441
rect 6251 15389 7041 15441
rect 7093 15389 7119 15441
rect 7171 15429 7961 15441
rect 8013 15429 8039 15441
rect 8091 15429 8881 15441
rect 8933 15429 8959 15441
rect 9011 15429 9801 15441
rect 7171 15389 7587 15429
rect 4964 15377 7587 15389
rect 4964 15325 5201 15377
rect 5253 15325 5279 15377
rect 5331 15325 6121 15377
rect 6173 15325 6199 15377
rect 6251 15325 7041 15377
rect 7093 15325 7119 15377
rect 7171 15373 7587 15377
rect 7643 15373 7669 15429
rect 7725 15373 7751 15429
rect 7807 15373 7833 15429
rect 7889 15373 7915 15429
rect 7971 15377 7997 15389
rect 8053 15377 8079 15389
rect 8135 15373 8161 15429
rect 8217 15373 8243 15429
rect 8299 15373 8325 15429
rect 8381 15373 8407 15429
rect 8463 15373 8489 15429
rect 8545 15373 8571 15429
rect 8627 15373 8653 15429
rect 8709 15373 8735 15429
rect 8791 15373 8817 15429
rect 8873 15389 8881 15429
rect 8955 15389 8959 15429
rect 8873 15377 8899 15389
rect 8955 15377 8981 15389
rect 8873 15373 8881 15377
rect 8955 15373 8959 15377
rect 9037 15373 9063 15429
rect 9119 15373 9145 15429
rect 9201 15373 9227 15429
rect 9283 15373 9308 15429
rect 9364 15373 9389 15429
rect 9445 15373 9470 15429
rect 9526 15373 9551 15429
rect 9607 15373 9632 15429
rect 9688 15373 9713 15429
rect 9769 15389 9801 15429
rect 9853 15389 9879 15441
rect 9931 15389 10721 15441
rect 10773 15389 10799 15441
rect 10851 15389 11641 15441
rect 11693 15389 11719 15441
rect 11771 15389 12561 15441
rect 12613 15389 12639 15441
rect 12691 15389 14858 15441
rect 9769 15377 14858 15389
rect 9769 15373 9801 15377
rect 7171 15349 7961 15373
rect 8013 15349 8039 15373
rect 8091 15349 8881 15373
rect 8933 15349 8959 15373
rect 9011 15349 9801 15373
rect 7171 15325 7587 15349
rect 4964 15313 7587 15325
rect 4964 15261 5201 15313
rect 5253 15261 5279 15313
rect 5331 15261 6121 15313
rect 6173 15261 6199 15313
rect 6251 15261 7041 15313
rect 7093 15261 7119 15313
rect 7171 15293 7587 15313
rect 7643 15293 7669 15349
rect 7725 15293 7751 15349
rect 7807 15293 7833 15349
rect 7889 15293 7915 15349
rect 7971 15313 7997 15325
rect 8053 15313 8079 15325
rect 8135 15293 8161 15349
rect 8217 15293 8243 15349
rect 8299 15293 8325 15349
rect 8381 15293 8407 15349
rect 8463 15293 8489 15349
rect 8545 15293 8571 15349
rect 8627 15293 8653 15349
rect 8709 15293 8735 15349
rect 8791 15293 8817 15349
rect 8873 15325 8881 15349
rect 8955 15325 8959 15349
rect 8873 15313 8899 15325
rect 8955 15313 8981 15325
rect 8873 15293 8881 15313
rect 8955 15293 8959 15313
rect 9037 15293 9063 15349
rect 9119 15293 9145 15349
rect 9201 15293 9227 15349
rect 9283 15293 9308 15349
rect 9364 15293 9389 15349
rect 9445 15293 9470 15349
rect 9526 15293 9551 15349
rect 9607 15293 9632 15349
rect 9688 15293 9713 15349
rect 9769 15325 9801 15349
rect 9853 15325 9879 15377
rect 9931 15325 10721 15377
rect 10773 15325 10799 15377
rect 10851 15325 11641 15377
rect 11693 15325 11719 15377
rect 11771 15325 12561 15377
rect 12613 15325 12639 15377
rect 12691 15325 14858 15377
rect 9769 15313 14858 15325
rect 9769 15293 9801 15313
rect 7171 15269 7961 15293
rect 8013 15269 8039 15293
rect 8091 15269 8881 15293
rect 8933 15269 8959 15293
rect 9011 15269 9801 15293
rect 7171 15261 7587 15269
rect 4964 15249 7587 15261
rect 4964 15197 5201 15249
rect 5253 15197 5279 15249
rect 5331 15197 6121 15249
rect 6173 15197 6199 15249
rect 6251 15197 7041 15249
rect 7093 15197 7119 15249
rect 7171 15213 7587 15249
rect 7643 15213 7669 15269
rect 7725 15213 7751 15269
rect 7807 15213 7833 15269
rect 7889 15213 7915 15269
rect 7971 15249 7997 15261
rect 8053 15249 8079 15261
rect 8135 15213 8161 15269
rect 8217 15213 8243 15269
rect 8299 15213 8325 15269
rect 8381 15213 8407 15269
rect 8463 15213 8489 15269
rect 8545 15213 8571 15269
rect 8627 15213 8653 15269
rect 8709 15213 8735 15269
rect 8791 15213 8817 15269
rect 8873 15261 8881 15269
rect 8955 15261 8959 15269
rect 8873 15249 8899 15261
rect 8955 15249 8981 15261
rect 8873 15213 8881 15249
rect 8955 15213 8959 15249
rect 9037 15213 9063 15269
rect 9119 15213 9145 15269
rect 9201 15213 9227 15269
rect 9283 15213 9308 15269
rect 9364 15213 9389 15269
rect 9445 15213 9470 15269
rect 9526 15213 9551 15269
rect 9607 15213 9632 15269
rect 9688 15213 9713 15269
rect 9769 15261 9801 15269
rect 9853 15261 9879 15313
rect 9931 15261 10721 15313
rect 10773 15261 10799 15313
rect 10851 15261 11641 15313
rect 11693 15261 11719 15313
rect 11771 15261 12561 15313
rect 12613 15261 12639 15313
rect 12691 15261 14858 15313
rect 9769 15249 14858 15261
rect 9769 15213 9801 15249
rect 7171 15197 7961 15213
rect 8013 15197 8039 15213
rect 8091 15197 8881 15213
rect 8933 15197 8959 15213
rect 9011 15197 9801 15213
rect 9853 15197 9879 15249
rect 9931 15197 10721 15249
rect 10773 15197 10799 15249
rect 10851 15197 11641 15249
rect 11693 15197 11719 15249
rect 11771 15197 12561 15249
rect 12613 15197 12639 15249
rect 12691 15197 14858 15249
rect 4964 15189 14858 15197
rect 4964 15185 7587 15189
rect 4964 15133 5201 15185
rect 5253 15133 5279 15185
rect 5331 15133 6121 15185
rect 6173 15133 6199 15185
rect 6251 15133 7041 15185
rect 7093 15133 7119 15185
rect 7171 15133 7587 15185
rect 7643 15133 7669 15189
rect 7725 15133 7751 15189
rect 7807 15133 7833 15189
rect 7889 15133 7915 15189
rect 7971 15185 7997 15189
rect 8053 15185 8079 15189
rect 8135 15133 8161 15189
rect 8217 15133 8243 15189
rect 8299 15133 8325 15189
rect 8381 15133 8407 15189
rect 8463 15133 8489 15189
rect 8545 15133 8571 15189
rect 8627 15133 8653 15189
rect 8709 15133 8735 15189
rect 8791 15133 8817 15189
rect 8873 15185 8899 15189
rect 8955 15185 8981 15189
rect 8873 15133 8881 15185
rect 8955 15133 8959 15185
rect 9037 15133 9063 15189
rect 9119 15133 9145 15189
rect 9201 15133 9227 15189
rect 9283 15133 9308 15189
rect 9364 15133 9389 15189
rect 9445 15133 9470 15189
rect 9526 15133 9551 15189
rect 9607 15133 9632 15189
rect 9688 15133 9713 15189
rect 9769 15185 14858 15189
rect 9769 15133 9801 15185
rect 9853 15133 9879 15185
rect 9931 15133 10721 15185
rect 10773 15133 10799 15185
rect 10851 15133 11641 15185
rect 11693 15133 11719 15185
rect 11771 15133 12561 15185
rect 12613 15133 12639 15185
rect 12691 15133 14858 15185
tri 4724 14883 4964 15123 se
rect 4964 15121 14858 15133
rect 4964 15069 5201 15121
rect 5253 15069 5279 15121
rect 5331 15069 6121 15121
rect 6173 15069 6199 15121
rect 6251 15069 7041 15121
rect 7093 15069 7119 15121
rect 7171 15109 7961 15121
rect 8013 15109 8039 15121
rect 8091 15109 8881 15121
rect 8933 15109 8959 15121
rect 9011 15109 9801 15121
rect 7171 15069 7587 15109
rect 4964 15057 7587 15069
rect 4964 15005 5201 15057
rect 5253 15005 5279 15057
rect 5331 15005 6121 15057
rect 6173 15005 6199 15057
rect 6251 15005 7041 15057
rect 7093 15005 7119 15057
rect 7171 15053 7587 15057
rect 7643 15053 7669 15109
rect 7725 15053 7751 15109
rect 7807 15053 7833 15109
rect 7889 15053 7915 15109
rect 7971 15057 7997 15069
rect 8053 15057 8079 15069
rect 8135 15053 8161 15109
rect 8217 15053 8243 15109
rect 8299 15053 8325 15109
rect 8381 15053 8407 15109
rect 8463 15053 8489 15109
rect 8545 15053 8571 15109
rect 8627 15053 8653 15109
rect 8709 15053 8735 15109
rect 8791 15053 8817 15109
rect 8873 15069 8881 15109
rect 8955 15069 8959 15109
rect 8873 15057 8899 15069
rect 8955 15057 8981 15069
rect 8873 15053 8881 15057
rect 8955 15053 8959 15057
rect 9037 15053 9063 15109
rect 9119 15053 9145 15109
rect 9201 15053 9227 15109
rect 9283 15053 9308 15109
rect 9364 15053 9389 15109
rect 9445 15053 9470 15109
rect 9526 15053 9551 15109
rect 9607 15053 9632 15109
rect 9688 15053 9713 15109
rect 9769 15069 9801 15109
rect 9853 15069 9879 15121
rect 9931 15069 10721 15121
rect 10773 15069 10799 15121
rect 10851 15069 11641 15121
rect 11693 15069 11719 15121
rect 11771 15069 12561 15121
rect 12613 15069 12639 15121
rect 12691 15069 14858 15121
rect 9769 15057 14858 15069
rect 9769 15053 9801 15057
rect 7171 15029 7961 15053
rect 8013 15029 8039 15053
rect 8091 15029 8881 15053
rect 8933 15029 8959 15053
rect 9011 15029 9801 15053
rect 7171 15005 7587 15029
rect 4964 14993 7587 15005
rect 4964 14941 5201 14993
rect 5253 14941 5279 14993
rect 5331 14941 6121 14993
rect 6173 14941 6199 14993
rect 6251 14941 7041 14993
rect 7093 14941 7119 14993
rect 7171 14973 7587 14993
rect 7643 14973 7669 15029
rect 7725 14973 7751 15029
rect 7807 14973 7833 15029
rect 7889 14973 7915 15029
rect 7971 14993 7997 15005
rect 8053 14993 8079 15005
rect 8135 14973 8161 15029
rect 8217 14973 8243 15029
rect 8299 14973 8325 15029
rect 8381 14973 8407 15029
rect 8463 14973 8489 15029
rect 8545 14973 8571 15029
rect 8627 14973 8653 15029
rect 8709 14973 8735 15029
rect 8791 14973 8817 15029
rect 8873 15005 8881 15029
rect 8955 15005 8959 15029
rect 8873 14993 8899 15005
rect 8955 14993 8981 15005
rect 8873 14973 8881 14993
rect 8955 14973 8959 14993
rect 9037 14973 9063 15029
rect 9119 14973 9145 15029
rect 9201 14973 9227 15029
rect 9283 14973 9308 15029
rect 9364 14973 9389 15029
rect 9445 14973 9470 15029
rect 9526 14973 9551 15029
rect 9607 14973 9632 15029
rect 9688 14973 9713 15029
rect 9769 15005 9801 15029
rect 9853 15005 9879 15057
rect 9931 15005 10721 15057
rect 10773 15005 10799 15057
rect 10851 15005 11641 15057
rect 11693 15005 11719 15057
rect 11771 15005 12561 15057
rect 12613 15005 12639 15057
rect 12691 15005 14858 15057
rect 9769 14993 14858 15005
rect 9769 14973 9801 14993
rect 7171 14949 7961 14973
rect 8013 14949 8039 14973
rect 8091 14949 8881 14973
rect 8933 14949 8959 14973
rect 9011 14949 9801 14973
rect 7171 14941 7587 14949
rect 4964 14929 7587 14941
rect 4964 14883 5201 14929
rect 3682 14831 3688 14883
rect 3740 14831 3754 14883
rect 3806 14877 5201 14883
rect 5253 14877 5279 14929
rect 5331 14877 6121 14929
rect 6173 14877 6199 14929
rect 6251 14877 7041 14929
rect 7093 14877 7119 14929
rect 7171 14893 7587 14929
rect 7643 14893 7669 14949
rect 7725 14893 7751 14949
rect 7807 14893 7833 14949
rect 7889 14893 7915 14949
rect 7971 14929 7997 14941
rect 8053 14929 8079 14941
rect 8135 14893 8161 14949
rect 8217 14893 8243 14949
rect 8299 14893 8325 14949
rect 8381 14893 8407 14949
rect 8463 14893 8489 14949
rect 8545 14893 8571 14949
rect 8627 14893 8653 14949
rect 8709 14893 8735 14949
rect 8791 14893 8817 14949
rect 8873 14941 8881 14949
rect 8955 14941 8959 14949
rect 8873 14929 8899 14941
rect 8955 14929 8981 14941
rect 8873 14893 8881 14929
rect 8955 14893 8959 14929
rect 9037 14893 9063 14949
rect 9119 14893 9145 14949
rect 9201 14893 9227 14949
rect 9283 14893 9308 14949
rect 9364 14893 9389 14949
rect 9445 14893 9470 14949
rect 9526 14893 9551 14949
rect 9607 14893 9632 14949
rect 9688 14893 9713 14949
rect 9769 14941 9801 14949
rect 9853 14941 9879 14993
rect 9931 14941 10721 14993
rect 10773 14941 10799 14993
rect 10851 14941 11641 14993
rect 11693 14941 11719 14993
rect 11771 14941 12561 14993
rect 12613 14941 12639 14993
rect 12691 14941 14858 14993
rect 9769 14929 14858 14941
rect 9769 14893 9801 14929
rect 7171 14877 7961 14893
rect 8013 14877 8039 14893
rect 8091 14877 8881 14893
rect 8933 14877 8959 14893
rect 9011 14877 9801 14893
rect 9853 14877 9879 14929
rect 9931 14877 10721 14929
rect 10773 14877 10799 14929
rect 10851 14877 11641 14929
rect 11693 14877 11719 14929
rect 11771 14877 12561 14929
rect 12613 14877 12639 14929
rect 12691 14877 14858 14929
rect 3806 14869 14858 14877
rect 3806 14864 7587 14869
rect 3806 14831 5201 14864
rect 3353 14650 3359 14702
rect 3411 14650 3448 14702
rect 3500 14650 3506 14702
tri 3353 14617 3386 14650 ne
rect 3386 14617 3434 14650
tri 3434 14617 3467 14650 nw
tri 3386 14616 3387 14617 ne
tri 2824 13599 3230 14005 sw
tri 3361 13651 3387 13677 se
rect 3387 13651 3433 14617
tri 3433 14616 3434 14617 nw
tri 4730 14597 4964 14831 ne
rect 4964 14812 5201 14831
rect 5253 14812 5279 14864
rect 5331 14812 6121 14864
rect 6173 14812 6199 14864
rect 6251 14812 7041 14864
rect 7093 14812 7119 14864
rect 7171 14813 7587 14864
rect 7643 14813 7669 14869
rect 7725 14813 7751 14869
rect 7807 14813 7833 14869
rect 7889 14813 7915 14869
rect 7971 14864 7997 14869
rect 8053 14864 8079 14869
rect 8135 14813 8161 14869
rect 8217 14813 8243 14869
rect 8299 14813 8325 14869
rect 8381 14813 8407 14869
rect 8463 14813 8489 14869
rect 8545 14813 8571 14869
rect 8627 14813 8653 14869
rect 8709 14813 8735 14869
rect 8791 14813 8817 14869
rect 8873 14864 8899 14869
rect 8955 14864 8981 14869
rect 8873 14813 8881 14864
rect 8955 14813 8959 14864
rect 9037 14813 9063 14869
rect 9119 14813 9145 14869
rect 9201 14813 9227 14869
rect 9283 14813 9308 14869
rect 9364 14813 9389 14869
rect 9445 14813 9470 14869
rect 9526 14813 9551 14869
rect 9607 14813 9632 14869
rect 9688 14813 9713 14869
rect 9769 14864 14858 14869
rect 9769 14813 9801 14864
rect 7171 14812 7961 14813
rect 8013 14812 8039 14813
rect 8091 14812 8881 14813
rect 8933 14812 8959 14813
rect 9011 14812 9801 14813
rect 9853 14812 9879 14864
rect 9931 14812 10721 14864
rect 10773 14812 10799 14864
rect 10851 14812 11641 14864
rect 11693 14812 11719 14864
rect 11771 14812 12561 14864
rect 12613 14812 12639 14864
rect 12691 14812 14858 14864
rect 4964 14799 14858 14812
rect 4964 14747 5201 14799
rect 5253 14747 5279 14799
rect 5331 14747 6121 14799
rect 6173 14747 6199 14799
rect 6251 14747 7041 14799
rect 7093 14747 7119 14799
rect 7171 14789 7961 14799
rect 8013 14789 8039 14799
rect 8091 14789 8881 14799
rect 8933 14789 8959 14799
rect 9011 14789 9801 14799
rect 7171 14747 7587 14789
rect 4964 14734 7587 14747
rect 4964 14682 5201 14734
rect 5253 14682 5279 14734
rect 5331 14682 6121 14734
rect 6173 14682 6199 14734
rect 6251 14682 7041 14734
rect 7093 14682 7119 14734
rect 7171 14733 7587 14734
rect 7643 14733 7669 14789
rect 7725 14733 7751 14789
rect 7807 14733 7833 14789
rect 7889 14733 7915 14789
rect 7971 14734 7997 14747
rect 8053 14734 8079 14747
rect 8135 14733 8161 14789
rect 8217 14733 8243 14789
rect 8299 14733 8325 14789
rect 8381 14733 8407 14789
rect 8463 14733 8489 14789
rect 8545 14733 8571 14789
rect 8627 14733 8653 14789
rect 8709 14733 8735 14789
rect 8791 14733 8817 14789
rect 8873 14747 8881 14789
rect 8955 14747 8959 14789
rect 8873 14734 8899 14747
rect 8955 14734 8981 14747
rect 8873 14733 8881 14734
rect 8955 14733 8959 14734
rect 9037 14733 9063 14789
rect 9119 14733 9145 14789
rect 9201 14733 9227 14789
rect 9283 14733 9308 14789
rect 9364 14733 9389 14789
rect 9445 14733 9470 14789
rect 9526 14733 9551 14789
rect 9607 14733 9632 14789
rect 9688 14733 9713 14789
rect 9769 14747 9801 14789
rect 9853 14747 9879 14799
rect 9931 14747 10721 14799
rect 10773 14747 10799 14799
rect 10851 14747 11641 14799
rect 11693 14747 11719 14799
rect 11771 14747 12561 14799
rect 12613 14747 12639 14799
rect 12691 14747 14858 14799
rect 9769 14734 14858 14747
rect 9769 14733 9801 14734
rect 7171 14709 7961 14733
rect 8013 14709 8039 14733
rect 8091 14709 8881 14733
rect 8933 14709 8959 14733
rect 9011 14709 9801 14733
rect 7171 14682 7587 14709
rect 4964 14669 7587 14682
rect 4964 14617 5201 14669
rect 5253 14617 5279 14669
rect 5331 14617 6121 14669
rect 6173 14617 6199 14669
rect 6251 14617 7041 14669
rect 7093 14617 7119 14669
rect 7171 14653 7587 14669
rect 7643 14653 7669 14709
rect 7725 14653 7751 14709
rect 7807 14653 7833 14709
rect 7889 14653 7915 14709
rect 7971 14669 7997 14682
rect 8053 14669 8079 14682
rect 8135 14653 8161 14709
rect 8217 14653 8243 14709
rect 8299 14653 8325 14709
rect 8381 14653 8407 14709
rect 8463 14653 8489 14709
rect 8545 14653 8571 14709
rect 8627 14653 8653 14709
rect 8709 14653 8735 14709
rect 8791 14653 8817 14709
rect 8873 14682 8881 14709
rect 8955 14682 8959 14709
rect 8873 14669 8899 14682
rect 8955 14669 8981 14682
rect 8873 14653 8881 14669
rect 8955 14653 8959 14669
rect 9037 14653 9063 14709
rect 9119 14653 9145 14709
rect 9201 14653 9227 14709
rect 9283 14653 9308 14709
rect 9364 14653 9389 14709
rect 9445 14653 9470 14709
rect 9526 14653 9551 14709
rect 9607 14653 9632 14709
rect 9688 14653 9713 14709
rect 9769 14682 9801 14709
rect 9853 14682 9879 14734
rect 9931 14682 10721 14734
rect 10773 14682 10799 14734
rect 10851 14682 11641 14734
rect 11693 14682 11719 14734
rect 11771 14682 12561 14734
rect 12613 14682 12639 14734
rect 12691 14682 14858 14734
rect 9769 14669 14858 14682
rect 9769 14653 9801 14669
rect 7171 14629 7961 14653
rect 8013 14629 8039 14653
rect 8091 14629 8881 14653
rect 8933 14629 8959 14653
rect 9011 14629 9801 14653
rect 7171 14617 7587 14629
rect 4964 14604 7587 14617
rect 4964 14552 5201 14604
rect 5253 14552 5279 14604
rect 5331 14552 6121 14604
rect 6173 14552 6199 14604
rect 6251 14552 7041 14604
rect 7093 14552 7119 14604
rect 7171 14573 7587 14604
rect 7643 14573 7669 14629
rect 7725 14573 7751 14629
rect 7807 14573 7833 14629
rect 7889 14573 7915 14629
rect 7971 14604 7997 14617
rect 8053 14604 8079 14617
rect 8135 14573 8161 14629
rect 8217 14573 8243 14629
rect 8299 14573 8325 14629
rect 8381 14573 8407 14629
rect 8463 14573 8489 14629
rect 8545 14573 8571 14629
rect 8627 14573 8653 14629
rect 8709 14573 8735 14629
rect 8791 14573 8817 14629
rect 8873 14617 8881 14629
rect 8955 14617 8959 14629
rect 8873 14604 8899 14617
rect 8955 14604 8981 14617
rect 8873 14573 8881 14604
rect 8955 14573 8959 14604
rect 9037 14573 9063 14629
rect 9119 14573 9145 14629
rect 9201 14573 9227 14629
rect 9283 14573 9308 14629
rect 9364 14573 9389 14629
rect 9445 14573 9470 14629
rect 9526 14573 9551 14629
rect 9607 14573 9632 14629
rect 9688 14573 9713 14629
rect 9769 14617 9801 14629
rect 9853 14617 9879 14669
rect 9931 14617 10721 14669
rect 10773 14617 10799 14669
rect 10851 14617 11641 14669
rect 11693 14617 11719 14669
rect 11771 14617 12561 14669
rect 12613 14617 12639 14669
rect 12691 14617 14858 14669
rect 9769 14604 14858 14617
rect 9769 14573 9801 14604
rect 7171 14552 7961 14573
rect 8013 14552 8039 14573
rect 8091 14552 8881 14573
rect 8933 14552 8959 14573
rect 9011 14552 9801 14573
rect 9853 14552 9879 14604
rect 9931 14552 10721 14604
rect 10773 14552 10799 14604
rect 10851 14552 11641 14604
rect 11693 14552 11719 14604
rect 11771 14552 12561 14604
rect 12613 14552 12639 14604
rect 12691 14552 14858 14604
rect 4964 14549 14858 14552
rect 4964 14539 7587 14549
rect 4964 14487 5201 14539
rect 5253 14487 5279 14539
rect 5331 14487 6121 14539
rect 6173 14487 6199 14539
rect 6251 14487 7041 14539
rect 7093 14487 7119 14539
rect 7171 14493 7587 14539
rect 7643 14493 7669 14549
rect 7725 14493 7751 14549
rect 7807 14493 7833 14549
rect 7889 14493 7915 14549
rect 7971 14539 7997 14549
rect 8053 14539 8079 14549
rect 8135 14493 8161 14549
rect 8217 14493 8243 14549
rect 8299 14493 8325 14549
rect 8381 14493 8407 14549
rect 8463 14493 8489 14549
rect 8545 14493 8571 14549
rect 8627 14493 8653 14549
rect 8709 14493 8735 14549
rect 8791 14493 8817 14549
rect 8873 14539 8899 14549
rect 8955 14539 8981 14549
rect 8873 14493 8881 14539
rect 8955 14493 8959 14539
rect 9037 14493 9063 14549
rect 9119 14493 9145 14549
rect 9201 14493 9227 14549
rect 9283 14493 9308 14549
rect 9364 14493 9389 14549
rect 9445 14493 9470 14549
rect 9526 14493 9551 14549
rect 9607 14493 9632 14549
rect 9688 14493 9713 14549
rect 9769 14539 14858 14549
rect 9769 14493 9801 14539
rect 7171 14487 7961 14493
rect 8013 14487 8039 14493
rect 8091 14487 8881 14493
rect 8933 14487 8959 14493
rect 9011 14487 9801 14493
rect 9853 14487 9879 14539
rect 9931 14487 10721 14539
rect 10773 14487 10799 14539
rect 10851 14487 11641 14539
rect 11693 14487 11719 14539
rect 11771 14487 12561 14539
rect 12613 14487 12639 14539
rect 12691 14487 14858 14539
rect 4964 14474 14858 14487
rect 4964 14422 5201 14474
rect 5253 14422 5279 14474
rect 5331 14422 6121 14474
rect 6173 14422 6199 14474
rect 6251 14422 7041 14474
rect 7093 14422 7119 14474
rect 7171 14469 7961 14474
rect 8013 14469 8039 14474
rect 8091 14469 8881 14474
rect 8933 14469 8959 14474
rect 9011 14469 9801 14474
rect 7171 14422 7587 14469
rect 4964 14413 7587 14422
rect 7643 14413 7669 14469
rect 7725 14413 7751 14469
rect 7807 14413 7833 14469
rect 7889 14413 7915 14469
rect 7971 14413 7997 14422
rect 8053 14413 8079 14422
rect 8135 14413 8161 14469
rect 8217 14413 8243 14469
rect 8299 14413 8325 14469
rect 8381 14413 8407 14469
rect 8463 14413 8489 14469
rect 8545 14413 8571 14469
rect 8627 14413 8653 14469
rect 8709 14413 8735 14469
rect 8791 14413 8817 14469
rect 8873 14422 8881 14469
rect 8955 14422 8959 14469
rect 8873 14413 8899 14422
rect 8955 14413 8981 14422
rect 9037 14413 9063 14469
rect 9119 14413 9145 14469
rect 9201 14413 9227 14469
rect 9283 14413 9308 14469
rect 9364 14413 9389 14469
rect 9445 14413 9470 14469
rect 9526 14413 9551 14469
rect 9607 14413 9632 14469
rect 9688 14413 9713 14469
rect 9769 14422 9801 14469
rect 9853 14422 9879 14474
rect 9931 14422 10721 14474
rect 10773 14422 10799 14474
rect 10851 14422 11641 14474
rect 11693 14422 11719 14474
rect 11771 14422 12561 14474
rect 12613 14422 12639 14474
rect 12691 14422 14858 14474
rect 9769 14413 14858 14422
rect 4964 14409 14858 14413
rect 4964 14357 5201 14409
rect 5253 14357 5279 14409
rect 5331 14357 6121 14409
rect 6173 14357 6199 14409
rect 6251 14357 7041 14409
rect 7093 14357 7119 14409
rect 7171 14389 7961 14409
rect 8013 14389 8039 14409
rect 8091 14389 8881 14409
rect 8933 14389 8959 14409
rect 9011 14389 9801 14409
rect 7171 14357 7587 14389
rect 4964 14344 7587 14357
rect 4964 14292 5201 14344
rect 5253 14292 5279 14344
rect 5331 14292 6121 14344
rect 6173 14292 6199 14344
rect 6251 14292 7041 14344
rect 7093 14292 7119 14344
rect 7171 14333 7587 14344
rect 7643 14333 7669 14389
rect 7725 14333 7751 14389
rect 7807 14333 7833 14389
rect 7889 14333 7915 14389
rect 7971 14344 7997 14357
rect 8053 14344 8079 14357
rect 8135 14333 8161 14389
rect 8217 14333 8243 14389
rect 8299 14333 8325 14389
rect 8381 14333 8407 14389
rect 8463 14333 8489 14389
rect 8545 14333 8571 14389
rect 8627 14333 8653 14389
rect 8709 14333 8735 14389
rect 8791 14333 8817 14389
rect 8873 14357 8881 14389
rect 8955 14357 8959 14389
rect 8873 14344 8899 14357
rect 8955 14344 8981 14357
rect 8873 14333 8881 14344
rect 8955 14333 8959 14344
rect 9037 14333 9063 14389
rect 9119 14333 9145 14389
rect 9201 14333 9227 14389
rect 9283 14333 9308 14389
rect 9364 14333 9389 14389
rect 9445 14333 9470 14389
rect 9526 14333 9551 14389
rect 9607 14333 9632 14389
rect 9688 14333 9713 14389
rect 9769 14357 9801 14389
rect 9853 14357 9879 14409
rect 9931 14357 10721 14409
rect 10773 14357 10799 14409
rect 10851 14357 11641 14409
rect 11693 14357 11719 14409
rect 11771 14357 12561 14409
rect 12613 14357 12639 14409
rect 12691 14357 14858 14409
rect 9769 14344 14858 14357
rect 9769 14333 9801 14344
rect 7171 14309 7961 14333
rect 8013 14309 8039 14333
rect 8091 14309 8881 14333
rect 8933 14309 8959 14333
rect 9011 14309 9801 14333
rect 7171 14292 7587 14309
rect 4964 14279 7587 14292
rect 4964 14227 5201 14279
rect 5253 14227 5279 14279
rect 5331 14227 6121 14279
rect 6173 14227 6199 14279
rect 6251 14227 7041 14279
rect 7093 14227 7119 14279
rect 7171 14253 7587 14279
rect 7643 14253 7669 14309
rect 7725 14253 7751 14309
rect 7807 14253 7833 14309
rect 7889 14253 7915 14309
rect 7971 14279 7997 14292
rect 8053 14279 8079 14292
rect 8135 14253 8161 14309
rect 8217 14253 8243 14309
rect 8299 14253 8325 14309
rect 8381 14253 8407 14309
rect 8463 14253 8489 14309
rect 8545 14253 8571 14309
rect 8627 14253 8653 14309
rect 8709 14253 8735 14309
rect 8791 14253 8817 14309
rect 8873 14292 8881 14309
rect 8955 14292 8959 14309
rect 8873 14279 8899 14292
rect 8955 14279 8981 14292
rect 8873 14253 8881 14279
rect 8955 14253 8959 14279
rect 9037 14253 9063 14309
rect 9119 14253 9145 14309
rect 9201 14253 9227 14309
rect 9283 14253 9308 14309
rect 9364 14253 9389 14309
rect 9445 14253 9470 14309
rect 9526 14253 9551 14309
rect 9607 14253 9632 14309
rect 9688 14253 9713 14309
rect 9769 14292 9801 14309
rect 9853 14292 9879 14344
rect 9931 14292 10721 14344
rect 10773 14292 10799 14344
rect 10851 14292 11641 14344
rect 11693 14292 11719 14344
rect 11771 14292 12561 14344
rect 12613 14292 12639 14344
rect 12691 14292 14858 14344
rect 9769 14279 14858 14292
rect 9769 14253 9801 14279
rect 7171 14229 7961 14253
rect 8013 14229 8039 14253
rect 8091 14229 8881 14253
rect 8933 14229 8959 14253
rect 9011 14229 9801 14253
rect 7171 14227 7587 14229
rect 4964 14214 7587 14227
rect 4964 14162 5201 14214
rect 5253 14162 5279 14214
rect 5331 14162 6121 14214
rect 6173 14162 6199 14214
rect 6251 14162 7041 14214
rect 7093 14162 7119 14214
rect 7171 14173 7587 14214
rect 7643 14173 7669 14229
rect 7725 14173 7751 14229
rect 7807 14173 7833 14229
rect 7889 14173 7915 14229
rect 7971 14214 7997 14227
rect 8053 14214 8079 14227
rect 8135 14173 8161 14229
rect 8217 14173 8243 14229
rect 8299 14173 8325 14229
rect 8381 14173 8407 14229
rect 8463 14173 8489 14229
rect 8545 14173 8571 14229
rect 8627 14173 8653 14229
rect 8709 14173 8735 14229
rect 8791 14173 8817 14229
rect 8873 14227 8881 14229
rect 8955 14227 8959 14229
rect 8873 14214 8899 14227
rect 8955 14214 8981 14227
rect 8873 14173 8881 14214
rect 8955 14173 8959 14214
rect 9037 14173 9063 14229
rect 9119 14173 9145 14229
rect 9201 14173 9227 14229
rect 9283 14173 9308 14229
rect 9364 14173 9389 14229
rect 9445 14173 9470 14229
rect 9526 14173 9551 14229
rect 9607 14173 9632 14229
rect 9688 14173 9713 14229
rect 9769 14227 9801 14229
rect 9853 14227 9879 14279
rect 9931 14227 10721 14279
rect 10773 14227 10799 14279
rect 10851 14227 11641 14279
rect 11693 14227 11719 14279
rect 11771 14227 12561 14279
rect 12613 14227 12639 14279
rect 12691 14227 14858 14279
rect 9769 14214 14858 14227
rect 9769 14173 9801 14214
rect 7171 14162 7961 14173
rect 8013 14162 8039 14173
rect 8091 14162 8881 14173
rect 8933 14162 8959 14173
rect 9011 14162 9801 14173
rect 9853 14162 9879 14214
rect 9931 14162 10721 14214
rect 10773 14162 10799 14214
rect 10851 14162 11641 14214
rect 11693 14162 11719 14214
rect 11771 14162 12561 14214
rect 12613 14162 12639 14214
rect 12691 14162 14858 14214
rect 4964 14149 14858 14162
rect 4964 14097 5201 14149
rect 5253 14097 5279 14149
rect 5331 14097 6121 14149
rect 6173 14097 6199 14149
rect 6251 14097 7041 14149
rect 7093 14097 7119 14149
rect 7171 14097 7587 14149
rect 4964 14093 7587 14097
rect 7643 14093 7669 14149
rect 7725 14093 7751 14149
rect 7807 14093 7833 14149
rect 7889 14093 7915 14149
rect 7971 14093 7997 14097
rect 8053 14093 8079 14097
rect 8135 14093 8161 14149
rect 8217 14093 8243 14149
rect 8299 14093 8325 14149
rect 8381 14093 8407 14149
rect 8463 14093 8489 14149
rect 8545 14093 8571 14149
rect 8627 14093 8653 14149
rect 8709 14093 8735 14149
rect 8791 14093 8817 14149
rect 8873 14097 8881 14149
rect 8955 14097 8959 14149
rect 8873 14093 8899 14097
rect 8955 14093 8981 14097
rect 9037 14093 9063 14149
rect 9119 14093 9145 14149
rect 9201 14093 9227 14149
rect 9283 14093 9308 14149
rect 9364 14093 9389 14149
rect 9445 14093 9470 14149
rect 9526 14093 9551 14149
rect 9607 14093 9632 14149
rect 9688 14093 9713 14149
rect 9769 14097 9801 14149
rect 9853 14097 9879 14149
rect 9931 14097 10721 14149
rect 10773 14097 10799 14149
rect 10851 14097 11641 14149
rect 11693 14097 11719 14149
rect 11771 14097 12561 14149
rect 12613 14097 12639 14149
rect 12691 14097 14858 14149
rect 9769 14093 14858 14097
rect 4964 14091 14858 14093
tri 3433 13651 3470 13688 sw
rect 3361 13599 3367 13651
rect 3419 13599 3456 13651
rect 3508 13599 3514 13651
rect 187 13550 3230 13599
rect 187 13498 2233 13550
rect 2285 13498 2335 13550
rect 2387 13498 3230 13550
rect 187 13486 3230 13498
rect 187 13434 2233 13486
rect 2285 13434 2335 13486
rect 2387 13434 3230 13486
rect 187 13422 3230 13434
rect 187 13370 2233 13422
rect 2285 13370 2335 13422
rect 2387 13377 3230 13422
rect 2387 13370 2872 13377
rect 187 13358 2872 13370
rect 187 13306 2233 13358
rect 2285 13306 2335 13358
rect 2387 13325 2872 13358
rect 2924 13325 2940 13377
rect 2992 13325 3008 13377
rect 3060 13325 3230 13377
rect 2387 13312 3230 13325
rect 2387 13306 2872 13312
rect 187 13294 2872 13306
rect 187 13242 2233 13294
rect 2285 13242 2335 13294
rect 2387 13260 2872 13294
rect 2924 13260 2940 13312
rect 2992 13260 3008 13312
rect 3060 13296 3230 13312
tri 3230 13296 3533 13599 sw
tri 11501 13370 12222 14091 ne
rect 3060 13294 11342 13296
rect 3060 13290 5188 13294
rect 3060 13260 3792 13290
rect 2387 13247 3792 13260
rect 2387 13242 2872 13247
rect 187 13230 2872 13242
rect 187 13178 2233 13230
rect 2285 13178 2335 13230
rect 2387 13195 2872 13230
rect 2924 13195 2940 13247
rect 2992 13195 3008 13247
rect 3060 13238 3792 13247
rect 3844 13238 3860 13290
rect 3912 13238 3928 13290
rect 3980 13238 4712 13290
rect 4764 13238 4780 13290
rect 4832 13238 4848 13290
rect 4900 13238 5188 13290
rect 5244 13238 5270 13294
rect 5326 13238 5352 13294
rect 5408 13238 5434 13294
rect 5490 13238 5516 13294
rect 5572 13238 5598 13294
rect 5654 13290 5680 13294
rect 5736 13290 5762 13294
rect 5818 13290 5844 13294
rect 5752 13238 5762 13290
rect 5820 13238 5844 13290
rect 5900 13238 5926 13294
rect 5982 13238 6008 13294
rect 6064 13238 6090 13294
rect 6146 13238 6172 13294
rect 6228 13238 6254 13294
rect 6310 13238 6336 13294
rect 6392 13238 6418 13294
rect 6474 13238 6500 13294
rect 6556 13290 6582 13294
rect 6638 13290 6664 13294
rect 6720 13290 6746 13294
rect 6740 13238 6746 13290
rect 6802 13238 6828 13294
rect 6884 13238 6909 13294
rect 6965 13238 6990 13294
rect 7046 13238 7071 13294
rect 7127 13238 7152 13294
rect 7208 13238 7233 13294
rect 7289 13238 7314 13294
rect 7370 13290 11342 13294
rect 7370 13238 7472 13290
rect 7524 13238 7540 13290
rect 7592 13238 7608 13290
rect 7660 13238 8392 13290
rect 8444 13238 8460 13290
rect 8512 13238 8528 13290
rect 8580 13238 9312 13290
rect 9364 13238 9380 13290
rect 9432 13238 9448 13290
rect 9500 13238 10232 13290
rect 10284 13238 10300 13290
rect 10352 13238 10368 13290
rect 10420 13238 11152 13290
rect 11204 13238 11220 13290
rect 11272 13238 11288 13290
rect 11340 13238 11342 13290
rect 3060 13226 11342 13238
rect 3060 13195 3792 13226
rect 2387 13182 3792 13195
rect 2387 13178 2872 13182
rect 187 13166 2872 13178
rect 187 13114 2233 13166
rect 2285 13114 2335 13166
rect 2387 13130 2872 13166
rect 2924 13130 2940 13182
rect 2992 13130 3008 13182
rect 3060 13174 3792 13182
rect 3844 13174 3860 13226
rect 3912 13174 3928 13226
rect 3980 13174 4712 13226
rect 4764 13174 4780 13226
rect 4832 13174 4848 13226
rect 4900 13214 5632 13226
rect 5684 13214 5700 13226
rect 5752 13214 5768 13226
rect 5820 13214 6552 13226
rect 6604 13214 6620 13226
rect 6672 13214 6688 13226
rect 6740 13214 7472 13226
rect 4900 13174 5188 13214
rect 3060 13162 5188 13174
rect 3060 13130 3792 13162
rect 2387 13117 3792 13130
rect 2387 13114 2872 13117
rect 187 13102 2872 13114
rect 187 13050 2233 13102
rect 2285 13050 2335 13102
rect 2387 13065 2872 13102
rect 2924 13065 2940 13117
rect 2992 13065 3008 13117
rect 3060 13110 3792 13117
rect 3844 13110 3860 13162
rect 3912 13110 3928 13162
rect 3980 13110 4712 13162
rect 4764 13110 4780 13162
rect 4832 13110 4848 13162
rect 4900 13158 5188 13162
rect 5244 13158 5270 13214
rect 5326 13158 5352 13214
rect 5408 13158 5434 13214
rect 5490 13158 5516 13214
rect 5572 13158 5598 13214
rect 5752 13174 5762 13214
rect 5820 13174 5844 13214
rect 5654 13162 5680 13174
rect 5736 13162 5762 13174
rect 5818 13162 5844 13174
rect 5752 13158 5762 13162
rect 5820 13158 5844 13162
rect 5900 13158 5926 13214
rect 5982 13158 6008 13214
rect 6064 13158 6090 13214
rect 6146 13158 6172 13214
rect 6228 13158 6254 13214
rect 6310 13158 6336 13214
rect 6392 13158 6418 13214
rect 6474 13158 6500 13214
rect 6740 13174 6746 13214
rect 6556 13162 6582 13174
rect 6638 13162 6664 13174
rect 6720 13162 6746 13174
rect 6740 13158 6746 13162
rect 6802 13158 6828 13214
rect 6884 13158 6909 13214
rect 6965 13158 6990 13214
rect 7046 13158 7071 13214
rect 7127 13158 7152 13214
rect 7208 13158 7233 13214
rect 7289 13158 7314 13214
rect 7370 13174 7472 13214
rect 7524 13174 7540 13226
rect 7592 13174 7608 13226
rect 7660 13174 8392 13226
rect 8444 13174 8460 13226
rect 8512 13174 8528 13226
rect 8580 13174 9312 13226
rect 9364 13174 9380 13226
rect 9432 13174 9448 13226
rect 9500 13174 10232 13226
rect 10284 13174 10300 13226
rect 10352 13174 10368 13226
rect 10420 13174 11152 13226
rect 11204 13174 11220 13226
rect 11272 13174 11288 13226
rect 11340 13174 11342 13226
rect 7370 13162 11342 13174
rect 7370 13158 7472 13162
rect 4900 13134 5632 13158
rect 5684 13134 5700 13158
rect 5752 13134 5768 13158
rect 5820 13134 6552 13158
rect 6604 13134 6620 13158
rect 6672 13134 6688 13158
rect 6740 13134 7472 13158
rect 4900 13110 5188 13134
rect 3060 13098 5188 13110
rect 3060 13065 3792 13098
rect 2387 13052 3792 13065
rect 2387 13050 2872 13052
rect 187 13038 2872 13050
rect 187 12986 2233 13038
rect 2285 12986 2335 13038
rect 2387 13000 2872 13038
rect 2924 13000 2940 13052
rect 2992 13000 3008 13052
rect 3060 13046 3792 13052
rect 3844 13046 3860 13098
rect 3912 13046 3928 13098
rect 3980 13046 4712 13098
rect 4764 13046 4780 13098
rect 4832 13046 4848 13098
rect 4900 13078 5188 13098
rect 5244 13078 5270 13134
rect 5326 13078 5352 13134
rect 5408 13078 5434 13134
rect 5490 13078 5516 13134
rect 5572 13078 5598 13134
rect 5752 13110 5762 13134
rect 5820 13110 5844 13134
rect 5654 13098 5680 13110
rect 5736 13098 5762 13110
rect 5818 13098 5844 13110
rect 5752 13078 5762 13098
rect 5820 13078 5844 13098
rect 5900 13078 5926 13134
rect 5982 13078 6008 13134
rect 6064 13078 6090 13134
rect 6146 13078 6172 13134
rect 6228 13078 6254 13134
rect 6310 13078 6336 13134
rect 6392 13078 6418 13134
rect 6474 13078 6500 13134
rect 6740 13110 6746 13134
rect 6556 13098 6582 13110
rect 6638 13098 6664 13110
rect 6720 13098 6746 13110
rect 6740 13078 6746 13098
rect 6802 13078 6828 13134
rect 6884 13078 6909 13134
rect 6965 13078 6990 13134
rect 7046 13078 7071 13134
rect 7127 13078 7152 13134
rect 7208 13078 7233 13134
rect 7289 13078 7314 13134
rect 7370 13110 7472 13134
rect 7524 13110 7540 13162
rect 7592 13110 7608 13162
rect 7660 13110 8392 13162
rect 8444 13110 8460 13162
rect 8512 13110 8528 13162
rect 8580 13110 9312 13162
rect 9364 13110 9380 13162
rect 9432 13110 9448 13162
rect 9500 13110 10232 13162
rect 10284 13110 10300 13162
rect 10352 13110 10368 13162
rect 10420 13110 11152 13162
rect 11204 13110 11220 13162
rect 11272 13110 11288 13162
rect 11340 13110 11342 13162
rect 7370 13098 11342 13110
rect 7370 13078 7472 13098
rect 4900 13054 5632 13078
rect 5684 13054 5700 13078
rect 5752 13054 5768 13078
rect 5820 13054 6552 13078
rect 6604 13054 6620 13078
rect 6672 13054 6688 13078
rect 6740 13054 7472 13078
rect 4900 13046 5188 13054
rect 3060 13034 5188 13046
rect 3060 13000 3792 13034
rect 2387 12987 3792 13000
rect 2387 12986 2872 12987
rect 187 12974 2872 12986
rect 187 12922 2233 12974
rect 2285 12922 2335 12974
rect 2387 12935 2872 12974
rect 2924 12935 2940 12987
rect 2992 12935 3008 12987
rect 3060 12982 3792 12987
rect 3844 12982 3860 13034
rect 3912 12982 3928 13034
rect 3980 12982 4712 13034
rect 4764 12982 4780 13034
rect 4832 12982 4848 13034
rect 4900 12998 5188 13034
rect 5244 12998 5270 13054
rect 5326 12998 5352 13054
rect 5408 12998 5434 13054
rect 5490 12998 5516 13054
rect 5572 12998 5598 13054
rect 5752 13046 5762 13054
rect 5820 13046 5844 13054
rect 5654 13034 5680 13046
rect 5736 13034 5762 13046
rect 5818 13034 5844 13046
rect 5752 12998 5762 13034
rect 5820 12998 5844 13034
rect 5900 12998 5926 13054
rect 5982 12998 6008 13054
rect 6064 12998 6090 13054
rect 6146 12998 6172 13054
rect 6228 12998 6254 13054
rect 6310 12998 6336 13054
rect 6392 12998 6418 13054
rect 6474 12998 6500 13054
rect 6740 13046 6746 13054
rect 6556 13034 6582 13046
rect 6638 13034 6664 13046
rect 6720 13034 6746 13046
rect 6740 12998 6746 13034
rect 6802 12998 6828 13054
rect 6884 12998 6909 13054
rect 6965 12998 6990 13054
rect 7046 12998 7071 13054
rect 7127 12998 7152 13054
rect 7208 12998 7233 13054
rect 7289 12998 7314 13054
rect 7370 13046 7472 13054
rect 7524 13046 7540 13098
rect 7592 13046 7608 13098
rect 7660 13046 8392 13098
rect 8444 13046 8460 13098
rect 8512 13046 8528 13098
rect 8580 13046 9312 13098
rect 9364 13046 9380 13098
rect 9432 13046 9448 13098
rect 9500 13046 10232 13098
rect 10284 13046 10300 13098
rect 10352 13046 10368 13098
rect 10420 13046 11152 13098
rect 11204 13046 11220 13098
rect 11272 13046 11288 13098
rect 11340 13046 11342 13098
rect 7370 13034 11342 13046
rect 7370 12998 7472 13034
rect 4900 12982 5632 12998
rect 5684 12982 5700 12998
rect 5752 12982 5768 12998
rect 5820 12982 6552 12998
rect 6604 12982 6620 12998
rect 6672 12982 6688 12998
rect 6740 12982 7472 12998
rect 7524 12982 7540 13034
rect 7592 12982 7608 13034
rect 7660 12982 8392 13034
rect 8444 12982 8460 13034
rect 8512 12982 8528 13034
rect 8580 12982 9312 13034
rect 9364 12982 9380 13034
rect 9432 12982 9448 13034
rect 9500 12982 10232 13034
rect 10284 12982 10300 13034
rect 10352 12982 10368 13034
rect 10420 12982 11152 13034
rect 11204 12982 11220 13034
rect 11272 12982 11288 13034
rect 11340 12982 11342 13034
rect 3060 12974 11342 12982
rect 3060 12970 5188 12974
rect 3060 12935 3792 12970
rect 2387 12922 3792 12935
rect 187 12910 2872 12922
rect 187 12858 2233 12910
rect 2285 12858 2335 12910
rect 2387 12870 2872 12910
rect 2924 12870 2940 12922
rect 2992 12870 3008 12922
rect 3060 12918 3792 12922
rect 3844 12918 3860 12970
rect 3912 12918 3928 12970
rect 3980 12918 4712 12970
rect 4764 12918 4780 12970
rect 4832 12918 4848 12970
rect 4900 12918 5188 12970
rect 5244 12918 5270 12974
rect 5326 12918 5352 12974
rect 5408 12918 5434 12974
rect 5490 12918 5516 12974
rect 5572 12918 5598 12974
rect 5654 12970 5680 12974
rect 5736 12970 5762 12974
rect 5818 12970 5844 12974
rect 5752 12918 5762 12970
rect 5820 12918 5844 12970
rect 5900 12918 5926 12974
rect 5982 12918 6008 12974
rect 6064 12918 6090 12974
rect 6146 12918 6172 12974
rect 6228 12918 6254 12974
rect 6310 12918 6336 12974
rect 6392 12918 6418 12974
rect 6474 12918 6500 12974
rect 6556 12970 6582 12974
rect 6638 12970 6664 12974
rect 6720 12970 6746 12974
rect 6740 12918 6746 12970
rect 6802 12918 6828 12974
rect 6884 12918 6909 12974
rect 6965 12918 6990 12974
rect 7046 12918 7071 12974
rect 7127 12918 7152 12974
rect 7208 12918 7233 12974
rect 7289 12918 7314 12974
rect 7370 12970 11342 12974
rect 7370 12918 7472 12970
rect 7524 12918 7540 12970
rect 7592 12918 7608 12970
rect 7660 12918 8392 12970
rect 8444 12918 8460 12970
rect 8512 12918 8528 12970
rect 8580 12918 9312 12970
rect 9364 12918 9380 12970
rect 9432 12918 9448 12970
rect 9500 12918 10232 12970
rect 10284 12918 10300 12970
rect 10352 12918 10368 12970
rect 10420 12918 11152 12970
rect 11204 12918 11220 12970
rect 11272 12918 11288 12970
rect 11340 12918 11342 12970
rect 3060 12906 11342 12918
rect 3060 12870 3792 12906
rect 2387 12858 3792 12870
rect 187 12857 3792 12858
rect 187 12846 2872 12857
rect 187 12794 2233 12846
rect 2285 12794 2335 12846
rect 2387 12805 2872 12846
rect 2924 12805 2940 12857
rect 2992 12805 3008 12857
rect 3060 12854 3792 12857
rect 3844 12854 3860 12906
rect 3912 12854 3928 12906
rect 3980 12854 4712 12906
rect 4764 12854 4780 12906
rect 4832 12854 4848 12906
rect 4900 12894 5632 12906
rect 5684 12894 5700 12906
rect 5752 12894 5768 12906
rect 5820 12894 6552 12906
rect 6604 12894 6620 12906
rect 6672 12894 6688 12906
rect 6740 12894 7472 12906
rect 4900 12854 5188 12894
rect 3060 12842 5188 12854
rect 3060 12805 3792 12842
rect 2387 12794 3792 12805
rect 187 12792 3792 12794
rect 187 12782 2872 12792
rect 187 12730 2233 12782
rect 2285 12730 2335 12782
rect 2387 12740 2872 12782
rect 2924 12740 2940 12792
rect 2992 12740 3008 12792
rect 3060 12790 3792 12792
rect 3844 12790 3860 12842
rect 3912 12790 3928 12842
rect 3980 12790 4712 12842
rect 4764 12790 4780 12842
rect 4832 12790 4848 12842
rect 4900 12838 5188 12842
rect 5244 12838 5270 12894
rect 5326 12838 5352 12894
rect 5408 12838 5434 12894
rect 5490 12838 5516 12894
rect 5572 12838 5598 12894
rect 5752 12854 5762 12894
rect 5820 12854 5844 12894
rect 5654 12842 5680 12854
rect 5736 12842 5762 12854
rect 5818 12842 5844 12854
rect 5752 12838 5762 12842
rect 5820 12838 5844 12842
rect 5900 12838 5926 12894
rect 5982 12838 6008 12894
rect 6064 12838 6090 12894
rect 6146 12838 6172 12894
rect 6228 12838 6254 12894
rect 6310 12838 6336 12894
rect 6392 12838 6418 12894
rect 6474 12838 6500 12894
rect 6740 12854 6746 12894
rect 6556 12842 6582 12854
rect 6638 12842 6664 12854
rect 6720 12842 6746 12854
rect 6740 12838 6746 12842
rect 6802 12838 6828 12894
rect 6884 12838 6909 12894
rect 6965 12838 6990 12894
rect 7046 12838 7071 12894
rect 7127 12838 7152 12894
rect 7208 12838 7233 12894
rect 7289 12838 7314 12894
rect 7370 12854 7472 12894
rect 7524 12854 7540 12906
rect 7592 12854 7608 12906
rect 7660 12854 8392 12906
rect 8444 12854 8460 12906
rect 8512 12854 8528 12906
rect 8580 12854 9312 12906
rect 9364 12854 9380 12906
rect 9432 12854 9448 12906
rect 9500 12854 10232 12906
rect 10284 12854 10300 12906
rect 10352 12854 10368 12906
rect 10420 12854 11152 12906
rect 11204 12854 11220 12906
rect 11272 12854 11288 12906
rect 11340 12854 11342 12906
rect 7370 12842 11342 12854
rect 7370 12838 7472 12842
rect 4900 12814 5632 12838
rect 5684 12814 5700 12838
rect 5752 12814 5768 12838
rect 5820 12814 6552 12838
rect 6604 12814 6620 12838
rect 6672 12814 6688 12838
rect 6740 12814 7472 12838
rect 4900 12790 5188 12814
rect 3060 12778 5188 12790
rect 3060 12740 3792 12778
rect 2387 12730 3792 12740
rect 187 12727 3792 12730
rect 187 12718 2872 12727
rect 187 12666 2233 12718
rect 2285 12666 2335 12718
rect 2387 12675 2872 12718
rect 2924 12675 2940 12727
rect 2992 12675 3008 12727
rect 3060 12726 3792 12727
rect 3844 12726 3860 12778
rect 3912 12726 3928 12778
rect 3980 12726 4712 12778
rect 4764 12726 4780 12778
rect 4832 12726 4848 12778
rect 4900 12758 5188 12778
rect 5244 12758 5270 12814
rect 5326 12758 5352 12814
rect 5408 12758 5434 12814
rect 5490 12758 5516 12814
rect 5572 12758 5598 12814
rect 5752 12790 5762 12814
rect 5820 12790 5844 12814
rect 5654 12778 5680 12790
rect 5736 12778 5762 12790
rect 5818 12778 5844 12790
rect 5752 12758 5762 12778
rect 5820 12758 5844 12778
rect 5900 12758 5926 12814
rect 5982 12758 6008 12814
rect 6064 12758 6090 12814
rect 6146 12758 6172 12814
rect 6228 12758 6254 12814
rect 6310 12758 6336 12814
rect 6392 12758 6418 12814
rect 6474 12758 6500 12814
rect 6740 12790 6746 12814
rect 6556 12778 6582 12790
rect 6638 12778 6664 12790
rect 6720 12778 6746 12790
rect 6740 12758 6746 12778
rect 6802 12758 6828 12814
rect 6884 12758 6909 12814
rect 6965 12758 6990 12814
rect 7046 12758 7071 12814
rect 7127 12758 7152 12814
rect 7208 12758 7233 12814
rect 7289 12758 7314 12814
rect 7370 12790 7472 12814
rect 7524 12790 7540 12842
rect 7592 12790 7608 12842
rect 7660 12790 8392 12842
rect 8444 12790 8460 12842
rect 8512 12790 8528 12842
rect 8580 12790 9312 12842
rect 9364 12790 9380 12842
rect 9432 12790 9448 12842
rect 9500 12790 10232 12842
rect 10284 12790 10300 12842
rect 10352 12790 10368 12842
rect 10420 12790 11152 12842
rect 11204 12790 11220 12842
rect 11272 12790 11288 12842
rect 11340 12790 11342 12842
rect 7370 12778 11342 12790
rect 7370 12758 7472 12778
rect 4900 12734 5632 12758
rect 5684 12734 5700 12758
rect 5752 12734 5768 12758
rect 5820 12734 6552 12758
rect 6604 12734 6620 12758
rect 6672 12734 6688 12758
rect 6740 12734 7472 12758
rect 4900 12726 5188 12734
rect 3060 12714 5188 12726
rect 3060 12675 3792 12714
rect 2387 12666 3792 12675
rect 187 12662 3792 12666
rect 3844 12662 3860 12714
rect 3912 12662 3928 12714
rect 3980 12662 4712 12714
rect 4764 12662 4780 12714
rect 4832 12662 4848 12714
rect 4900 12678 5188 12714
rect 5244 12678 5270 12734
rect 5326 12678 5352 12734
rect 5408 12678 5434 12734
rect 5490 12678 5516 12734
rect 5572 12678 5598 12734
rect 5752 12726 5762 12734
rect 5820 12726 5844 12734
rect 5654 12714 5680 12726
rect 5736 12714 5762 12726
rect 5818 12714 5844 12726
rect 5752 12678 5762 12714
rect 5820 12678 5844 12714
rect 5900 12678 5926 12734
rect 5982 12678 6008 12734
rect 6064 12678 6090 12734
rect 6146 12678 6172 12734
rect 6228 12678 6254 12734
rect 6310 12678 6336 12734
rect 6392 12678 6418 12734
rect 6474 12678 6500 12734
rect 6740 12726 6746 12734
rect 6556 12714 6582 12726
rect 6638 12714 6664 12726
rect 6720 12714 6746 12726
rect 6740 12678 6746 12714
rect 6802 12678 6828 12734
rect 6884 12678 6909 12734
rect 6965 12678 6990 12734
rect 7046 12678 7071 12734
rect 7127 12678 7152 12734
rect 7208 12678 7233 12734
rect 7289 12678 7314 12734
rect 7370 12726 7472 12734
rect 7524 12726 7540 12778
rect 7592 12726 7608 12778
rect 7660 12726 8392 12778
rect 8444 12726 8460 12778
rect 8512 12726 8528 12778
rect 8580 12726 9312 12778
rect 9364 12726 9380 12778
rect 9432 12726 9448 12778
rect 9500 12726 10232 12778
rect 10284 12726 10300 12778
rect 10352 12726 10368 12778
rect 10420 12726 11152 12778
rect 11204 12726 11220 12778
rect 11272 12726 11288 12778
rect 11340 12726 11342 12778
rect 7370 12714 11342 12726
rect 7370 12678 7472 12714
rect 4900 12662 5632 12678
rect 5684 12662 5700 12678
rect 5752 12662 5768 12678
rect 5820 12662 6552 12678
rect 6604 12662 6620 12678
rect 6672 12662 6688 12678
rect 6740 12662 7472 12678
rect 7524 12662 7540 12714
rect 7592 12662 7608 12714
rect 7660 12662 8392 12714
rect 8444 12662 8460 12714
rect 8512 12662 8528 12714
rect 8580 12662 9312 12714
rect 9364 12662 9380 12714
rect 9432 12662 9448 12714
rect 9500 12662 10232 12714
rect 10284 12662 10300 12714
rect 10352 12662 10368 12714
rect 10420 12662 11152 12714
rect 11204 12662 11220 12714
rect 11272 12662 11288 12714
rect 11340 12662 11342 12714
rect 187 12654 2872 12662
rect 187 12602 2233 12654
rect 2285 12602 2335 12654
rect 2387 12610 2872 12654
rect 2924 12610 2940 12662
rect 2992 12610 3008 12662
rect 3060 12654 11342 12662
rect 3060 12650 5188 12654
rect 3060 12610 3792 12650
rect 2387 12602 3792 12610
rect 187 12598 3792 12602
rect 3844 12598 3860 12650
rect 3912 12598 3928 12650
rect 3980 12598 4712 12650
rect 4764 12598 4780 12650
rect 4832 12598 4848 12650
rect 4900 12598 5188 12650
rect 5244 12598 5270 12654
rect 5326 12598 5352 12654
rect 5408 12598 5434 12654
rect 5490 12598 5516 12654
rect 5572 12598 5598 12654
rect 5654 12650 5680 12654
rect 5736 12650 5762 12654
rect 5818 12650 5844 12654
rect 5752 12598 5762 12650
rect 5820 12598 5844 12650
rect 5900 12598 5926 12654
rect 5982 12598 6008 12654
rect 6064 12598 6090 12654
rect 6146 12598 6172 12654
rect 6228 12598 6254 12654
rect 6310 12598 6336 12654
rect 6392 12598 6418 12654
rect 6474 12598 6500 12654
rect 6556 12650 6582 12654
rect 6638 12650 6664 12654
rect 6720 12650 6746 12654
rect 6740 12598 6746 12650
rect 6802 12598 6828 12654
rect 6884 12598 6909 12654
rect 6965 12598 6990 12654
rect 7046 12598 7071 12654
rect 7127 12598 7152 12654
rect 7208 12598 7233 12654
rect 7289 12598 7314 12654
rect 7370 12650 11342 12654
rect 7370 12598 7472 12650
rect 7524 12598 7540 12650
rect 7592 12598 7608 12650
rect 7660 12598 8392 12650
rect 8444 12598 8460 12650
rect 8512 12598 8528 12650
rect 8580 12598 9312 12650
rect 9364 12598 9380 12650
rect 9432 12598 9448 12650
rect 9500 12598 10232 12650
rect 10284 12598 10300 12650
rect 10352 12598 10368 12650
rect 10420 12598 11152 12650
rect 11204 12598 11220 12650
rect 11272 12598 11288 12650
rect 11340 12598 11342 12650
rect 187 12597 11342 12598
rect 187 12590 2872 12597
rect 187 12538 2233 12590
rect 2285 12538 2335 12590
rect 2387 12545 2872 12590
rect 2924 12545 2940 12597
rect 2992 12545 3008 12597
rect 3060 12586 11342 12597
rect 3060 12545 3792 12586
rect 2387 12538 3792 12545
rect 187 12534 3792 12538
rect 3844 12534 3860 12586
rect 3912 12534 3928 12586
rect 3980 12534 4712 12586
rect 4764 12534 4780 12586
rect 4832 12534 4848 12586
rect 4900 12574 5632 12586
rect 5684 12574 5700 12586
rect 5752 12574 5768 12586
rect 5820 12574 6552 12586
rect 6604 12574 6620 12586
rect 6672 12574 6688 12586
rect 6740 12574 7472 12586
rect 4900 12534 5188 12574
rect 187 12532 5188 12534
rect 187 12526 2872 12532
rect 187 12474 2233 12526
rect 2285 12474 2335 12526
rect 2387 12480 2872 12526
rect 2924 12480 2940 12532
rect 2992 12480 3008 12532
rect 3060 12522 5188 12532
rect 3060 12480 3792 12522
rect 2387 12474 3792 12480
rect 187 12470 3792 12474
rect 3844 12470 3860 12522
rect 3912 12470 3928 12522
rect 3980 12470 4712 12522
rect 4764 12470 4780 12522
rect 4832 12470 4848 12522
rect 4900 12518 5188 12522
rect 5244 12518 5270 12574
rect 5326 12518 5352 12574
rect 5408 12518 5434 12574
rect 5490 12518 5516 12574
rect 5572 12518 5598 12574
rect 5752 12534 5762 12574
rect 5820 12534 5844 12574
rect 5654 12522 5680 12534
rect 5736 12522 5762 12534
rect 5818 12522 5844 12534
rect 5752 12518 5762 12522
rect 5820 12518 5844 12522
rect 5900 12518 5926 12574
rect 5982 12518 6008 12574
rect 6064 12518 6090 12574
rect 6146 12518 6172 12574
rect 6228 12518 6254 12574
rect 6310 12518 6336 12574
rect 6392 12518 6418 12574
rect 6474 12518 6500 12574
rect 6740 12534 6746 12574
rect 6556 12522 6582 12534
rect 6638 12522 6664 12534
rect 6720 12522 6746 12534
rect 6740 12518 6746 12522
rect 6802 12518 6828 12574
rect 6884 12518 6909 12574
rect 6965 12518 6990 12574
rect 7046 12518 7071 12574
rect 7127 12518 7152 12574
rect 7208 12518 7233 12574
rect 7289 12518 7314 12574
rect 7370 12534 7472 12574
rect 7524 12534 7540 12586
rect 7592 12534 7608 12586
rect 7660 12534 8392 12586
rect 8444 12534 8460 12586
rect 8512 12534 8528 12586
rect 8580 12534 9312 12586
rect 9364 12534 9380 12586
rect 9432 12534 9448 12586
rect 9500 12534 10232 12586
rect 10284 12534 10300 12586
rect 10352 12534 10368 12586
rect 10420 12534 11152 12586
rect 11204 12534 11220 12586
rect 11272 12534 11288 12586
rect 11340 12534 11342 12586
rect 7370 12522 11342 12534
rect 7370 12518 7472 12522
rect 4900 12494 5632 12518
rect 5684 12494 5700 12518
rect 5752 12494 5768 12518
rect 5820 12494 6552 12518
rect 6604 12494 6620 12518
rect 6672 12494 6688 12518
rect 6740 12494 7472 12518
rect 4900 12470 5188 12494
rect 187 12467 5188 12470
rect 187 12462 2872 12467
rect 187 12410 2233 12462
rect 2285 12410 2335 12462
rect 2387 12415 2872 12462
rect 2924 12415 2940 12467
rect 2992 12415 3008 12467
rect 3060 12458 5188 12467
rect 3060 12415 3792 12458
rect 2387 12410 3792 12415
rect 187 12406 3792 12410
rect 3844 12406 3860 12458
rect 3912 12406 3928 12458
rect 3980 12406 4712 12458
rect 4764 12406 4780 12458
rect 4832 12406 4848 12458
rect 4900 12438 5188 12458
rect 5244 12438 5270 12494
rect 5326 12438 5352 12494
rect 5408 12438 5434 12494
rect 5490 12438 5516 12494
rect 5572 12438 5598 12494
rect 5752 12470 5762 12494
rect 5820 12470 5844 12494
rect 5654 12458 5680 12470
rect 5736 12458 5762 12470
rect 5818 12458 5844 12470
rect 5752 12438 5762 12458
rect 5820 12438 5844 12458
rect 5900 12438 5926 12494
rect 5982 12438 6008 12494
rect 6064 12438 6090 12494
rect 6146 12438 6172 12494
rect 6228 12438 6254 12494
rect 6310 12438 6336 12494
rect 6392 12438 6418 12494
rect 6474 12438 6500 12494
rect 6740 12470 6746 12494
rect 6556 12458 6582 12470
rect 6638 12458 6664 12470
rect 6720 12458 6746 12470
rect 6740 12438 6746 12458
rect 6802 12438 6828 12494
rect 6884 12438 6909 12494
rect 6965 12438 6990 12494
rect 7046 12438 7071 12494
rect 7127 12438 7152 12494
rect 7208 12438 7233 12494
rect 7289 12438 7314 12494
rect 7370 12470 7472 12494
rect 7524 12470 7540 12522
rect 7592 12470 7608 12522
rect 7660 12470 8392 12522
rect 8444 12470 8460 12522
rect 8512 12470 8528 12522
rect 8580 12470 9312 12522
rect 9364 12470 9380 12522
rect 9432 12470 9448 12522
rect 9500 12470 10232 12522
rect 10284 12470 10300 12522
rect 10352 12470 10368 12522
rect 10420 12470 11152 12522
rect 11204 12470 11220 12522
rect 11272 12470 11288 12522
rect 11340 12470 11342 12522
rect 7370 12458 11342 12470
rect 7370 12438 7472 12458
rect 4900 12414 5632 12438
rect 5684 12414 5700 12438
rect 5752 12414 5768 12438
rect 5820 12414 6552 12438
rect 6604 12414 6620 12438
rect 6672 12414 6688 12438
rect 6740 12414 7472 12438
rect 4900 12406 5188 12414
rect 187 12402 5188 12406
rect 187 12398 2872 12402
rect 187 12346 2233 12398
rect 2285 12346 2335 12398
rect 2387 12350 2872 12398
rect 2924 12350 2940 12402
rect 2992 12350 3008 12402
rect 3060 12394 5188 12402
rect 3060 12350 3792 12394
rect 2387 12346 3792 12350
rect 187 12342 3792 12346
rect 3844 12342 3860 12394
rect 3912 12342 3928 12394
rect 3980 12342 4712 12394
rect 4764 12342 4780 12394
rect 4832 12342 4848 12394
rect 4900 12358 5188 12394
rect 5244 12358 5270 12414
rect 5326 12358 5352 12414
rect 5408 12358 5434 12414
rect 5490 12358 5516 12414
rect 5572 12358 5598 12414
rect 5752 12406 5762 12414
rect 5820 12406 5844 12414
rect 5654 12394 5680 12406
rect 5736 12394 5762 12406
rect 5818 12394 5844 12406
rect 5752 12358 5762 12394
rect 5820 12358 5844 12394
rect 5900 12358 5926 12414
rect 5982 12358 6008 12414
rect 6064 12358 6090 12414
rect 6146 12358 6172 12414
rect 6228 12358 6254 12414
rect 6310 12358 6336 12414
rect 6392 12358 6418 12414
rect 6474 12358 6500 12414
rect 6740 12406 6746 12414
rect 6556 12394 6582 12406
rect 6638 12394 6664 12406
rect 6720 12394 6746 12406
rect 6740 12358 6746 12394
rect 6802 12358 6828 12414
rect 6884 12358 6909 12414
rect 6965 12358 6990 12414
rect 7046 12358 7071 12414
rect 7127 12358 7152 12414
rect 7208 12358 7233 12414
rect 7289 12358 7314 12414
rect 7370 12406 7472 12414
rect 7524 12406 7540 12458
rect 7592 12406 7608 12458
rect 7660 12406 8392 12458
rect 8444 12406 8460 12458
rect 8512 12406 8528 12458
rect 8580 12406 9312 12458
rect 9364 12406 9380 12458
rect 9432 12406 9448 12458
rect 9500 12406 10232 12458
rect 10284 12406 10300 12458
rect 10352 12406 10368 12458
rect 10420 12406 11152 12458
rect 11204 12406 11220 12458
rect 11272 12406 11288 12458
rect 11340 12406 11342 12458
rect 7370 12394 11342 12406
rect 7370 12358 7472 12394
rect 4900 12342 5632 12358
rect 5684 12342 5700 12358
rect 5752 12342 5768 12358
rect 5820 12342 6552 12358
rect 6604 12342 6620 12358
rect 6672 12342 6688 12358
rect 6740 12342 7472 12358
rect 7524 12342 7540 12394
rect 7592 12342 7608 12394
rect 7660 12342 8392 12394
rect 8444 12342 8460 12394
rect 8512 12342 8528 12394
rect 8580 12342 9312 12394
rect 9364 12342 9380 12394
rect 9432 12342 9448 12394
rect 9500 12342 10232 12394
rect 10284 12342 10300 12394
rect 10352 12342 10368 12394
rect 10420 12342 11152 12394
rect 11204 12342 11220 12394
rect 11272 12342 11288 12394
rect 11340 12342 11342 12394
rect 187 12337 11342 12342
rect 187 12334 2872 12337
rect 187 12282 2233 12334
rect 2285 12282 2335 12334
rect 2387 12285 2872 12334
rect 2924 12285 2940 12337
rect 2992 12285 3008 12337
rect 3060 12334 11342 12337
rect 3060 12329 5188 12334
rect 3060 12285 3792 12329
rect 2387 12282 3792 12285
rect 187 12277 3792 12282
rect 3844 12277 3860 12329
rect 3912 12277 3928 12329
rect 3980 12277 4712 12329
rect 4764 12277 4780 12329
rect 4832 12277 4848 12329
rect 4900 12278 5188 12329
rect 5244 12278 5270 12334
rect 5326 12278 5352 12334
rect 5408 12278 5434 12334
rect 5490 12278 5516 12334
rect 5572 12278 5598 12334
rect 5654 12329 5680 12334
rect 5736 12329 5762 12334
rect 5818 12329 5844 12334
rect 5752 12278 5762 12329
rect 5820 12278 5844 12329
rect 5900 12278 5926 12334
rect 5982 12278 6008 12334
rect 6064 12278 6090 12334
rect 6146 12278 6172 12334
rect 6228 12278 6254 12334
rect 6310 12278 6336 12334
rect 6392 12278 6418 12334
rect 6474 12278 6500 12334
rect 6556 12329 6582 12334
rect 6638 12329 6664 12334
rect 6720 12329 6746 12334
rect 6740 12278 6746 12329
rect 6802 12278 6828 12334
rect 6884 12278 6909 12334
rect 6965 12278 6990 12334
rect 7046 12278 7071 12334
rect 7127 12278 7152 12334
rect 7208 12278 7233 12334
rect 7289 12278 7314 12334
rect 7370 12329 11342 12334
rect 7370 12278 7472 12329
rect 4900 12277 5632 12278
rect 5684 12277 5700 12278
rect 5752 12277 5768 12278
rect 5820 12277 6552 12278
rect 6604 12277 6620 12278
rect 6672 12277 6688 12278
rect 6740 12277 7472 12278
rect 7524 12277 7540 12329
rect 7592 12277 7608 12329
rect 7660 12277 8392 12329
rect 8444 12277 8460 12329
rect 8512 12277 8528 12329
rect 8580 12277 9312 12329
rect 9364 12277 9380 12329
rect 9432 12277 9448 12329
rect 9500 12277 10232 12329
rect 10284 12277 10300 12329
rect 10352 12277 10368 12329
rect 10420 12277 11152 12329
rect 11204 12277 11220 12329
rect 11272 12277 11288 12329
rect 11340 12277 11342 12329
rect 187 12272 11342 12277
rect 187 12270 2872 12272
rect 187 12218 2233 12270
rect 2285 12218 2335 12270
rect 2387 12220 2872 12270
rect 2924 12220 2940 12272
rect 2992 12220 3008 12272
rect 3060 12264 11342 12272
rect 3060 12220 3792 12264
rect 2387 12218 3792 12220
rect 187 12212 3792 12218
rect 3844 12212 3860 12264
rect 3912 12212 3928 12264
rect 3980 12212 4712 12264
rect 4764 12212 4780 12264
rect 4832 12212 4848 12264
rect 4900 12254 5632 12264
rect 5684 12254 5700 12264
rect 5752 12254 5768 12264
rect 5820 12254 6552 12264
rect 6604 12254 6620 12264
rect 6672 12254 6688 12264
rect 6740 12254 7472 12264
rect 4900 12212 5188 12254
rect 187 12207 5188 12212
rect 187 12206 2872 12207
rect 187 12154 2233 12206
rect 2285 12154 2335 12206
rect 2387 12155 2872 12206
rect 2924 12155 2940 12207
rect 2992 12155 3008 12207
rect 3060 12199 5188 12207
rect 3060 12155 3792 12199
rect 2387 12154 3792 12155
rect 187 12147 3792 12154
rect 3844 12147 3860 12199
rect 3912 12147 3928 12199
rect 3980 12147 4712 12199
rect 4764 12147 4780 12199
rect 4832 12147 4848 12199
rect 4900 12198 5188 12199
rect 5244 12198 5270 12254
rect 5326 12198 5352 12254
rect 5408 12198 5434 12254
rect 5490 12198 5516 12254
rect 5572 12198 5598 12254
rect 5752 12212 5762 12254
rect 5820 12212 5844 12254
rect 5654 12199 5680 12212
rect 5736 12199 5762 12212
rect 5818 12199 5844 12212
rect 5752 12198 5762 12199
rect 5820 12198 5844 12199
rect 5900 12198 5926 12254
rect 5982 12198 6008 12254
rect 6064 12198 6090 12254
rect 6146 12198 6172 12254
rect 6228 12198 6254 12254
rect 6310 12198 6336 12254
rect 6392 12198 6418 12254
rect 6474 12198 6500 12254
rect 6740 12212 6746 12254
rect 6556 12199 6582 12212
rect 6638 12199 6664 12212
rect 6720 12199 6746 12212
rect 6740 12198 6746 12199
rect 6802 12198 6828 12254
rect 6884 12198 6909 12254
rect 6965 12198 6990 12254
rect 7046 12198 7071 12254
rect 7127 12198 7152 12254
rect 7208 12198 7233 12254
rect 7289 12198 7314 12254
rect 7370 12212 7472 12254
rect 7524 12212 7540 12264
rect 7592 12212 7608 12264
rect 7660 12212 8392 12264
rect 8444 12212 8460 12264
rect 8512 12212 8528 12264
rect 8580 12212 9312 12264
rect 9364 12212 9380 12264
rect 9432 12212 9448 12264
rect 9500 12212 10232 12264
rect 10284 12212 10300 12264
rect 10352 12212 10368 12264
rect 10420 12212 11152 12264
rect 11204 12212 11220 12264
rect 11272 12212 11288 12264
rect 11340 12212 11342 12264
rect 7370 12199 11342 12212
rect 7370 12198 7472 12199
rect 4900 12174 5632 12198
rect 5684 12174 5700 12198
rect 5752 12174 5768 12198
rect 5820 12174 6552 12198
rect 6604 12174 6620 12198
rect 6672 12174 6688 12198
rect 6740 12174 7472 12198
rect 4900 12147 5188 12174
rect 187 12142 5188 12147
rect 187 12090 2233 12142
rect 2285 12090 2335 12142
rect 2387 12090 2872 12142
rect 2924 12090 2940 12142
rect 2992 12090 3008 12142
rect 3060 12134 5188 12142
rect 3060 12090 3792 12134
rect 187 12082 3792 12090
rect 3844 12082 3860 12134
rect 3912 12082 3928 12134
rect 3980 12082 4712 12134
rect 4764 12082 4780 12134
rect 4832 12082 4848 12134
rect 4900 12118 5188 12134
rect 5244 12118 5270 12174
rect 5326 12118 5352 12174
rect 5408 12118 5434 12174
rect 5490 12118 5516 12174
rect 5572 12118 5598 12174
rect 5752 12147 5762 12174
rect 5820 12147 5844 12174
rect 5654 12134 5680 12147
rect 5736 12134 5762 12147
rect 5818 12134 5844 12147
rect 5752 12118 5762 12134
rect 5820 12118 5844 12134
rect 5900 12118 5926 12174
rect 5982 12118 6008 12174
rect 6064 12118 6090 12174
rect 6146 12118 6172 12174
rect 6228 12118 6254 12174
rect 6310 12118 6336 12174
rect 6392 12118 6418 12174
rect 6474 12118 6500 12174
rect 6740 12147 6746 12174
rect 6556 12134 6582 12147
rect 6638 12134 6664 12147
rect 6720 12134 6746 12147
rect 6740 12118 6746 12134
rect 6802 12118 6828 12174
rect 6884 12118 6909 12174
rect 6965 12118 6990 12174
rect 7046 12118 7071 12174
rect 7127 12118 7152 12174
rect 7208 12118 7233 12174
rect 7289 12118 7314 12174
rect 7370 12147 7472 12174
rect 7524 12147 7540 12199
rect 7592 12147 7608 12199
rect 7660 12147 8392 12199
rect 8444 12147 8460 12199
rect 8512 12147 8528 12199
rect 8580 12147 9312 12199
rect 9364 12147 9380 12199
rect 9432 12147 9448 12199
rect 9500 12147 10232 12199
rect 10284 12147 10300 12199
rect 10352 12147 10368 12199
rect 10420 12147 11152 12199
rect 11204 12147 11220 12199
rect 11272 12147 11288 12199
rect 11340 12147 11342 12199
rect 7370 12134 11342 12147
rect 7370 12118 7472 12134
rect 4900 12094 5632 12118
rect 5684 12094 5700 12118
rect 5752 12094 5768 12118
rect 5820 12094 6552 12118
rect 6604 12094 6620 12118
rect 6672 12094 6688 12118
rect 6740 12094 7472 12118
rect 4900 12082 5188 12094
rect 187 12078 5188 12082
rect 187 12026 2233 12078
rect 2285 12026 2335 12078
rect 2387 12076 5188 12078
rect 2387 12026 2872 12076
rect 187 12024 2872 12026
rect 2924 12024 2940 12076
rect 2992 12024 3008 12076
rect 3060 12069 5188 12076
rect 3060 12024 3792 12069
rect 187 12017 3792 12024
rect 3844 12017 3860 12069
rect 3912 12017 3928 12069
rect 3980 12017 4712 12069
rect 4764 12017 4780 12069
rect 4832 12017 4848 12069
rect 4900 12038 5188 12069
rect 5244 12038 5270 12094
rect 5326 12038 5352 12094
rect 5408 12038 5434 12094
rect 5490 12038 5516 12094
rect 5572 12038 5598 12094
rect 5752 12082 5762 12094
rect 5820 12082 5844 12094
rect 5654 12069 5680 12082
rect 5736 12069 5762 12082
rect 5818 12069 5844 12082
rect 5752 12038 5762 12069
rect 5820 12038 5844 12069
rect 5900 12038 5926 12094
rect 5982 12038 6008 12094
rect 6064 12038 6090 12094
rect 6146 12038 6172 12094
rect 6228 12038 6254 12094
rect 6310 12038 6336 12094
rect 6392 12038 6418 12094
rect 6474 12038 6500 12094
rect 6740 12082 6746 12094
rect 6556 12069 6582 12082
rect 6638 12069 6664 12082
rect 6720 12069 6746 12082
rect 6740 12038 6746 12069
rect 6802 12038 6828 12094
rect 6884 12038 6909 12094
rect 6965 12038 6990 12094
rect 7046 12038 7071 12094
rect 7127 12038 7152 12094
rect 7208 12038 7233 12094
rect 7289 12038 7314 12094
rect 7370 12082 7472 12094
rect 7524 12082 7540 12134
rect 7592 12082 7608 12134
rect 7660 12082 8392 12134
rect 8444 12082 8460 12134
rect 8512 12082 8528 12134
rect 8580 12082 9312 12134
rect 9364 12082 9380 12134
rect 9432 12082 9448 12134
rect 9500 12082 10232 12134
rect 10284 12082 10300 12134
rect 10352 12082 10368 12134
rect 10420 12082 11152 12134
rect 11204 12082 11220 12134
rect 11272 12082 11288 12134
rect 11340 12082 11342 12134
rect 7370 12069 11342 12082
rect 7370 12038 7472 12069
rect 4900 12017 5632 12038
rect 5684 12017 5700 12038
rect 5752 12017 5768 12038
rect 5820 12017 6552 12038
rect 6604 12017 6620 12038
rect 6672 12017 6688 12038
rect 6740 12017 7472 12038
rect 7524 12017 7540 12069
rect 7592 12017 7608 12069
rect 7660 12017 8392 12069
rect 8444 12017 8460 12069
rect 8512 12017 8528 12069
rect 8580 12017 9312 12069
rect 9364 12017 9380 12069
rect 9432 12017 9448 12069
rect 9500 12017 10232 12069
rect 10284 12017 10300 12069
rect 10352 12017 10368 12069
rect 10420 12017 11152 12069
rect 11204 12017 11220 12069
rect 11272 12017 11288 12069
rect 11340 12017 11342 12069
rect 187 12014 11342 12017
rect 187 11962 2233 12014
rect 2285 11962 2335 12014
rect 2387 12010 5188 12014
rect 2387 11962 2872 12010
rect 187 11958 2872 11962
rect 2924 11958 2940 12010
rect 2992 11958 3008 12010
rect 3060 12004 5188 12010
rect 3060 11958 3792 12004
rect 187 11952 3792 11958
rect 3844 11952 3860 12004
rect 3912 11952 3928 12004
rect 3980 11952 4712 12004
rect 4764 11952 4780 12004
rect 4832 11952 4848 12004
rect 4900 11958 5188 12004
rect 5244 11958 5270 12014
rect 5326 11958 5352 12014
rect 5408 11958 5434 12014
rect 5490 11958 5516 12014
rect 5572 11958 5598 12014
rect 5654 12004 5680 12014
rect 5736 12004 5762 12014
rect 5818 12004 5844 12014
rect 5752 11958 5762 12004
rect 5820 11958 5844 12004
rect 5900 11958 5926 12014
rect 5982 11958 6008 12014
rect 6064 11958 6090 12014
rect 6146 11958 6172 12014
rect 6228 11958 6254 12014
rect 6310 11958 6336 12014
rect 6392 11958 6418 12014
rect 6474 11958 6500 12014
rect 6556 12004 6582 12014
rect 6638 12004 6664 12014
rect 6720 12004 6746 12014
rect 6740 11958 6746 12004
rect 6802 11958 6828 12014
rect 6884 11958 6909 12014
rect 6965 11958 6990 12014
rect 7046 11958 7071 12014
rect 7127 11958 7152 12014
rect 7208 11958 7233 12014
rect 7289 11958 7314 12014
rect 7370 12004 11342 12014
rect 7370 11958 7472 12004
rect 4900 11952 5632 11958
rect 5684 11952 5700 11958
rect 5752 11952 5768 11958
rect 5820 11952 6552 11958
rect 6604 11952 6620 11958
rect 6672 11952 6688 11958
rect 6740 11952 7472 11958
rect 7524 11952 7540 12004
rect 7592 11952 7608 12004
rect 7660 11952 8392 12004
rect 8444 11952 8460 12004
rect 8512 11952 8528 12004
rect 8580 11952 9312 12004
rect 9364 11952 9380 12004
rect 9432 11952 9448 12004
rect 9500 11952 10232 12004
rect 10284 11952 10300 12004
rect 10352 11952 10368 12004
rect 10420 11952 11152 12004
rect 11204 11952 11220 12004
rect 11272 11952 11288 12004
rect 11340 11952 11342 12004
rect 187 11950 11342 11952
rect 187 11898 2233 11950
rect 2285 11898 2335 11950
rect 2387 11944 11342 11950
rect 2387 11898 2872 11944
rect 187 11892 2872 11898
rect 2924 11892 2940 11944
rect 2992 11892 3008 11944
rect 3060 11939 11342 11944
rect 3060 11892 3792 11939
rect 187 11887 3792 11892
rect 3844 11887 3860 11939
rect 3912 11887 3928 11939
rect 3980 11887 4712 11939
rect 4764 11887 4780 11939
rect 4832 11887 4848 11939
rect 4900 11934 5632 11939
rect 5684 11934 5700 11939
rect 5752 11934 5768 11939
rect 5820 11934 6552 11939
rect 6604 11934 6620 11939
rect 6672 11934 6688 11939
rect 6740 11934 7472 11939
rect 4900 11887 5188 11934
rect 187 11886 5188 11887
rect 187 11834 2233 11886
rect 2285 11834 2335 11886
rect 2387 11878 5188 11886
rect 5244 11878 5270 11934
rect 5326 11878 5352 11934
rect 5408 11878 5434 11934
rect 5490 11878 5516 11934
rect 5572 11878 5598 11934
rect 5752 11887 5762 11934
rect 5820 11887 5844 11934
rect 5654 11878 5680 11887
rect 5736 11878 5762 11887
rect 5818 11878 5844 11887
rect 5900 11878 5926 11934
rect 5982 11878 6008 11934
rect 6064 11878 6090 11934
rect 6146 11878 6172 11934
rect 6228 11878 6254 11934
rect 6310 11878 6336 11934
rect 6392 11878 6418 11934
rect 6474 11878 6500 11934
rect 6740 11887 6746 11934
rect 6556 11878 6582 11887
rect 6638 11878 6664 11887
rect 6720 11878 6746 11887
rect 6802 11878 6828 11934
rect 6884 11878 6909 11934
rect 6965 11878 6990 11934
rect 7046 11878 7071 11934
rect 7127 11878 7152 11934
rect 7208 11878 7233 11934
rect 7289 11878 7314 11934
rect 7370 11887 7472 11934
rect 7524 11887 7540 11939
rect 7592 11887 7608 11939
rect 7660 11887 8392 11939
rect 8444 11887 8460 11939
rect 8512 11887 8528 11939
rect 8580 11887 9312 11939
rect 9364 11887 9380 11939
rect 9432 11887 9448 11939
rect 9500 11887 10232 11939
rect 10284 11887 10300 11939
rect 10352 11887 10368 11939
rect 10420 11887 11152 11939
rect 11204 11887 11220 11939
rect 11272 11887 11288 11939
rect 11340 11887 11342 11939
rect 7370 11878 11342 11887
rect 2387 11834 2872 11878
rect 187 11826 2872 11834
rect 2924 11826 2940 11878
rect 2992 11826 3008 11878
rect 3060 11874 11342 11878
rect 3060 11826 3792 11874
rect 187 11822 3792 11826
rect 3844 11822 3860 11874
rect 3912 11822 3928 11874
rect 3980 11822 4712 11874
rect 4764 11822 4780 11874
rect 4832 11822 4848 11874
rect 4900 11854 5632 11874
rect 5684 11854 5700 11874
rect 5752 11854 5768 11874
rect 5820 11854 6552 11874
rect 6604 11854 6620 11874
rect 6672 11854 6688 11874
rect 6740 11854 7472 11874
rect 4900 11822 5188 11854
rect 187 11770 2233 11822
rect 2285 11770 2335 11822
rect 2387 11812 5188 11822
rect 2387 11770 2872 11812
rect 187 11760 2872 11770
rect 2924 11760 2940 11812
rect 2992 11760 3008 11812
rect 3060 11809 5188 11812
rect 3060 11760 3792 11809
rect 187 11757 3792 11760
rect 3844 11757 3860 11809
rect 3912 11757 3928 11809
rect 3980 11757 4712 11809
rect 4764 11757 4780 11809
rect 4832 11757 4848 11809
rect 4900 11798 5188 11809
rect 5244 11798 5270 11854
rect 5326 11798 5352 11854
rect 5408 11798 5434 11854
rect 5490 11798 5516 11854
rect 5572 11798 5598 11854
rect 5752 11822 5762 11854
rect 5820 11822 5844 11854
rect 5654 11809 5680 11822
rect 5736 11809 5762 11822
rect 5818 11809 5844 11822
rect 5752 11798 5762 11809
rect 5820 11798 5844 11809
rect 5900 11798 5926 11854
rect 5982 11798 6008 11854
rect 6064 11798 6090 11854
rect 6146 11798 6172 11854
rect 6228 11798 6254 11854
rect 6310 11798 6336 11854
rect 6392 11798 6418 11854
rect 6474 11798 6500 11854
rect 6740 11822 6746 11854
rect 6556 11809 6582 11822
rect 6638 11809 6664 11822
rect 6720 11809 6746 11822
rect 6740 11798 6746 11809
rect 6802 11798 6828 11854
rect 6884 11798 6909 11854
rect 6965 11798 6990 11854
rect 7046 11798 7071 11854
rect 7127 11798 7152 11854
rect 7208 11798 7233 11854
rect 7289 11798 7314 11854
rect 7370 11822 7472 11854
rect 7524 11822 7540 11874
rect 7592 11822 7608 11874
rect 7660 11822 8392 11874
rect 8444 11822 8460 11874
rect 8512 11822 8528 11874
rect 8580 11822 9312 11874
rect 9364 11822 9380 11874
rect 9432 11822 9448 11874
rect 9500 11822 10232 11874
rect 10284 11822 10300 11874
rect 10352 11822 10368 11874
rect 10420 11822 11152 11874
rect 11204 11822 11220 11874
rect 11272 11822 11288 11874
rect 11340 11822 11342 11874
rect 7370 11809 11342 11822
rect 7370 11798 7472 11809
rect 4900 11774 5632 11798
rect 5684 11774 5700 11798
rect 5752 11774 5768 11798
rect 5820 11774 6552 11798
rect 6604 11774 6620 11798
rect 6672 11774 6688 11798
rect 6740 11774 7472 11798
rect 4900 11757 5188 11774
rect 187 11705 2233 11757
rect 2285 11705 2335 11757
rect 2387 11746 5188 11757
rect 2387 11705 2872 11746
rect 187 11694 2872 11705
rect 2924 11694 2940 11746
rect 2992 11694 3008 11746
rect 3060 11744 5188 11746
rect 3060 11694 3792 11744
rect 187 11692 3792 11694
rect 3844 11692 3860 11744
rect 3912 11692 3928 11744
rect 3980 11692 4712 11744
rect 4764 11692 4780 11744
rect 4832 11692 4848 11744
rect 4900 11718 5188 11744
rect 5244 11718 5270 11774
rect 5326 11718 5352 11774
rect 5408 11718 5434 11774
rect 5490 11718 5516 11774
rect 5572 11718 5598 11774
rect 5752 11757 5762 11774
rect 5820 11757 5844 11774
rect 5654 11744 5680 11757
rect 5736 11744 5762 11757
rect 5818 11744 5844 11757
rect 5752 11718 5762 11744
rect 5820 11718 5844 11744
rect 5900 11718 5926 11774
rect 5982 11718 6008 11774
rect 6064 11718 6090 11774
rect 6146 11718 6172 11774
rect 6228 11718 6254 11774
rect 6310 11718 6336 11774
rect 6392 11718 6418 11774
rect 6474 11718 6500 11774
rect 6740 11757 6746 11774
rect 6556 11744 6582 11757
rect 6638 11744 6664 11757
rect 6720 11744 6746 11757
rect 6740 11718 6746 11744
rect 6802 11718 6828 11774
rect 6884 11718 6909 11774
rect 6965 11718 6990 11774
rect 7046 11718 7071 11774
rect 7127 11718 7152 11774
rect 7208 11718 7233 11774
rect 7289 11718 7314 11774
rect 7370 11757 7472 11774
rect 7524 11757 7540 11809
rect 7592 11757 7608 11809
rect 7660 11757 8392 11809
rect 8444 11757 8460 11809
rect 8512 11757 8528 11809
rect 8580 11757 9312 11809
rect 9364 11757 9380 11809
rect 9432 11757 9448 11809
rect 9500 11757 10232 11809
rect 10284 11757 10300 11809
rect 10352 11757 10368 11809
rect 10420 11757 11152 11809
rect 11204 11757 11220 11809
rect 11272 11757 11288 11809
rect 11340 11757 11342 11809
rect 7370 11744 11342 11757
rect 7370 11718 7472 11744
rect 4900 11694 5632 11718
rect 5684 11694 5700 11718
rect 5752 11694 5768 11718
rect 5820 11694 6552 11718
rect 6604 11694 6620 11718
rect 6672 11694 6688 11718
rect 6740 11694 7472 11718
rect 4900 11692 5188 11694
rect 187 11640 2233 11692
rect 2285 11640 2335 11692
rect 2387 11680 5188 11692
rect 2387 11640 2872 11680
rect 187 11628 2872 11640
rect 2924 11628 2940 11680
rect 2992 11628 3008 11680
rect 3060 11679 5188 11680
rect 3060 11628 3792 11679
rect 187 11627 3792 11628
rect 3844 11627 3860 11679
rect 3912 11627 3928 11679
rect 3980 11627 4712 11679
rect 4764 11627 4780 11679
rect 4832 11627 4848 11679
rect 4900 11638 5188 11679
rect 5244 11638 5270 11694
rect 5326 11638 5352 11694
rect 5408 11638 5434 11694
rect 5490 11638 5516 11694
rect 5572 11638 5598 11694
rect 5752 11692 5762 11694
rect 5820 11692 5844 11694
rect 5654 11679 5680 11692
rect 5736 11679 5762 11692
rect 5818 11679 5844 11692
rect 5752 11638 5762 11679
rect 5820 11638 5844 11679
rect 5900 11638 5926 11694
rect 5982 11638 6008 11694
rect 6064 11638 6090 11694
rect 6146 11638 6172 11694
rect 6228 11638 6254 11694
rect 6310 11638 6336 11694
rect 6392 11638 6418 11694
rect 6474 11638 6500 11694
rect 6740 11692 6746 11694
rect 6556 11679 6582 11692
rect 6638 11679 6664 11692
rect 6720 11679 6746 11692
rect 6740 11638 6746 11679
rect 6802 11638 6828 11694
rect 6884 11638 6909 11694
rect 6965 11638 6990 11694
rect 7046 11638 7071 11694
rect 7127 11638 7152 11694
rect 7208 11638 7233 11694
rect 7289 11638 7314 11694
rect 7370 11692 7472 11694
rect 7524 11692 7540 11744
rect 7592 11692 7608 11744
rect 7660 11692 8392 11744
rect 8444 11692 8460 11744
rect 8512 11692 8528 11744
rect 8580 11692 9312 11744
rect 9364 11692 9380 11744
rect 9432 11692 9448 11744
rect 9500 11692 10232 11744
rect 10284 11692 10300 11744
rect 10352 11692 10368 11744
rect 10420 11692 11152 11744
rect 11204 11692 11220 11744
rect 11272 11692 11288 11744
rect 11340 11692 11342 11744
rect 7370 11679 11342 11692
rect 7370 11638 7472 11679
rect 4900 11627 5632 11638
rect 5684 11627 5700 11638
rect 5752 11627 5768 11638
rect 5820 11627 6552 11638
rect 6604 11627 6620 11638
rect 6672 11627 6688 11638
rect 6740 11627 7472 11638
rect 7524 11627 7540 11679
rect 7592 11627 7608 11679
rect 7660 11627 8392 11679
rect 8444 11627 8460 11679
rect 8512 11627 8528 11679
rect 8580 11627 9312 11679
rect 9364 11627 9380 11679
rect 9432 11627 9448 11679
rect 9500 11627 10232 11679
rect 10284 11627 10300 11679
rect 10352 11627 10368 11679
rect 10420 11627 11152 11679
rect 11204 11627 11220 11679
rect 11272 11627 11288 11679
rect 11340 11627 11342 11679
rect 187 11575 2233 11627
rect 2285 11575 2335 11627
rect 2387 11614 11342 11627
rect 2387 11575 2872 11614
rect 187 11562 2872 11575
rect 2924 11562 2940 11614
rect 2992 11562 3008 11614
rect 3060 11562 3792 11614
rect 3844 11562 3860 11614
rect 3912 11562 3928 11614
rect 3980 11562 4712 11614
rect 4764 11562 4780 11614
rect 4832 11562 4848 11614
rect 4900 11562 5188 11614
rect 187 11510 2233 11562
rect 2285 11510 2335 11562
rect 2387 11558 5188 11562
rect 5244 11558 5270 11614
rect 5326 11558 5352 11614
rect 5408 11558 5434 11614
rect 5490 11558 5516 11614
rect 5572 11558 5598 11614
rect 5752 11562 5762 11614
rect 5820 11562 5844 11614
rect 5654 11558 5680 11562
rect 5736 11558 5762 11562
rect 5818 11558 5844 11562
rect 5900 11558 5926 11614
rect 5982 11558 6008 11614
rect 6064 11558 6090 11614
rect 6146 11558 6172 11614
rect 6228 11558 6254 11614
rect 6310 11558 6336 11614
rect 6392 11558 6418 11614
rect 6474 11558 6500 11614
rect 6740 11562 6746 11614
rect 6556 11558 6582 11562
rect 6638 11558 6664 11562
rect 6720 11558 6746 11562
rect 6802 11558 6828 11614
rect 6884 11558 6909 11614
rect 6965 11558 6990 11614
rect 7046 11558 7071 11614
rect 7127 11558 7152 11614
rect 7208 11558 7233 11614
rect 7289 11558 7314 11614
rect 7370 11562 7472 11614
rect 7524 11562 7540 11614
rect 7592 11562 7608 11614
rect 7660 11562 8392 11614
rect 8444 11562 8460 11614
rect 8512 11562 8528 11614
rect 8580 11562 9312 11614
rect 9364 11562 9380 11614
rect 9432 11562 9448 11614
rect 9500 11562 10232 11614
rect 10284 11562 10300 11614
rect 10352 11562 10368 11614
rect 10420 11562 11152 11614
rect 11204 11562 11220 11614
rect 11272 11562 11288 11614
rect 11340 11562 11342 11614
rect 7370 11558 11342 11562
rect 2387 11556 11342 11558
rect 2387 11510 3342 11556
rect 187 11497 3342 11510
rect 187 11445 2233 11497
rect 2285 11445 2335 11497
rect 2387 11445 3342 11497
rect 187 11432 3342 11445
rect 187 11380 2233 11432
rect 2285 11380 2335 11432
rect 2387 11380 3342 11432
rect 187 11367 3342 11380
rect 187 11315 2233 11367
rect 2285 11315 2335 11367
rect 2387 11361 3342 11367
tri 3342 11361 3537 11556 nw
rect 2387 11315 2824 11361
rect 187 11302 2824 11315
rect 187 11250 2233 11302
rect 2285 11250 2335 11302
rect 2387 11250 2824 11302
rect 187 11237 2824 11250
rect 187 11185 2233 11237
rect 2285 11185 2335 11237
rect 2387 11185 2824 11237
rect 187 11172 2824 11185
rect 187 11120 2233 11172
rect 2285 11120 2335 11172
rect 2387 11120 2824 11172
rect 187 11107 2824 11120
rect 187 11055 2233 11107
rect 2285 11055 2335 11107
rect 2387 11055 2824 11107
rect 187 11042 2824 11055
rect 187 10990 2233 11042
rect 2285 10990 2335 11042
rect 2387 10990 2824 11042
rect 187 10977 2824 10990
rect 187 10925 2233 10977
rect 2285 10925 2335 10977
rect 2387 10925 2824 10977
rect 187 10912 2824 10925
rect 187 10860 2233 10912
rect 2285 10860 2335 10912
rect 2387 10860 2824 10912
rect 187 10847 2824 10860
rect 187 10795 2233 10847
rect 2285 10795 2335 10847
rect 2387 10795 2824 10847
tri 2824 10843 3342 11361 nw
tri 11505 11231 12222 11948 se
rect 12222 11231 14858 14091
tri 3492 10953 3770 11231 se
rect 3770 11229 14858 11231
rect 3770 11225 7587 11229
rect 3770 11173 4281 11225
rect 4333 11173 4359 11225
rect 4411 11173 5201 11225
rect 5253 11173 5279 11225
rect 5331 11173 6121 11225
rect 6173 11173 6199 11225
rect 6251 11173 7041 11225
rect 7093 11173 7119 11225
rect 7171 11173 7587 11225
rect 7643 11173 7669 11229
rect 7725 11173 7751 11229
rect 7807 11173 7833 11229
rect 7889 11173 7915 11229
rect 7971 11225 7997 11229
rect 8053 11225 8079 11229
rect 8135 11173 8161 11229
rect 8217 11173 8243 11229
rect 8299 11173 8325 11229
rect 8381 11173 8407 11229
rect 8463 11173 8489 11229
rect 8545 11173 8571 11229
rect 8627 11173 8653 11229
rect 8709 11173 8735 11229
rect 8791 11173 8817 11229
rect 8873 11225 8899 11229
rect 8955 11225 8981 11229
rect 8873 11173 8881 11225
rect 8955 11173 8959 11225
rect 9037 11173 9063 11229
rect 9119 11173 9145 11229
rect 9201 11173 9227 11229
rect 9283 11173 9308 11229
rect 9364 11173 9389 11229
rect 9445 11173 9470 11229
rect 9526 11173 9551 11229
rect 9607 11173 9632 11229
rect 9688 11173 9713 11229
rect 9769 11225 14858 11229
rect 9769 11173 9801 11225
rect 9853 11173 9879 11225
rect 9931 11173 10721 11225
rect 10773 11173 10799 11225
rect 10851 11173 11641 11225
rect 11693 11173 11719 11225
rect 11771 11173 12561 11225
rect 12613 11173 12639 11225
rect 12691 11173 14858 11225
rect 3770 11161 14858 11173
rect 3770 11109 4281 11161
rect 4333 11109 4359 11161
rect 4411 11109 5201 11161
rect 5253 11109 5279 11161
rect 5331 11109 6121 11161
rect 6173 11109 6199 11161
rect 6251 11109 7041 11161
rect 7093 11109 7119 11161
rect 7171 11149 7961 11161
rect 8013 11149 8039 11161
rect 8091 11149 8881 11161
rect 8933 11149 8959 11161
rect 9011 11149 9801 11161
rect 7171 11109 7587 11149
rect 3770 11097 7587 11109
rect 3770 11045 4281 11097
rect 4333 11045 4359 11097
rect 4411 11045 5201 11097
rect 5253 11045 5279 11097
rect 5331 11045 6121 11097
rect 6173 11045 6199 11097
rect 6251 11045 7041 11097
rect 7093 11045 7119 11097
rect 7171 11093 7587 11097
rect 7643 11093 7669 11149
rect 7725 11093 7751 11149
rect 7807 11093 7833 11149
rect 7889 11093 7915 11149
rect 7971 11097 7997 11109
rect 8053 11097 8079 11109
rect 8135 11093 8161 11149
rect 8217 11093 8243 11149
rect 8299 11093 8325 11149
rect 8381 11093 8407 11149
rect 8463 11093 8489 11149
rect 8545 11093 8571 11149
rect 8627 11093 8653 11149
rect 8709 11093 8735 11149
rect 8791 11093 8817 11149
rect 8873 11109 8881 11149
rect 8955 11109 8959 11149
rect 8873 11097 8899 11109
rect 8955 11097 8981 11109
rect 8873 11093 8881 11097
rect 8955 11093 8959 11097
rect 9037 11093 9063 11149
rect 9119 11093 9145 11149
rect 9201 11093 9227 11149
rect 9283 11093 9308 11149
rect 9364 11093 9389 11149
rect 9445 11093 9470 11149
rect 9526 11093 9551 11149
rect 9607 11093 9632 11149
rect 9688 11093 9713 11149
rect 9769 11109 9801 11149
rect 9853 11109 9879 11161
rect 9931 11109 10721 11161
rect 10773 11109 10799 11161
rect 10851 11109 11641 11161
rect 11693 11109 11719 11161
rect 11771 11109 12561 11161
rect 12613 11109 12639 11161
rect 12691 11109 14858 11161
rect 9769 11097 14858 11109
rect 9769 11093 9801 11097
rect 7171 11069 7961 11093
rect 8013 11069 8039 11093
rect 8091 11069 8881 11093
rect 8933 11069 8959 11093
rect 9011 11069 9801 11093
rect 7171 11045 7587 11069
rect 3770 11033 7587 11045
rect 3770 10981 4281 11033
rect 4333 10981 4359 11033
rect 4411 10981 5201 11033
rect 5253 10981 5279 11033
rect 5331 10981 6121 11033
rect 6173 10981 6199 11033
rect 6251 10981 7041 11033
rect 7093 10981 7119 11033
rect 7171 11013 7587 11033
rect 7643 11013 7669 11069
rect 7725 11013 7751 11069
rect 7807 11013 7833 11069
rect 7889 11013 7915 11069
rect 7971 11033 7997 11045
rect 8053 11033 8079 11045
rect 8135 11013 8161 11069
rect 8217 11013 8243 11069
rect 8299 11013 8325 11069
rect 8381 11013 8407 11069
rect 8463 11013 8489 11069
rect 8545 11013 8571 11069
rect 8627 11013 8653 11069
rect 8709 11013 8735 11069
rect 8791 11013 8817 11069
rect 8873 11045 8881 11069
rect 8955 11045 8959 11069
rect 8873 11033 8899 11045
rect 8955 11033 8981 11045
rect 8873 11013 8881 11033
rect 8955 11013 8959 11033
rect 9037 11013 9063 11069
rect 9119 11013 9145 11069
rect 9201 11013 9227 11069
rect 9283 11013 9308 11069
rect 9364 11013 9389 11069
rect 9445 11013 9470 11069
rect 9526 11013 9551 11069
rect 9607 11013 9632 11069
rect 9688 11013 9713 11069
rect 9769 11045 9801 11069
rect 9853 11045 9879 11097
rect 9931 11045 10721 11097
rect 10773 11045 10799 11097
rect 10851 11045 11641 11097
rect 11693 11045 11719 11097
rect 11771 11045 12561 11097
rect 12613 11045 12639 11097
rect 12691 11045 14858 11097
rect 9769 11033 14858 11045
rect 9769 11013 9801 11033
rect 7171 10989 7961 11013
rect 8013 10989 8039 11013
rect 8091 10989 8881 11013
rect 8933 10989 8959 11013
rect 9011 10989 9801 11013
rect 7171 10981 7587 10989
rect 3770 10969 7587 10981
rect 3770 10953 4281 10969
rect 3361 10947 4281 10953
rect 3413 10895 3439 10947
rect 3491 10917 4281 10947
rect 4333 10917 4359 10969
rect 4411 10917 5201 10969
rect 5253 10917 5279 10969
rect 5331 10917 6121 10969
rect 6173 10917 6199 10969
rect 6251 10917 7041 10969
rect 7093 10917 7119 10969
rect 7171 10933 7587 10969
rect 7643 10933 7669 10989
rect 7725 10933 7751 10989
rect 7807 10933 7833 10989
rect 7889 10933 7915 10989
rect 7971 10969 7997 10981
rect 8053 10969 8079 10981
rect 8135 10933 8161 10989
rect 8217 10933 8243 10989
rect 8299 10933 8325 10989
rect 8381 10933 8407 10989
rect 8463 10933 8489 10989
rect 8545 10933 8571 10989
rect 8627 10933 8653 10989
rect 8709 10933 8735 10989
rect 8791 10933 8817 10989
rect 8873 10981 8881 10989
rect 8955 10981 8959 10989
rect 8873 10969 8899 10981
rect 8955 10969 8981 10981
rect 8873 10933 8881 10969
rect 8955 10933 8959 10969
rect 9037 10933 9063 10989
rect 9119 10933 9145 10989
rect 9201 10933 9227 10989
rect 9283 10933 9308 10989
rect 9364 10933 9389 10989
rect 9445 10933 9470 10989
rect 9526 10933 9551 10989
rect 9607 10933 9632 10989
rect 9688 10933 9713 10989
rect 9769 10981 9801 10989
rect 9853 10981 9879 11033
rect 9931 10981 10721 11033
rect 10773 10981 10799 11033
rect 10851 10981 11641 11033
rect 11693 10981 11719 11033
rect 11771 10981 12561 11033
rect 12613 10981 12639 11033
rect 12691 10981 14858 11033
rect 9769 10969 14858 10981
rect 9769 10933 9801 10969
rect 7171 10917 7961 10933
rect 8013 10917 8039 10933
rect 8091 10917 8881 10933
rect 8933 10917 8959 10933
rect 9011 10917 9801 10933
rect 9853 10917 9879 10969
rect 9931 10917 10721 10969
rect 10773 10917 10799 10969
rect 10851 10917 11641 10969
rect 11693 10917 11719 10969
rect 11771 10917 12561 10969
rect 12613 10917 12639 10969
rect 12691 10917 14858 10969
rect 3491 10909 14858 10917
rect 3491 10905 7587 10909
rect 3491 10895 4281 10905
rect 3361 10881 4281 10895
rect 187 10782 2824 10795
rect 187 10730 2233 10782
rect 2285 10730 2335 10782
rect 2387 10730 2824 10782
rect 187 10717 2824 10730
rect 187 10665 2233 10717
rect 2285 10665 2335 10717
rect 2387 10665 2824 10717
rect 187 10652 2824 10665
rect 187 10600 2233 10652
rect 2285 10600 2335 10652
rect 2387 10600 2824 10652
rect 187 10587 2824 10600
rect 187 10535 2233 10587
rect 2285 10535 2335 10587
rect 2387 10535 2824 10587
rect 187 10522 2824 10535
rect 187 10470 2233 10522
rect 2285 10470 2335 10522
rect 2387 10470 2824 10522
rect 187 10457 2824 10470
rect 187 10405 2233 10457
rect 2285 10405 2335 10457
rect 2387 10405 2824 10457
rect 187 10392 2824 10405
rect 187 10340 2233 10392
rect 2285 10340 2335 10392
rect 2387 10340 2824 10392
rect 187 10327 2824 10340
rect 187 10275 2233 10327
rect 2285 10275 2335 10327
rect 2387 10275 2824 10327
rect 187 10262 2824 10275
rect 187 10210 2233 10262
rect 2285 10210 2335 10262
rect 2387 10210 2824 10262
rect 187 10197 2824 10210
rect 187 10145 2233 10197
rect 2285 10145 2335 10197
rect 2387 10145 2824 10197
rect 187 10132 2824 10145
rect 187 10080 2233 10132
rect 2285 10080 2335 10132
rect 2387 10080 2824 10132
rect 187 10067 2824 10080
rect 187 10015 2233 10067
rect 2285 10015 2335 10067
rect 2387 10015 2824 10067
rect 187 10002 2824 10015
rect 187 9950 2233 10002
rect 2285 9950 2335 10002
rect 2387 9950 2824 10002
rect 187 9937 2824 9950
rect 187 9885 2233 9937
rect 2285 9885 2335 9937
rect 2387 9885 2824 9937
rect 187 9872 2824 9885
rect 187 9820 2233 9872
rect 2285 9820 2335 9872
rect 2387 9820 2824 9872
rect 187 9807 2824 9820
rect 187 9755 2233 9807
rect 2285 9755 2335 9807
rect 2387 9755 2824 9807
rect 187 9742 2824 9755
rect 187 9690 2233 9742
rect 2285 9690 2335 9742
rect 2387 9690 2824 9742
rect 187 9677 2824 9690
rect 187 9625 2233 9677
rect 2285 9625 2335 9677
rect 2387 9625 2824 9677
rect 187 9612 2824 9625
rect 187 9560 2233 9612
rect 2285 9560 2335 9612
rect 2387 9560 2824 9612
rect 187 9547 2824 9560
rect 187 9495 2233 9547
rect 2285 9495 2335 9547
rect 2387 9495 2824 9547
rect 187 9482 2824 9495
rect 3413 10829 3439 10881
rect 3491 10853 4281 10881
rect 4333 10853 4359 10905
rect 4411 10853 5201 10905
rect 5253 10853 5279 10905
rect 5331 10853 6121 10905
rect 6173 10853 6199 10905
rect 6251 10853 7041 10905
rect 7093 10853 7119 10905
rect 7171 10853 7587 10905
rect 7643 10853 7669 10909
rect 7725 10853 7751 10909
rect 7807 10853 7833 10909
rect 7889 10853 7915 10909
rect 7971 10905 7997 10909
rect 8053 10905 8079 10909
rect 8135 10853 8161 10909
rect 8217 10853 8243 10909
rect 8299 10853 8325 10909
rect 8381 10853 8407 10909
rect 8463 10853 8489 10909
rect 8545 10853 8571 10909
rect 8627 10853 8653 10909
rect 8709 10853 8735 10909
rect 8791 10853 8817 10909
rect 8873 10905 8899 10909
rect 8955 10905 8981 10909
rect 8873 10853 8881 10905
rect 8955 10853 8959 10905
rect 9037 10853 9063 10909
rect 9119 10853 9145 10909
rect 9201 10853 9227 10909
rect 9283 10853 9308 10909
rect 9364 10853 9389 10909
rect 9445 10853 9470 10909
rect 9526 10853 9551 10909
rect 9607 10853 9632 10909
rect 9688 10853 9713 10909
rect 9769 10905 14858 10909
rect 9769 10853 9801 10905
rect 9853 10853 9879 10905
rect 9931 10853 10721 10905
rect 10773 10853 10799 10905
rect 10851 10853 11641 10905
rect 11693 10853 11719 10905
rect 11771 10853 12561 10905
rect 12613 10853 12639 10905
rect 12691 10853 14858 10905
rect 3491 10841 14858 10853
rect 3491 10829 4281 10841
rect 3361 10815 4281 10829
rect 3413 10763 3439 10815
rect 3491 10789 4281 10815
rect 4333 10789 4359 10841
rect 4411 10789 5201 10841
rect 5253 10789 5279 10841
rect 5331 10789 6121 10841
rect 6173 10789 6199 10841
rect 6251 10789 7041 10841
rect 7093 10789 7119 10841
rect 7171 10829 7961 10841
rect 8013 10829 8039 10841
rect 8091 10829 8881 10841
rect 8933 10829 8959 10841
rect 9011 10829 9801 10841
rect 7171 10789 7587 10829
rect 3491 10777 7587 10789
rect 3491 10763 4281 10777
rect 3361 10749 4281 10763
rect 3413 10697 3439 10749
rect 3491 10725 4281 10749
rect 4333 10725 4359 10777
rect 4411 10725 5201 10777
rect 5253 10725 5279 10777
rect 5331 10725 6121 10777
rect 6173 10725 6199 10777
rect 6251 10725 7041 10777
rect 7093 10725 7119 10777
rect 7171 10773 7587 10777
rect 7643 10773 7669 10829
rect 7725 10773 7751 10829
rect 7807 10773 7833 10829
rect 7889 10773 7915 10829
rect 7971 10777 7997 10789
rect 8053 10777 8079 10789
rect 8135 10773 8161 10829
rect 8217 10773 8243 10829
rect 8299 10773 8325 10829
rect 8381 10773 8407 10829
rect 8463 10773 8489 10829
rect 8545 10773 8571 10829
rect 8627 10773 8653 10829
rect 8709 10773 8735 10829
rect 8791 10773 8817 10829
rect 8873 10789 8881 10829
rect 8955 10789 8959 10829
rect 8873 10777 8899 10789
rect 8955 10777 8981 10789
rect 8873 10773 8881 10777
rect 8955 10773 8959 10777
rect 9037 10773 9063 10829
rect 9119 10773 9145 10829
rect 9201 10773 9227 10829
rect 9283 10773 9308 10829
rect 9364 10773 9389 10829
rect 9445 10773 9470 10829
rect 9526 10773 9551 10829
rect 9607 10773 9632 10829
rect 9688 10773 9713 10829
rect 9769 10789 9801 10829
rect 9853 10789 9879 10841
rect 9931 10789 10721 10841
rect 10773 10789 10799 10841
rect 10851 10789 11641 10841
rect 11693 10789 11719 10841
rect 11771 10789 12561 10841
rect 12613 10789 12639 10841
rect 12691 10789 14858 10841
rect 9769 10777 14858 10789
rect 9769 10773 9801 10777
rect 7171 10749 7961 10773
rect 8013 10749 8039 10773
rect 8091 10749 8881 10773
rect 8933 10749 8959 10773
rect 9011 10749 9801 10773
rect 7171 10725 7587 10749
rect 3491 10713 7587 10725
rect 3491 10697 4281 10713
rect 3361 10683 4281 10697
rect 3413 10631 3439 10683
rect 3491 10661 4281 10683
rect 4333 10661 4359 10713
rect 4411 10661 5201 10713
rect 5253 10661 5279 10713
rect 5331 10661 6121 10713
rect 6173 10661 6199 10713
rect 6251 10661 7041 10713
rect 7093 10661 7119 10713
rect 7171 10693 7587 10713
rect 7643 10693 7669 10749
rect 7725 10693 7751 10749
rect 7807 10693 7833 10749
rect 7889 10693 7915 10749
rect 7971 10713 7997 10725
rect 8053 10713 8079 10725
rect 8135 10693 8161 10749
rect 8217 10693 8243 10749
rect 8299 10693 8325 10749
rect 8381 10693 8407 10749
rect 8463 10693 8489 10749
rect 8545 10693 8571 10749
rect 8627 10693 8653 10749
rect 8709 10693 8735 10749
rect 8791 10693 8817 10749
rect 8873 10725 8881 10749
rect 8955 10725 8959 10749
rect 8873 10713 8899 10725
rect 8955 10713 8981 10725
rect 8873 10693 8881 10713
rect 8955 10693 8959 10713
rect 9037 10693 9063 10749
rect 9119 10693 9145 10749
rect 9201 10693 9227 10749
rect 9283 10693 9308 10749
rect 9364 10693 9389 10749
rect 9445 10693 9470 10749
rect 9526 10693 9551 10749
rect 9607 10693 9632 10749
rect 9688 10693 9713 10749
rect 9769 10725 9801 10749
rect 9853 10725 9879 10777
rect 9931 10725 10721 10777
rect 10773 10725 10799 10777
rect 10851 10725 11641 10777
rect 11693 10725 11719 10777
rect 11771 10725 12561 10777
rect 12613 10725 12639 10777
rect 12691 10725 14858 10777
rect 9769 10713 14858 10725
rect 9769 10693 9801 10713
rect 7171 10669 7961 10693
rect 8013 10669 8039 10693
rect 8091 10669 8881 10693
rect 8933 10669 8959 10693
rect 9011 10669 9801 10693
rect 7171 10661 7587 10669
rect 3491 10649 7587 10661
rect 3491 10631 4281 10649
rect 3361 10617 4281 10631
rect 3413 10565 3439 10617
rect 3491 10597 4281 10617
rect 4333 10597 4359 10649
rect 4411 10597 5201 10649
rect 5253 10597 5279 10649
rect 5331 10597 6121 10649
rect 6173 10597 6199 10649
rect 6251 10597 7041 10649
rect 7093 10597 7119 10649
rect 7171 10613 7587 10649
rect 7643 10613 7669 10669
rect 7725 10613 7751 10669
rect 7807 10613 7833 10669
rect 7889 10613 7915 10669
rect 7971 10649 7997 10661
rect 8053 10649 8079 10661
rect 8135 10613 8161 10669
rect 8217 10613 8243 10669
rect 8299 10613 8325 10669
rect 8381 10613 8407 10669
rect 8463 10613 8489 10669
rect 8545 10613 8571 10669
rect 8627 10613 8653 10669
rect 8709 10613 8735 10669
rect 8791 10613 8817 10669
rect 8873 10661 8881 10669
rect 8955 10661 8959 10669
rect 8873 10649 8899 10661
rect 8955 10649 8981 10661
rect 8873 10613 8881 10649
rect 8955 10613 8959 10649
rect 9037 10613 9063 10669
rect 9119 10613 9145 10669
rect 9201 10613 9227 10669
rect 9283 10613 9308 10669
rect 9364 10613 9389 10669
rect 9445 10613 9470 10669
rect 9526 10613 9551 10669
rect 9607 10613 9632 10669
rect 9688 10613 9713 10669
rect 9769 10661 9801 10669
rect 9853 10661 9879 10713
rect 9931 10661 10721 10713
rect 10773 10661 10799 10713
rect 10851 10661 11641 10713
rect 11693 10661 11719 10713
rect 11771 10661 12561 10713
rect 12613 10661 12639 10713
rect 12691 10661 14858 10713
rect 9769 10649 14858 10661
rect 9769 10613 9801 10649
rect 7171 10597 7961 10613
rect 8013 10597 8039 10613
rect 8091 10597 8881 10613
rect 8933 10597 8959 10613
rect 9011 10597 9801 10613
rect 9853 10597 9879 10649
rect 9931 10597 10721 10649
rect 10773 10597 10799 10649
rect 10851 10597 11641 10649
rect 11693 10597 11719 10649
rect 11771 10597 12561 10649
rect 12613 10597 12639 10649
rect 12691 10597 14858 10649
rect 3491 10589 14858 10597
rect 3491 10585 7587 10589
rect 3491 10565 4281 10585
rect 3361 10551 4281 10565
rect 3413 10499 3439 10551
rect 3491 10533 4281 10551
rect 4333 10533 4359 10585
rect 4411 10533 5201 10585
rect 5253 10533 5279 10585
rect 5331 10533 6121 10585
rect 6173 10533 6199 10585
rect 6251 10533 7041 10585
rect 7093 10533 7119 10585
rect 7171 10533 7587 10585
rect 7643 10533 7669 10589
rect 7725 10533 7751 10589
rect 7807 10533 7833 10589
rect 7889 10533 7915 10589
rect 7971 10585 7997 10589
rect 8053 10585 8079 10589
rect 8135 10533 8161 10589
rect 8217 10533 8243 10589
rect 8299 10533 8325 10589
rect 8381 10533 8407 10589
rect 8463 10533 8489 10589
rect 8545 10533 8571 10589
rect 8627 10533 8653 10589
rect 8709 10533 8735 10589
rect 8791 10533 8817 10589
rect 8873 10585 8899 10589
rect 8955 10585 8981 10589
rect 8873 10533 8881 10585
rect 8955 10533 8959 10585
rect 9037 10533 9063 10589
rect 9119 10533 9145 10589
rect 9201 10533 9227 10589
rect 9283 10533 9308 10589
rect 9364 10533 9389 10589
rect 9445 10533 9470 10589
rect 9526 10533 9551 10589
rect 9607 10533 9632 10589
rect 9688 10533 9713 10589
rect 9769 10585 14858 10589
rect 9769 10533 9801 10585
rect 9853 10533 9879 10585
rect 9931 10533 10721 10585
rect 10773 10533 10799 10585
rect 10851 10533 11641 10585
rect 11693 10533 11719 10585
rect 11771 10533 12561 10585
rect 12613 10533 12639 10585
rect 12691 10533 14858 10585
rect 3491 10521 14858 10533
rect 3491 10499 4281 10521
rect 3361 10485 4281 10499
rect 3413 10433 3439 10485
rect 3491 10469 4281 10485
rect 4333 10469 4359 10521
rect 4411 10469 5201 10521
rect 5253 10469 5279 10521
rect 5331 10469 6121 10521
rect 6173 10469 6199 10521
rect 6251 10469 7041 10521
rect 7093 10469 7119 10521
rect 7171 10509 7961 10521
rect 8013 10509 8039 10521
rect 8091 10509 8881 10521
rect 8933 10509 8959 10521
rect 9011 10509 9801 10521
rect 7171 10469 7587 10509
rect 3491 10457 7587 10469
rect 3491 10433 4281 10457
rect 3361 10419 4281 10433
rect 3413 10367 3439 10419
rect 3491 10405 4281 10419
rect 4333 10405 4359 10457
rect 4411 10405 5201 10457
rect 5253 10405 5279 10457
rect 5331 10405 6121 10457
rect 6173 10405 6199 10457
rect 6251 10405 7041 10457
rect 7093 10405 7119 10457
rect 7171 10453 7587 10457
rect 7643 10453 7669 10509
rect 7725 10453 7751 10509
rect 7807 10453 7833 10509
rect 7889 10453 7915 10509
rect 7971 10457 7997 10469
rect 8053 10457 8079 10469
rect 8135 10453 8161 10509
rect 8217 10453 8243 10509
rect 8299 10453 8325 10509
rect 8381 10453 8407 10509
rect 8463 10453 8489 10509
rect 8545 10453 8571 10509
rect 8627 10453 8653 10509
rect 8709 10453 8735 10509
rect 8791 10453 8817 10509
rect 8873 10469 8881 10509
rect 8955 10469 8959 10509
rect 8873 10457 8899 10469
rect 8955 10457 8981 10469
rect 8873 10453 8881 10457
rect 8955 10453 8959 10457
rect 9037 10453 9063 10509
rect 9119 10453 9145 10509
rect 9201 10453 9227 10509
rect 9283 10453 9308 10509
rect 9364 10453 9389 10509
rect 9445 10453 9470 10509
rect 9526 10453 9551 10509
rect 9607 10453 9632 10509
rect 9688 10453 9713 10509
rect 9769 10469 9801 10509
rect 9853 10469 9879 10521
rect 9931 10469 10721 10521
rect 10773 10469 10799 10521
rect 10851 10469 11641 10521
rect 11693 10469 11719 10521
rect 11771 10469 12561 10521
rect 12613 10469 12639 10521
rect 12691 10469 14858 10521
rect 9769 10457 14858 10469
rect 9769 10453 9801 10457
rect 7171 10429 7961 10453
rect 8013 10429 8039 10453
rect 8091 10429 8881 10453
rect 8933 10429 8959 10453
rect 9011 10429 9801 10453
rect 7171 10405 7587 10429
rect 3491 10393 7587 10405
rect 3491 10367 4281 10393
rect 3361 10353 4281 10367
rect 3413 10301 3439 10353
rect 3491 10341 4281 10353
rect 4333 10341 4359 10393
rect 4411 10341 5201 10393
rect 5253 10341 5279 10393
rect 5331 10341 6121 10393
rect 6173 10341 6199 10393
rect 6251 10341 7041 10393
rect 7093 10341 7119 10393
rect 7171 10373 7587 10393
rect 7643 10373 7669 10429
rect 7725 10373 7751 10429
rect 7807 10373 7833 10429
rect 7889 10373 7915 10429
rect 7971 10393 7997 10405
rect 8053 10393 8079 10405
rect 8135 10373 8161 10429
rect 8217 10373 8243 10429
rect 8299 10373 8325 10429
rect 8381 10373 8407 10429
rect 8463 10373 8489 10429
rect 8545 10373 8571 10429
rect 8627 10373 8653 10429
rect 8709 10373 8735 10429
rect 8791 10373 8817 10429
rect 8873 10405 8881 10429
rect 8955 10405 8959 10429
rect 8873 10393 8899 10405
rect 8955 10393 8981 10405
rect 8873 10373 8881 10393
rect 8955 10373 8959 10393
rect 9037 10373 9063 10429
rect 9119 10373 9145 10429
rect 9201 10373 9227 10429
rect 9283 10373 9308 10429
rect 9364 10373 9389 10429
rect 9445 10373 9470 10429
rect 9526 10373 9551 10429
rect 9607 10373 9632 10429
rect 9688 10373 9713 10429
rect 9769 10405 9801 10429
rect 9853 10405 9879 10457
rect 9931 10405 10721 10457
rect 10773 10405 10799 10457
rect 10851 10405 11641 10457
rect 11693 10405 11719 10457
rect 11771 10405 12561 10457
rect 12613 10405 12639 10457
rect 12691 10405 14858 10457
rect 9769 10393 14858 10405
rect 9769 10373 9801 10393
rect 7171 10349 7961 10373
rect 8013 10349 8039 10373
rect 8091 10349 8881 10373
rect 8933 10349 8959 10373
rect 9011 10349 9801 10373
rect 7171 10341 7587 10349
rect 3491 10329 7587 10341
rect 3491 10301 4281 10329
rect 3361 10286 4281 10301
rect 3413 10234 3439 10286
rect 3491 10277 4281 10286
rect 4333 10277 4359 10329
rect 4411 10277 5201 10329
rect 5253 10277 5279 10329
rect 5331 10277 6121 10329
rect 6173 10277 6199 10329
rect 6251 10277 7041 10329
rect 7093 10277 7119 10329
rect 7171 10293 7587 10329
rect 7643 10293 7669 10349
rect 7725 10293 7751 10349
rect 7807 10293 7833 10349
rect 7889 10293 7915 10349
rect 7971 10329 7997 10341
rect 8053 10329 8079 10341
rect 8135 10293 8161 10349
rect 8217 10293 8243 10349
rect 8299 10293 8325 10349
rect 8381 10293 8407 10349
rect 8463 10293 8489 10349
rect 8545 10293 8571 10349
rect 8627 10293 8653 10349
rect 8709 10293 8735 10349
rect 8791 10293 8817 10349
rect 8873 10341 8881 10349
rect 8955 10341 8959 10349
rect 8873 10329 8899 10341
rect 8955 10329 8981 10341
rect 8873 10293 8881 10329
rect 8955 10293 8959 10329
rect 9037 10293 9063 10349
rect 9119 10293 9145 10349
rect 9201 10293 9227 10349
rect 9283 10293 9308 10349
rect 9364 10293 9389 10349
rect 9445 10293 9470 10349
rect 9526 10293 9551 10349
rect 9607 10293 9632 10349
rect 9688 10293 9713 10349
rect 9769 10341 9801 10349
rect 9853 10341 9879 10393
rect 9931 10341 10721 10393
rect 10773 10341 10799 10393
rect 10851 10341 11641 10393
rect 11693 10341 11719 10393
rect 11771 10341 12561 10393
rect 12613 10341 12639 10393
rect 12691 10341 14858 10393
rect 9769 10329 14858 10341
rect 9769 10293 9801 10329
rect 7171 10277 7961 10293
rect 8013 10277 8039 10293
rect 8091 10277 8881 10293
rect 8933 10277 8959 10293
rect 9011 10277 9801 10293
rect 9853 10277 9879 10329
rect 9931 10277 10721 10329
rect 10773 10277 10799 10329
rect 10851 10277 11641 10329
rect 11693 10277 11719 10329
rect 11771 10277 12561 10329
rect 12613 10277 12639 10329
rect 12691 10277 14858 10329
rect 3491 10269 14858 10277
rect 3491 10264 7587 10269
rect 3491 10234 4281 10264
rect 3361 10219 4281 10234
rect 3413 10167 3439 10219
rect 3491 10212 4281 10219
rect 4333 10212 4359 10264
rect 4411 10212 5201 10264
rect 5253 10212 5279 10264
rect 5331 10212 6121 10264
rect 6173 10212 6199 10264
rect 6251 10212 7041 10264
rect 7093 10212 7119 10264
rect 7171 10213 7587 10264
rect 7643 10213 7669 10269
rect 7725 10213 7751 10269
rect 7807 10213 7833 10269
rect 7889 10213 7915 10269
rect 7971 10264 7997 10269
rect 8053 10264 8079 10269
rect 8135 10213 8161 10269
rect 8217 10213 8243 10269
rect 8299 10213 8325 10269
rect 8381 10213 8407 10269
rect 8463 10213 8489 10269
rect 8545 10213 8571 10269
rect 8627 10213 8653 10269
rect 8709 10213 8735 10269
rect 8791 10213 8817 10269
rect 8873 10264 8899 10269
rect 8955 10264 8981 10269
rect 8873 10213 8881 10264
rect 8955 10213 8959 10264
rect 9037 10213 9063 10269
rect 9119 10213 9145 10269
rect 9201 10213 9227 10269
rect 9283 10213 9308 10269
rect 9364 10213 9389 10269
rect 9445 10213 9470 10269
rect 9526 10213 9551 10269
rect 9607 10213 9632 10269
rect 9688 10213 9713 10269
rect 9769 10264 14858 10269
rect 9769 10213 9801 10264
rect 7171 10212 7961 10213
rect 8013 10212 8039 10213
rect 8091 10212 8881 10213
rect 8933 10212 8959 10213
rect 9011 10212 9801 10213
rect 9853 10212 9879 10264
rect 9931 10212 10721 10264
rect 10773 10212 10799 10264
rect 10851 10212 11641 10264
rect 11693 10212 11719 10264
rect 11771 10212 12561 10264
rect 12613 10212 12639 10264
rect 12691 10212 14858 10264
rect 3491 10199 14858 10212
rect 3491 10167 4281 10199
rect 3361 10152 4281 10167
rect 3413 10100 3439 10152
rect 3491 10147 4281 10152
rect 4333 10147 4359 10199
rect 4411 10147 5201 10199
rect 5253 10147 5279 10199
rect 5331 10147 6121 10199
rect 6173 10147 6199 10199
rect 6251 10147 7041 10199
rect 7093 10147 7119 10199
rect 7171 10189 7961 10199
rect 8013 10189 8039 10199
rect 8091 10189 8881 10199
rect 8933 10189 8959 10199
rect 9011 10189 9801 10199
rect 7171 10147 7587 10189
rect 3491 10134 7587 10147
rect 3491 10100 4281 10134
rect 3361 10085 4281 10100
rect 3413 10033 3439 10085
rect 3491 10082 4281 10085
rect 4333 10082 4359 10134
rect 4411 10082 5201 10134
rect 5253 10082 5279 10134
rect 5331 10082 6121 10134
rect 6173 10082 6199 10134
rect 6251 10082 7041 10134
rect 7093 10082 7119 10134
rect 7171 10133 7587 10134
rect 7643 10133 7669 10189
rect 7725 10133 7751 10189
rect 7807 10133 7833 10189
rect 7889 10133 7915 10189
rect 7971 10134 7997 10147
rect 8053 10134 8079 10147
rect 8135 10133 8161 10189
rect 8217 10133 8243 10189
rect 8299 10133 8325 10189
rect 8381 10133 8407 10189
rect 8463 10133 8489 10189
rect 8545 10133 8571 10189
rect 8627 10133 8653 10189
rect 8709 10133 8735 10189
rect 8791 10133 8817 10189
rect 8873 10147 8881 10189
rect 8955 10147 8959 10189
rect 8873 10134 8899 10147
rect 8955 10134 8981 10147
rect 8873 10133 8881 10134
rect 8955 10133 8959 10134
rect 9037 10133 9063 10189
rect 9119 10133 9145 10189
rect 9201 10133 9227 10189
rect 9283 10133 9308 10189
rect 9364 10133 9389 10189
rect 9445 10133 9470 10189
rect 9526 10133 9551 10189
rect 9607 10133 9632 10189
rect 9688 10133 9713 10189
rect 9769 10147 9801 10189
rect 9853 10147 9879 10199
rect 9931 10147 10721 10199
rect 10773 10147 10799 10199
rect 10851 10147 11641 10199
rect 11693 10147 11719 10199
rect 11771 10147 12561 10199
rect 12613 10147 12639 10199
rect 12691 10147 14858 10199
rect 9769 10134 14858 10147
rect 9769 10133 9801 10134
rect 7171 10109 7961 10133
rect 8013 10109 8039 10133
rect 8091 10109 8881 10133
rect 8933 10109 8959 10133
rect 9011 10109 9801 10133
rect 7171 10082 7587 10109
rect 3491 10069 7587 10082
rect 3491 10033 4281 10069
rect 3361 10018 4281 10033
rect 3413 9966 3439 10018
rect 3491 10017 4281 10018
rect 4333 10017 4359 10069
rect 4411 10017 5201 10069
rect 5253 10017 5279 10069
rect 5331 10017 6121 10069
rect 6173 10017 6199 10069
rect 6251 10017 7041 10069
rect 7093 10017 7119 10069
rect 7171 10053 7587 10069
rect 7643 10053 7669 10109
rect 7725 10053 7751 10109
rect 7807 10053 7833 10109
rect 7889 10053 7915 10109
rect 7971 10069 7997 10082
rect 8053 10069 8079 10082
rect 8135 10053 8161 10109
rect 8217 10053 8243 10109
rect 8299 10053 8325 10109
rect 8381 10053 8407 10109
rect 8463 10053 8489 10109
rect 8545 10053 8571 10109
rect 8627 10053 8653 10109
rect 8709 10053 8735 10109
rect 8791 10053 8817 10109
rect 8873 10082 8881 10109
rect 8955 10082 8959 10109
rect 8873 10069 8899 10082
rect 8955 10069 8981 10082
rect 8873 10053 8881 10069
rect 8955 10053 8959 10069
rect 9037 10053 9063 10109
rect 9119 10053 9145 10109
rect 9201 10053 9227 10109
rect 9283 10053 9308 10109
rect 9364 10053 9389 10109
rect 9445 10053 9470 10109
rect 9526 10053 9551 10109
rect 9607 10053 9632 10109
rect 9688 10053 9713 10109
rect 9769 10082 9801 10109
rect 9853 10082 9879 10134
rect 9931 10082 10721 10134
rect 10773 10082 10799 10134
rect 10851 10082 11641 10134
rect 11693 10082 11719 10134
rect 11771 10082 12561 10134
rect 12613 10082 12639 10134
rect 12691 10082 14858 10134
rect 9769 10069 14858 10082
rect 9769 10053 9801 10069
rect 7171 10029 7961 10053
rect 8013 10029 8039 10053
rect 8091 10029 8881 10053
rect 8933 10029 8959 10053
rect 9011 10029 9801 10053
rect 7171 10017 7587 10029
rect 3491 10004 7587 10017
rect 3491 9966 4281 10004
rect 3361 9952 4281 9966
rect 4333 9952 4359 10004
rect 4411 9952 5201 10004
rect 5253 9952 5279 10004
rect 5331 9952 6121 10004
rect 6173 9952 6199 10004
rect 6251 9952 7041 10004
rect 7093 9952 7119 10004
rect 7171 9973 7587 10004
rect 7643 9973 7669 10029
rect 7725 9973 7751 10029
rect 7807 9973 7833 10029
rect 7889 9973 7915 10029
rect 7971 10004 7997 10017
rect 8053 10004 8079 10017
rect 8135 9973 8161 10029
rect 8217 9973 8243 10029
rect 8299 9973 8325 10029
rect 8381 9973 8407 10029
rect 8463 9973 8489 10029
rect 8545 9973 8571 10029
rect 8627 9973 8653 10029
rect 8709 9973 8735 10029
rect 8791 9973 8817 10029
rect 8873 10017 8881 10029
rect 8955 10017 8959 10029
rect 8873 10004 8899 10017
rect 8955 10004 8981 10017
rect 8873 9973 8881 10004
rect 8955 9973 8959 10004
rect 9037 9973 9063 10029
rect 9119 9973 9145 10029
rect 9201 9973 9227 10029
rect 9283 9973 9308 10029
rect 9364 9973 9389 10029
rect 9445 9973 9470 10029
rect 9526 9973 9551 10029
rect 9607 9973 9632 10029
rect 9688 9973 9713 10029
rect 9769 10017 9801 10029
rect 9853 10017 9879 10069
rect 9931 10017 10721 10069
rect 10773 10017 10799 10069
rect 10851 10017 11641 10069
rect 11693 10017 11719 10069
rect 11771 10017 12561 10069
rect 12613 10017 12639 10069
rect 12691 10017 14858 10069
rect 9769 10004 14858 10017
rect 9769 9973 9801 10004
rect 7171 9952 7961 9973
rect 8013 9952 8039 9973
rect 8091 9952 8881 9973
rect 8933 9952 8959 9973
rect 9011 9952 9801 9973
rect 9853 9952 9879 10004
rect 9931 9952 10721 10004
rect 10773 9952 10799 10004
rect 10851 9952 11641 10004
rect 11693 9952 11719 10004
rect 11771 9952 12561 10004
rect 12613 9952 12639 10004
rect 12691 9952 14858 10004
rect 3361 9951 14858 9952
rect 3413 9899 3439 9951
rect 3491 9949 14858 9951
rect 3491 9939 7587 9949
rect 3491 9899 4281 9939
rect 3361 9887 4281 9899
rect 4333 9887 4359 9939
rect 4411 9887 5201 9939
rect 5253 9887 5279 9939
rect 5331 9887 6121 9939
rect 6173 9887 6199 9939
rect 6251 9887 7041 9939
rect 7093 9887 7119 9939
rect 7171 9893 7587 9939
rect 7643 9893 7669 9949
rect 7725 9893 7751 9949
rect 7807 9893 7833 9949
rect 7889 9893 7915 9949
rect 7971 9939 7997 9949
rect 8053 9939 8079 9949
rect 8135 9893 8161 9949
rect 8217 9893 8243 9949
rect 8299 9893 8325 9949
rect 8381 9893 8407 9949
rect 8463 9893 8489 9949
rect 8545 9893 8571 9949
rect 8627 9893 8653 9949
rect 8709 9893 8735 9949
rect 8791 9893 8817 9949
rect 8873 9939 8899 9949
rect 8955 9939 8981 9949
rect 8873 9893 8881 9939
rect 8955 9893 8959 9939
rect 9037 9893 9063 9949
rect 9119 9893 9145 9949
rect 9201 9893 9227 9949
rect 9283 9893 9308 9949
rect 9364 9893 9389 9949
rect 9445 9893 9470 9949
rect 9526 9893 9551 9949
rect 9607 9893 9632 9949
rect 9688 9893 9713 9949
rect 9769 9939 14858 9949
rect 9769 9893 9801 9939
rect 7171 9887 7961 9893
rect 8013 9887 8039 9893
rect 8091 9887 8881 9893
rect 8933 9887 8959 9893
rect 9011 9887 9801 9893
rect 9853 9887 9879 9939
rect 9931 9887 10721 9939
rect 10773 9887 10799 9939
rect 10851 9887 11641 9939
rect 11693 9887 11719 9939
rect 11771 9887 12561 9939
rect 12613 9887 12639 9939
rect 12691 9887 14858 9939
rect 3361 9884 14858 9887
rect 3413 9832 3439 9884
rect 3491 9874 14858 9884
rect 3491 9832 4281 9874
rect 3361 9822 4281 9832
rect 4333 9822 4359 9874
rect 4411 9822 5201 9874
rect 5253 9822 5279 9874
rect 5331 9822 6121 9874
rect 6173 9822 6199 9874
rect 6251 9822 7041 9874
rect 7093 9822 7119 9874
rect 7171 9869 7961 9874
rect 8013 9869 8039 9874
rect 8091 9869 8881 9874
rect 8933 9869 8959 9874
rect 9011 9869 9801 9874
rect 7171 9822 7587 9869
rect 3361 9817 7587 9822
rect 3413 9765 3439 9817
rect 3491 9813 7587 9817
rect 7643 9813 7669 9869
rect 7725 9813 7751 9869
rect 7807 9813 7833 9869
rect 7889 9813 7915 9869
rect 7971 9813 7997 9822
rect 8053 9813 8079 9822
rect 8135 9813 8161 9869
rect 8217 9813 8243 9869
rect 8299 9813 8325 9869
rect 8381 9813 8407 9869
rect 8463 9813 8489 9869
rect 8545 9813 8571 9869
rect 8627 9813 8653 9869
rect 8709 9813 8735 9869
rect 8791 9813 8817 9869
rect 8873 9822 8881 9869
rect 8955 9822 8959 9869
rect 8873 9813 8899 9822
rect 8955 9813 8981 9822
rect 9037 9813 9063 9869
rect 9119 9813 9145 9869
rect 9201 9813 9227 9869
rect 9283 9813 9308 9869
rect 9364 9813 9389 9869
rect 9445 9813 9470 9869
rect 9526 9813 9551 9869
rect 9607 9813 9632 9869
rect 9688 9813 9713 9869
rect 9769 9822 9801 9869
rect 9853 9822 9879 9874
rect 9931 9822 10721 9874
rect 10773 9822 10799 9874
rect 10851 9822 11641 9874
rect 11693 9822 11719 9874
rect 11771 9822 12561 9874
rect 12613 9822 12639 9874
rect 12691 9822 14858 9874
rect 9769 9813 14858 9822
rect 3491 9809 14858 9813
rect 3491 9765 4281 9809
rect 3361 9757 4281 9765
rect 4333 9757 4359 9809
rect 4411 9757 5201 9809
rect 5253 9757 5279 9809
rect 5331 9757 6121 9809
rect 6173 9757 6199 9809
rect 6251 9757 7041 9809
rect 7093 9757 7119 9809
rect 7171 9789 7961 9809
rect 8013 9789 8039 9809
rect 8091 9789 8881 9809
rect 8933 9789 8959 9809
rect 9011 9789 9801 9809
rect 7171 9757 7587 9789
rect 3361 9750 7587 9757
rect 3413 9698 3439 9750
rect 3491 9744 7587 9750
rect 3491 9698 4281 9744
rect 3361 9692 4281 9698
rect 4333 9692 4359 9744
rect 4411 9692 5201 9744
rect 5253 9692 5279 9744
rect 5331 9692 6121 9744
rect 6173 9692 6199 9744
rect 6251 9692 7041 9744
rect 7093 9692 7119 9744
rect 7171 9733 7587 9744
rect 7643 9733 7669 9789
rect 7725 9733 7751 9789
rect 7807 9733 7833 9789
rect 7889 9733 7915 9789
rect 7971 9744 7997 9757
rect 8053 9744 8079 9757
rect 8135 9733 8161 9789
rect 8217 9733 8243 9789
rect 8299 9733 8325 9789
rect 8381 9733 8407 9789
rect 8463 9733 8489 9789
rect 8545 9733 8571 9789
rect 8627 9733 8653 9789
rect 8709 9733 8735 9789
rect 8791 9733 8817 9789
rect 8873 9757 8881 9789
rect 8955 9757 8959 9789
rect 8873 9744 8899 9757
rect 8955 9744 8981 9757
rect 8873 9733 8881 9744
rect 8955 9733 8959 9744
rect 9037 9733 9063 9789
rect 9119 9733 9145 9789
rect 9201 9733 9227 9789
rect 9283 9733 9308 9789
rect 9364 9733 9389 9789
rect 9445 9733 9470 9789
rect 9526 9733 9551 9789
rect 9607 9733 9632 9789
rect 9688 9733 9713 9789
rect 9769 9757 9801 9789
rect 9853 9757 9879 9809
rect 9931 9757 10721 9809
rect 10773 9757 10799 9809
rect 10851 9757 11641 9809
rect 11693 9757 11719 9809
rect 11771 9757 12561 9809
rect 12613 9757 12639 9809
rect 12691 9757 14858 9809
rect 9769 9744 14858 9757
rect 9769 9733 9801 9744
rect 7171 9709 7961 9733
rect 8013 9709 8039 9733
rect 8091 9709 8881 9733
rect 8933 9709 8959 9733
rect 9011 9709 9801 9733
rect 7171 9692 7587 9709
rect 3361 9683 7587 9692
rect 3413 9631 3439 9683
rect 3491 9679 7587 9683
rect 3491 9631 4281 9679
rect 3361 9627 4281 9631
rect 4333 9627 4359 9679
rect 4411 9627 5201 9679
rect 5253 9627 5279 9679
rect 5331 9627 6121 9679
rect 6173 9627 6199 9679
rect 6251 9627 7041 9679
rect 7093 9627 7119 9679
rect 7171 9653 7587 9679
rect 7643 9653 7669 9709
rect 7725 9653 7751 9709
rect 7807 9653 7833 9709
rect 7889 9653 7915 9709
rect 7971 9679 7997 9692
rect 8053 9679 8079 9692
rect 8135 9653 8161 9709
rect 8217 9653 8243 9709
rect 8299 9653 8325 9709
rect 8381 9653 8407 9709
rect 8463 9653 8489 9709
rect 8545 9653 8571 9709
rect 8627 9653 8653 9709
rect 8709 9653 8735 9709
rect 8791 9653 8817 9709
rect 8873 9692 8881 9709
rect 8955 9692 8959 9709
rect 8873 9679 8899 9692
rect 8955 9679 8981 9692
rect 8873 9653 8881 9679
rect 8955 9653 8959 9679
rect 9037 9653 9063 9709
rect 9119 9653 9145 9709
rect 9201 9653 9227 9709
rect 9283 9653 9308 9709
rect 9364 9653 9389 9709
rect 9445 9653 9470 9709
rect 9526 9653 9551 9709
rect 9607 9653 9632 9709
rect 9688 9653 9713 9709
rect 9769 9692 9801 9709
rect 9853 9692 9879 9744
rect 9931 9692 10721 9744
rect 10773 9692 10799 9744
rect 10851 9692 11641 9744
rect 11693 9692 11719 9744
rect 11771 9692 12561 9744
rect 12613 9692 12639 9744
rect 12691 9692 14858 9744
rect 9769 9679 14858 9692
rect 9769 9653 9801 9679
rect 7171 9629 7961 9653
rect 8013 9629 8039 9653
rect 8091 9629 8881 9653
rect 8933 9629 8959 9653
rect 9011 9629 9801 9653
rect 7171 9627 7587 9629
rect 3361 9616 7587 9627
rect 3413 9564 3439 9616
rect 3491 9614 7587 9616
rect 3491 9564 4281 9614
rect 3361 9562 4281 9564
rect 4333 9562 4359 9614
rect 4411 9562 5201 9614
rect 5253 9562 5279 9614
rect 5331 9562 6121 9614
rect 6173 9562 6199 9614
rect 6251 9562 7041 9614
rect 7093 9562 7119 9614
rect 7171 9573 7587 9614
rect 7643 9573 7669 9629
rect 7725 9573 7751 9629
rect 7807 9573 7833 9629
rect 7889 9573 7915 9629
rect 7971 9614 7997 9627
rect 8053 9614 8079 9627
rect 8135 9573 8161 9629
rect 8217 9573 8243 9629
rect 8299 9573 8325 9629
rect 8381 9573 8407 9629
rect 8463 9573 8489 9629
rect 8545 9573 8571 9629
rect 8627 9573 8653 9629
rect 8709 9573 8735 9629
rect 8791 9573 8817 9629
rect 8873 9627 8881 9629
rect 8955 9627 8959 9629
rect 8873 9614 8899 9627
rect 8955 9614 8981 9627
rect 8873 9573 8881 9614
rect 8955 9573 8959 9614
rect 9037 9573 9063 9629
rect 9119 9573 9145 9629
rect 9201 9573 9227 9629
rect 9283 9573 9308 9629
rect 9364 9573 9389 9629
rect 9445 9573 9470 9629
rect 9526 9573 9551 9629
rect 9607 9573 9632 9629
rect 9688 9573 9713 9629
rect 9769 9627 9801 9629
rect 9853 9627 9879 9679
rect 9931 9627 10721 9679
rect 10773 9627 10799 9679
rect 10851 9627 11641 9679
rect 11693 9627 11719 9679
rect 11771 9627 12561 9679
rect 12613 9627 12639 9679
rect 12691 9627 14858 9679
rect 9769 9614 14858 9627
rect 9769 9573 9801 9614
rect 7171 9562 7961 9573
rect 8013 9562 8039 9573
rect 8091 9562 8881 9573
rect 8933 9562 8959 9573
rect 9011 9562 9801 9573
rect 9853 9562 9879 9614
rect 9931 9562 10721 9614
rect 10773 9562 10799 9614
rect 10851 9562 11641 9614
rect 11693 9562 11719 9614
rect 11771 9562 12561 9614
rect 12613 9562 12639 9614
rect 12691 9562 14858 9614
rect 3361 9549 14858 9562
rect 3413 9497 3439 9549
rect 3491 9497 4281 9549
rect 4333 9497 4359 9549
rect 4411 9497 5201 9549
rect 5253 9497 5279 9549
rect 5331 9497 6121 9549
rect 6173 9497 6199 9549
rect 6251 9497 7041 9549
rect 7093 9497 7119 9549
rect 7171 9497 7587 9549
rect 3361 9493 7587 9497
rect 7643 9493 7669 9549
rect 7725 9493 7751 9549
rect 7807 9493 7833 9549
rect 7889 9493 7915 9549
rect 7971 9493 7997 9497
rect 8053 9493 8079 9497
rect 8135 9493 8161 9549
rect 8217 9493 8243 9549
rect 8299 9493 8325 9549
rect 8381 9493 8407 9549
rect 8463 9493 8489 9549
rect 8545 9493 8571 9549
rect 8627 9493 8653 9549
rect 8709 9493 8735 9549
rect 8791 9493 8817 9549
rect 8873 9497 8881 9549
rect 8955 9497 8959 9549
rect 8873 9493 8899 9497
rect 8955 9493 8981 9497
rect 9037 9493 9063 9549
rect 9119 9493 9145 9549
rect 9201 9493 9227 9549
rect 9283 9493 9308 9549
rect 9364 9493 9389 9549
rect 9445 9493 9470 9549
rect 9526 9493 9551 9549
rect 9607 9493 9632 9549
rect 9688 9493 9713 9549
rect 9769 9497 9801 9549
rect 9853 9497 9879 9549
rect 9931 9497 10721 9549
rect 10773 9497 10799 9549
rect 10851 9497 11641 9549
rect 11693 9497 11719 9549
rect 11771 9497 12561 9549
rect 12613 9497 12639 9549
rect 12691 9497 14858 9549
rect 9769 9493 14858 9497
rect 3361 9491 14858 9493
rect 187 9430 2233 9482
rect 2285 9430 2335 9482
rect 2387 9430 2824 9482
rect 187 9417 2824 9430
rect 187 9365 2233 9417
rect 2285 9365 2335 9417
rect 2387 9365 2824 9417
rect 187 9352 2824 9365
rect 187 9300 2233 9352
rect 2285 9300 2335 9352
rect 2387 9300 2824 9352
rect 187 9287 2824 9300
rect 187 9235 2233 9287
rect 2285 9235 2335 9287
rect 2387 9235 2824 9287
rect 187 9222 2824 9235
rect 187 9170 2233 9222
rect 2285 9170 2335 9222
rect 2387 9170 2824 9222
rect 187 9157 2824 9170
rect 187 9105 2233 9157
rect 2285 9105 2335 9157
rect 2387 9105 2824 9157
rect 187 8476 2824 9105
tri 2824 8476 3411 9063 sw
tri 11495 9016 11970 9491 ne
rect 11970 9016 14858 9491
rect 11191 8881 11964 8887
rect 11191 8829 11204 8881
rect 11256 8829 11274 8881
rect 11326 8829 11344 8881
rect 11396 8829 11414 8881
rect 11466 8829 11483 8881
rect 11535 8829 11552 8881
rect 11604 8829 11621 8881
rect 11673 8829 11690 8881
rect 11742 8829 11759 8881
rect 11811 8829 11828 8881
rect 11880 8829 11897 8881
rect 11949 8829 11964 8881
rect 11191 8759 11964 8829
tri 11970 8764 12222 9016 ne
rect 11191 8707 11204 8759
rect 11256 8707 11274 8759
rect 11326 8707 11344 8759
rect 11396 8707 11414 8759
rect 11466 8707 11483 8759
rect 11535 8707 11552 8759
rect 11604 8707 11621 8759
rect 11673 8707 11690 8759
rect 11742 8707 11759 8759
rect 11811 8707 11828 8759
rect 11880 8707 11897 8759
rect 11949 8707 11964 8759
rect 11191 8495 11964 8707
rect 187 8314 10840 8476
tri 10840 8314 11002 8476 sw
rect 11191 8443 11204 8495
rect 11256 8443 11274 8495
rect 11326 8443 11344 8495
rect 11396 8443 11414 8495
rect 11466 8443 11483 8495
rect 11535 8443 11552 8495
rect 11604 8443 11621 8495
rect 11673 8443 11690 8495
rect 11742 8443 11759 8495
rect 11811 8443 11828 8495
rect 11880 8443 11897 8495
rect 11949 8443 11964 8495
rect 11191 8373 11964 8443
rect 11191 8321 11204 8373
rect 11256 8321 11274 8373
rect 11326 8321 11344 8373
rect 11396 8321 11414 8373
rect 11466 8321 11483 8373
rect 11535 8321 11552 8373
rect 11604 8321 11621 8373
rect 11673 8321 11690 8373
rect 11742 8321 11759 8373
rect 11811 8321 11828 8373
rect 11880 8321 11897 8373
rect 11949 8321 11964 8373
rect 11191 8314 11964 8321
rect 187 8070 11002 8314
rect 187 8057 3965 8070
tri 3965 8057 3978 8070 nw
tri 10515 8059 10526 8070 ne
rect 10526 8059 11002 8070
rect 187 8043 3951 8057
tri 3951 8043 3965 8057 nw
tri 10526 8045 10540 8059 ne
rect 10540 8045 11002 8059
rect 187 8029 3937 8043
tri 3937 8029 3951 8043 nw
rect 187 8015 3923 8029
tri 3923 8015 3937 8029 nw
rect 187 8001 3909 8015
tri 3909 8001 3923 8015 nw
rect 187 7987 3895 8001
tri 3895 7987 3909 8001 nw
rect 187 7973 3881 7987
tri 3881 7973 3895 7987 nw
rect 187 7959 3867 7973
tri 3867 7959 3881 7973 nw
rect 187 7945 3853 7959
tri 3853 7945 3867 7959 nw
rect 187 7931 3839 7945
tri 3839 7931 3853 7945 nw
tri 10540 7933 10652 8045 ne
rect 10652 7933 11002 8045
tri 11002 7933 11383 8314 sw
rect 187 7917 3825 7931
tri 3825 7917 3839 7931 nw
rect 187 7914 3811 7917
rect 187 7862 695 7914
rect 747 7862 761 7914
rect 813 7862 827 7914
rect 879 7862 893 7914
rect 945 7862 959 7914
rect 1011 7862 1025 7914
rect 1077 7862 1091 7914
rect 1143 7862 1157 7914
rect 1209 7862 1223 7914
rect 1275 7862 1289 7914
rect 1341 7862 1355 7914
rect 1407 7862 1421 7914
rect 1473 7862 1487 7914
rect 1539 7862 1553 7914
rect 1605 7862 1619 7914
rect 1671 7862 1684 7914
rect 1736 7862 1749 7914
rect 1801 7862 1814 7914
rect 1866 7862 1879 7914
rect 1931 7862 1944 7914
rect 1996 7862 2009 7914
rect 2061 7862 2074 7914
rect 2126 7862 2139 7914
rect 2191 7862 2204 7914
rect 2256 7862 2269 7914
rect 2321 7862 2334 7914
rect 2386 7862 2399 7914
rect 2451 7862 2464 7914
rect 2516 7862 2529 7914
rect 2581 7862 2594 7914
rect 2646 7862 2659 7914
rect 2711 7862 2724 7914
rect 2776 7862 2789 7914
rect 2841 7862 2854 7914
rect 2906 7862 2919 7914
rect 2971 7862 2984 7914
rect 3036 7862 3049 7914
rect 3101 7862 3114 7914
rect 3166 7862 3179 7914
rect 3231 7862 3244 7914
rect 3296 7862 3309 7914
rect 3361 7862 3374 7914
rect 3426 7862 3439 7914
rect 3491 7862 3504 7914
rect 3556 7862 3569 7914
rect 3621 7903 3811 7914
tri 3811 7903 3825 7917 nw
rect 3621 7889 3797 7903
tri 3797 7889 3811 7903 nw
rect 3621 7875 3783 7889
tri 3783 7875 3797 7889 nw
rect 3621 7862 3769 7875
rect 187 7861 3769 7862
tri 3769 7861 3783 7875 nw
rect 187 7850 3755 7861
rect 187 7798 631 7850
rect 683 7847 3755 7850
tri 3755 7847 3769 7861 nw
rect 683 7833 3741 7847
tri 3741 7833 3755 7847 nw
tri 10652 7833 10752 7933 ne
rect 10752 7864 11383 7933
rect 10752 7833 10934 7864
rect 683 7819 3727 7833
tri 3727 7819 3741 7833 nw
rect 683 7805 3713 7819
tri 3713 7805 3727 7819 nw
rect 683 7798 3699 7805
rect 187 7796 3699 7798
rect 187 7786 749 7796
rect 187 7734 631 7786
rect 683 7744 749 7786
rect 801 7744 814 7796
rect 866 7744 879 7796
rect 931 7744 944 7796
rect 996 7744 1009 7796
rect 1061 7744 1073 7796
rect 1125 7744 1137 7796
rect 1189 7744 1201 7796
rect 1253 7744 1265 7796
rect 1317 7744 1329 7796
rect 1381 7744 1393 7796
rect 1445 7744 1457 7796
rect 1509 7744 1521 7796
rect 1573 7744 1585 7796
rect 1637 7744 1649 7796
rect 1701 7744 1713 7796
rect 1765 7744 1777 7796
rect 1829 7744 1841 7796
rect 1893 7744 1905 7796
rect 1957 7744 1969 7796
rect 2021 7744 2033 7796
rect 2085 7744 2097 7796
rect 2149 7744 2161 7796
rect 2213 7744 2225 7796
rect 2277 7744 2289 7796
rect 2341 7744 2353 7796
rect 2405 7744 2417 7796
rect 2469 7744 2481 7796
rect 2533 7744 2545 7796
rect 2597 7744 2609 7796
rect 2661 7744 2673 7796
rect 2725 7744 2737 7796
rect 2789 7744 2801 7796
rect 2853 7744 2865 7796
rect 2917 7744 2929 7796
rect 2981 7744 2993 7796
rect 3045 7744 3057 7796
rect 3109 7744 3121 7796
rect 3173 7744 3185 7796
rect 3237 7744 3249 7796
rect 3301 7744 3313 7796
rect 3365 7744 3377 7796
rect 3429 7744 3441 7796
rect 3493 7744 3505 7796
rect 3557 7744 3569 7796
rect 3621 7791 3699 7796
tri 3699 7791 3713 7805 nw
rect 3621 7777 3685 7791
tri 3685 7777 3699 7791 nw
rect 3621 7763 3671 7777
tri 3671 7763 3685 7777 nw
rect 3621 7744 3652 7763
tri 3652 7744 3671 7763 nw
rect 9727 7750 10729 7756
rect 683 7735 3643 7744
tri 3643 7735 3652 7744 nw
rect 683 7734 3629 7735
rect 187 7732 3629 7734
rect 187 7722 749 7732
rect 187 7670 631 7722
rect 683 7680 749 7722
rect 801 7721 3629 7732
tri 3629 7721 3643 7735 nw
rect 801 7707 3615 7721
tri 3615 7707 3629 7721 nw
rect 801 7693 3601 7707
tri 3601 7693 3615 7707 nw
rect 9727 7704 10677 7750
rect 9727 7698 9807 7704
tri 9807 7698 9813 7704 nw
tri 10646 7698 10652 7704 ne
rect 10652 7698 10677 7704
rect 801 7680 3587 7693
rect 683 7679 3587 7680
tri 3587 7679 3601 7693 nw
rect 9727 7686 9795 7698
tri 9795 7686 9807 7698 nw
tri 10652 7686 10664 7698 ne
rect 10664 7686 10729 7698
rect 683 7670 3573 7679
rect 187 7668 3573 7670
rect 187 7658 749 7668
rect 187 7606 631 7658
rect 683 7616 749 7658
rect 801 7665 3573 7668
tri 3573 7665 3587 7679 nw
rect 801 7651 3559 7665
tri 3559 7651 3573 7665 nw
rect 801 7637 3545 7651
tri 3545 7637 3559 7651 nw
rect 801 7623 3531 7637
tri 3531 7623 3545 7637 nw
rect 801 7616 3517 7623
rect 683 7609 3517 7616
tri 3517 7609 3531 7623 nw
rect 683 7606 3503 7609
rect 187 7604 3503 7606
rect 187 7594 749 7604
rect 187 7542 631 7594
rect 683 7552 749 7594
rect 801 7595 3503 7604
tri 3503 7595 3517 7609 nw
rect 801 7581 3489 7595
tri 3489 7581 3503 7595 nw
rect 801 7567 3475 7581
tri 3475 7567 3489 7581 nw
rect 801 7553 3461 7567
tri 3461 7553 3475 7567 nw
rect 801 7552 3447 7553
rect 683 7542 3447 7552
rect 187 7540 3447 7542
rect 187 7530 749 7540
rect 187 7478 631 7530
rect 683 7488 749 7530
rect 801 7539 3447 7540
tri 3447 7539 3461 7553 nw
rect 801 7525 3433 7539
tri 3433 7525 3447 7539 nw
rect 801 7511 3419 7525
tri 3419 7511 3433 7525 nw
rect 801 7497 3405 7511
tri 3405 7497 3419 7511 nw
rect 801 7488 3391 7497
rect 683 7483 3391 7488
tri 3391 7483 3405 7497 nw
rect 683 7478 3377 7483
rect 187 7476 3377 7478
rect 187 7466 749 7476
rect 187 7414 631 7466
rect 683 7424 749 7466
rect 801 7469 3377 7476
tri 3377 7469 3391 7483 nw
rect 801 7455 3363 7469
tri 3363 7455 3377 7469 nw
tri 9714 7455 9727 7468 se
rect 9727 7455 9779 7686
tri 9779 7670 9795 7686 nw
tri 10664 7673 10677 7686 ne
tri 10752 7651 10934 7833 ne
rect 10986 7812 11000 7864
rect 11052 7812 11066 7864
rect 11118 7812 11132 7864
rect 11184 7812 11198 7864
rect 11250 7812 11264 7864
rect 11316 7812 11330 7864
rect 11382 7812 11383 7864
rect 10934 7793 11383 7812
rect 10986 7741 11000 7793
rect 11052 7741 11066 7793
rect 11118 7741 11132 7793
rect 11184 7741 11198 7793
rect 11250 7741 11264 7793
rect 11316 7741 11330 7793
rect 11382 7741 11383 7793
rect 10934 7722 11383 7741
rect 10986 7670 11000 7722
rect 11052 7670 11066 7722
rect 11118 7670 11132 7722
rect 11184 7670 11198 7722
rect 11250 7670 11264 7722
rect 11316 7670 11330 7722
rect 11382 7670 11383 7722
rect 10934 7651 11383 7670
rect 10677 7628 10729 7634
rect 801 7441 3349 7455
tri 3349 7441 3363 7455 nw
rect 801 7427 3335 7441
tri 3335 7427 3349 7441 nw
tri 9694 7435 9714 7455 se
rect 9714 7435 9779 7455
tri 9693 7434 9694 7435 se
rect 9694 7434 9779 7435
rect 801 7424 3321 7427
rect 683 7414 3321 7424
rect 187 7413 3321 7414
tri 3321 7413 3335 7427 nw
rect 187 7412 3307 7413
rect 187 7402 749 7412
rect 187 7350 631 7402
rect 683 7360 749 7402
rect 801 7399 3307 7412
tri 3307 7399 3321 7413 nw
rect 801 7385 3293 7399
tri 3293 7385 3307 7399 nw
rect 801 7371 3279 7385
tri 3279 7371 3293 7385 nw
rect 8889 7382 8895 7434
rect 8947 7382 8959 7434
rect 9011 7382 9779 7434
rect 10986 7599 11000 7651
rect 11052 7599 11066 7651
rect 11118 7599 11132 7651
rect 11184 7599 11198 7651
rect 11250 7599 11264 7651
rect 11316 7599 11330 7651
rect 11382 7599 11383 7651
rect 10934 7579 11383 7599
rect 10986 7527 11000 7579
rect 11052 7527 11066 7579
rect 11118 7527 11132 7579
rect 11184 7527 11198 7579
rect 11250 7527 11264 7579
rect 11316 7527 11330 7579
rect 11382 7527 11383 7579
rect 10934 7507 11383 7527
rect 10986 7455 11000 7507
rect 11052 7455 11066 7507
rect 11118 7455 11132 7507
rect 11184 7455 11198 7507
rect 11250 7455 11264 7507
rect 11316 7455 11330 7507
rect 11382 7455 11383 7507
rect 10934 7435 11383 7455
rect 10986 7383 11000 7435
rect 11052 7383 11066 7435
rect 11118 7383 11132 7435
rect 11184 7383 11198 7435
rect 11250 7383 11264 7435
rect 11316 7383 11330 7435
rect 11382 7383 11383 7435
rect 801 7360 3265 7371
rect 683 7357 3265 7360
tri 3265 7357 3279 7371 nw
rect 10934 7363 11383 7383
rect 683 7350 3251 7357
rect 187 7348 3251 7350
rect 187 7338 749 7348
rect 187 7286 631 7338
rect 683 7296 749 7338
rect 801 7343 3251 7348
tri 3251 7343 3265 7357 nw
rect 801 7329 3237 7343
tri 3237 7329 3251 7343 nw
rect 801 7315 3223 7329
tri 3223 7315 3237 7329 nw
rect 801 7301 3209 7315
tri 3209 7301 3223 7315 nw
rect 10986 7311 11000 7363
rect 11052 7311 11066 7363
rect 11118 7311 11132 7363
rect 11184 7311 11198 7363
rect 11250 7311 11264 7363
rect 11316 7311 11330 7363
rect 11382 7311 11383 7363
rect 801 7296 3195 7301
rect 683 7287 3195 7296
tri 3195 7287 3209 7301 nw
rect 3440 7296 9112 7297
rect 3440 7295 7588 7296
rect 7644 7295 7670 7296
rect 7726 7295 7751 7296
rect 7807 7295 7832 7296
rect 7888 7295 7913 7296
rect 7969 7295 7994 7296
rect 8050 7295 8075 7296
rect 8131 7295 8156 7296
rect 8212 7295 8237 7296
rect 8293 7295 8318 7296
rect 8374 7295 8399 7296
rect 8455 7295 8480 7296
rect 8536 7295 8561 7296
rect 8617 7295 8642 7296
rect 8698 7295 8723 7296
rect 8779 7295 8804 7296
rect 8860 7295 8885 7296
rect 8941 7295 8966 7296
rect 9022 7295 9047 7296
rect 683 7286 3181 7287
rect 187 7283 3181 7286
rect 187 7274 749 7283
rect 187 7222 631 7274
rect 683 7231 749 7274
rect 801 7273 3181 7283
tri 3181 7273 3195 7287 nw
rect 801 7259 3167 7273
tri 3167 7259 3181 7273 nw
rect 801 7245 3153 7259
tri 3153 7245 3167 7259 nw
rect 801 7231 3139 7245
tri 3139 7231 3153 7245 nw
rect 3440 7243 3446 7295
rect 3498 7243 3511 7295
rect 3563 7243 3576 7295
rect 3628 7243 3641 7295
rect 3693 7243 3706 7295
rect 3758 7243 3771 7295
rect 3823 7243 3836 7295
rect 3888 7243 3901 7295
rect 3953 7243 3966 7295
rect 4018 7243 4031 7295
rect 4083 7243 4096 7295
rect 4148 7243 4161 7295
rect 4213 7243 4226 7295
rect 4278 7243 4291 7295
rect 4343 7243 4356 7295
rect 4408 7243 4421 7295
rect 4473 7243 4486 7295
rect 4538 7243 4551 7295
rect 4603 7243 4616 7295
rect 4668 7243 4681 7295
rect 4733 7243 4746 7295
rect 4798 7243 4811 7295
rect 4863 7243 4876 7295
rect 4928 7243 4941 7295
rect 4993 7243 5006 7295
rect 5058 7243 5071 7295
rect 5123 7243 5136 7295
rect 5188 7243 5201 7295
rect 5253 7243 5266 7295
rect 5318 7243 5331 7295
rect 5383 7243 5396 7295
rect 5448 7243 5461 7295
rect 5513 7243 5526 7295
rect 5578 7243 5591 7295
rect 3440 7231 5591 7243
rect 9103 7240 9112 7296
rect 683 7222 3125 7231
rect 187 7218 3125 7222
rect 187 7210 749 7218
rect 187 7158 631 7210
rect 683 7166 749 7210
rect 801 7217 3125 7218
tri 3125 7217 3139 7231 nw
rect 801 7203 3111 7217
tri 3111 7203 3125 7217 nw
rect 801 7189 3097 7203
tri 3097 7189 3111 7203 nw
rect 801 7175 3083 7189
tri 3083 7175 3097 7189 nw
rect 3440 7179 3446 7231
rect 3498 7179 3511 7231
rect 3563 7179 3576 7231
rect 3628 7179 3641 7231
rect 3693 7179 3706 7231
rect 3758 7179 3771 7231
rect 3823 7179 3836 7231
rect 3888 7179 3901 7231
rect 3953 7179 3966 7231
rect 4018 7179 4031 7231
rect 4083 7179 4096 7231
rect 4148 7179 4161 7231
rect 4213 7179 4226 7231
rect 4278 7179 4291 7231
rect 4343 7179 4356 7231
rect 4408 7179 4421 7231
rect 4473 7179 4486 7231
rect 4538 7179 4551 7231
rect 4603 7179 4616 7231
rect 4668 7179 4681 7231
rect 4733 7179 4746 7231
rect 4798 7179 4811 7231
rect 4863 7179 4876 7231
rect 4928 7179 4941 7231
rect 4993 7179 5006 7231
rect 5058 7179 5071 7231
rect 5123 7179 5136 7231
rect 5188 7179 5201 7231
rect 5253 7179 5266 7231
rect 5318 7179 5331 7231
rect 5383 7179 5396 7231
rect 5448 7179 5461 7231
rect 5513 7179 5526 7231
rect 5578 7179 5591 7231
rect 9099 7214 9112 7240
rect 10934 7291 11383 7311
rect 10986 7239 11000 7291
rect 11052 7239 11066 7291
rect 11118 7239 11132 7291
rect 11184 7239 11198 7291
rect 11250 7239 11264 7291
rect 11316 7239 11330 7291
rect 11382 7239 11383 7291
rect 10934 7223 11383 7239
rect 801 7166 3069 7175
rect 683 7161 3069 7166
tri 3069 7161 3083 7175 nw
rect 3440 7167 5591 7179
rect 683 7158 3041 7161
rect 187 7153 3041 7158
rect 187 7146 749 7153
rect 187 7094 631 7146
rect 683 7101 749 7146
rect 801 7101 3041 7153
tri 3041 7133 3069 7161 nw
rect 683 7094 3041 7101
rect 187 7088 3041 7094
rect 187 7082 749 7088
rect 187 7030 631 7082
rect 683 7036 749 7082
rect 801 7036 3041 7088
rect 683 7030 3041 7036
rect 187 7023 3041 7030
rect 187 7018 749 7023
rect 187 6966 631 7018
rect 683 6971 749 7018
rect 801 6971 3041 7023
rect 683 6966 3041 6971
rect 187 6958 3041 6966
rect 187 6954 749 6958
rect 187 6902 631 6954
rect 683 6906 749 6954
rect 801 6906 3041 6958
rect 683 6902 3041 6906
rect 187 6893 3041 6902
rect 187 6890 749 6893
rect 187 6838 631 6890
rect 683 6841 749 6890
rect 801 6841 3041 6893
rect 683 6838 3041 6841
rect 187 6828 3041 6838
rect 187 6826 749 6828
rect 187 6774 631 6826
rect 683 6776 749 6826
rect 801 6776 3041 6828
rect 683 6774 3041 6776
rect 187 6763 3041 6774
rect 187 6762 749 6763
rect 187 6710 631 6762
rect 683 6711 749 6762
rect 801 6711 3041 6763
rect 683 6710 3041 6711
rect 187 6698 3041 6710
rect 187 6646 631 6698
rect 683 6646 749 6698
rect 801 6646 3041 6698
rect 3440 7115 3446 7167
rect 3498 7115 3511 7167
rect 3563 7115 3576 7167
rect 3628 7115 3641 7167
rect 3693 7115 3706 7167
rect 3758 7115 3771 7167
rect 3823 7115 3836 7167
rect 3888 7115 3901 7167
rect 3953 7115 3966 7167
rect 4018 7115 4031 7167
rect 4083 7115 4096 7167
rect 4148 7115 4161 7167
rect 4213 7115 4226 7167
rect 4278 7115 4291 7167
rect 4343 7115 4356 7167
rect 4408 7115 4421 7167
rect 4473 7115 4486 7167
rect 4538 7115 4551 7167
rect 4603 7115 4616 7167
rect 4668 7115 4681 7167
rect 4733 7115 4746 7167
rect 4798 7115 4811 7167
rect 4863 7115 4876 7167
rect 4928 7115 4941 7167
rect 4993 7115 5006 7167
rect 5058 7115 5071 7167
rect 5123 7115 5136 7167
rect 5188 7115 5201 7167
rect 5253 7115 5266 7167
rect 5318 7115 5331 7167
rect 5383 7115 5396 7167
rect 5448 7115 5461 7167
rect 5513 7115 5526 7167
rect 5578 7115 5591 7167
rect 9103 7158 9112 7214
tri 9938 7160 9940 7162 se
rect 9940 7160 11164 7166
rect 9099 7132 9112 7158
rect 3440 7103 5591 7115
rect 3440 7051 3446 7103
rect 3498 7051 3511 7103
rect 3563 7051 3576 7103
rect 3628 7051 3641 7103
rect 3693 7051 3706 7103
rect 3758 7051 3771 7103
rect 3823 7051 3836 7103
rect 3888 7051 3901 7103
rect 3953 7051 3966 7103
rect 4018 7051 4031 7103
rect 4083 7051 4096 7103
rect 4148 7051 4161 7103
rect 4213 7051 4226 7103
rect 4278 7051 4291 7103
rect 4343 7051 4356 7103
rect 4408 7051 4421 7103
rect 4473 7051 4486 7103
rect 4538 7051 4551 7103
rect 4603 7051 4616 7103
rect 4668 7051 4681 7103
rect 4733 7051 4746 7103
rect 4798 7051 4811 7103
rect 4863 7051 4876 7103
rect 4928 7051 4941 7103
rect 4993 7051 5006 7103
rect 5058 7051 5071 7103
rect 5123 7051 5136 7103
rect 5188 7051 5201 7103
rect 5253 7051 5266 7103
rect 5318 7051 5331 7103
rect 5383 7051 5396 7103
rect 5448 7051 5461 7103
rect 5513 7051 5526 7103
rect 5578 7051 5591 7103
rect 9103 7076 9112 7132
tri 9886 7108 9938 7160 se
rect 9938 7108 10985 7160
rect 11037 7108 11111 7160
rect 11163 7108 11164 7160
tri 9873 7095 9886 7108 se
rect 9886 7095 11164 7108
rect 3440 7039 5591 7051
rect 9099 7050 9112 7076
rect 3440 6987 3446 7039
rect 3498 6987 3511 7039
rect 3563 6987 3576 7039
rect 3628 6987 3641 7039
rect 3693 6987 3706 7039
rect 3758 6987 3771 7039
rect 3823 6987 3836 7039
rect 3888 6987 3901 7039
rect 3953 6987 3966 7039
rect 4018 6987 4031 7039
rect 4083 6987 4096 7039
rect 4148 6987 4161 7039
rect 4213 6987 4226 7039
rect 4278 6987 4291 7039
rect 4343 6987 4356 7039
rect 4408 6987 4421 7039
rect 4473 6987 4486 7039
rect 4538 6987 4551 7039
rect 4603 6987 4616 7039
rect 4668 6987 4681 7039
rect 4733 6987 4746 7039
rect 4798 6987 4811 7039
rect 4863 6987 4876 7039
rect 4928 6987 4941 7039
rect 4993 6987 5006 7039
rect 5058 6987 5071 7039
rect 5123 6987 5136 7039
rect 5188 6987 5201 7039
rect 5253 6987 5266 7039
rect 5318 6987 5331 7039
rect 5383 6987 5396 7039
rect 5448 6987 5461 7039
rect 5513 6987 5526 7039
rect 5578 6987 5591 7039
rect 9103 6994 9112 7050
tri 9821 7043 9873 7095 se
rect 9873 7043 10985 7095
rect 11037 7043 11111 7095
rect 11163 7043 11164 7095
tri 9808 7030 9821 7043 se
rect 9821 7030 11164 7043
rect 3440 6975 5591 6987
rect 3440 6923 3446 6975
rect 3498 6923 3511 6975
rect 3563 6923 3576 6975
rect 3628 6923 3641 6975
rect 3693 6923 3706 6975
rect 3758 6923 3771 6975
rect 3823 6923 3836 6975
rect 3888 6923 3901 6975
rect 3953 6923 3966 6975
rect 4018 6923 4031 6975
rect 4083 6923 4096 6975
rect 4148 6923 4161 6975
rect 4213 6923 4226 6975
rect 4278 6923 4291 6975
rect 4343 6923 4356 6975
rect 4408 6923 4421 6975
rect 4473 6923 4486 6975
rect 4538 6923 4551 6975
rect 4603 6923 4616 6975
rect 4668 6923 4681 6975
rect 4733 6923 4746 6975
rect 4798 6923 4811 6975
rect 4863 6923 4876 6975
rect 4928 6923 4941 6975
rect 4993 6923 5006 6975
rect 5058 6923 5071 6975
rect 5123 6923 5136 6975
rect 5188 6923 5201 6975
rect 5253 6923 5266 6975
rect 5318 6923 5331 6975
rect 5383 6923 5396 6975
rect 5448 6923 5461 6975
rect 5513 6923 5526 6975
rect 5578 6923 5591 6975
rect 9099 6968 9112 6994
tri 9756 6978 9808 7030 se
rect 9808 6978 10985 7030
rect 11037 6978 11111 7030
rect 11163 6978 11164 7030
rect 3440 6911 5591 6923
rect 9103 6912 9112 6968
tri 9743 6965 9756 6978 se
rect 9756 6965 11164 6978
tri 9691 6913 9743 6965 se
rect 9743 6913 10985 6965
rect 11037 6913 11111 6965
rect 11163 6913 11164 6965
rect 3440 6859 3446 6911
rect 3498 6859 3511 6911
rect 3563 6859 3576 6911
rect 3628 6859 3641 6911
rect 3693 6859 3706 6911
rect 3758 6859 3771 6911
rect 3823 6859 3836 6911
rect 3888 6859 3901 6911
rect 3953 6859 3966 6911
rect 4018 6859 4031 6911
rect 4083 6859 4096 6911
rect 4148 6859 4161 6911
rect 4213 6859 4226 6911
rect 4278 6859 4291 6911
rect 4343 6859 4356 6911
rect 4408 6859 4421 6911
rect 4473 6859 4486 6911
rect 4538 6859 4551 6911
rect 4603 6859 4616 6911
rect 4668 6859 4681 6911
rect 4733 6859 4746 6911
rect 4798 6859 4811 6911
rect 4863 6859 4876 6911
rect 4928 6859 4941 6911
rect 4993 6859 5006 6911
rect 5058 6859 5071 6911
rect 5123 6859 5136 6911
rect 5188 6859 5201 6911
rect 5253 6859 5266 6911
rect 5318 6859 5331 6911
rect 5383 6859 5396 6911
rect 5448 6859 5461 6911
rect 5513 6859 5526 6911
rect 5578 6859 5591 6911
rect 9099 6886 9112 6912
tri 9677 6899 9691 6913 se
rect 9691 6899 11164 6913
rect 3440 6847 5591 6859
rect 3440 6795 3446 6847
rect 3498 6795 3511 6847
rect 3563 6795 3576 6847
rect 3628 6795 3641 6847
rect 3693 6795 3706 6847
rect 3758 6795 3771 6847
rect 3823 6795 3836 6847
rect 3888 6795 3901 6847
rect 3953 6795 3966 6847
rect 4018 6795 4031 6847
rect 4083 6795 4096 6847
rect 4148 6795 4161 6847
rect 4213 6795 4226 6847
rect 4278 6795 4291 6847
rect 4343 6795 4356 6847
rect 4408 6795 4421 6847
rect 4473 6795 4486 6847
rect 4538 6795 4551 6847
rect 4603 6795 4616 6847
rect 4668 6795 4681 6847
rect 4733 6795 4746 6847
rect 4798 6795 4811 6847
rect 4863 6795 4876 6847
rect 4928 6795 4941 6847
rect 4993 6795 5006 6847
rect 5058 6795 5071 6847
rect 5123 6795 5136 6847
rect 5188 6795 5201 6847
rect 5253 6795 5266 6847
rect 5318 6795 5331 6847
rect 5383 6795 5396 6847
rect 5448 6795 5461 6847
rect 5513 6795 5526 6847
rect 5578 6795 5591 6847
rect 9103 6830 9112 6886
tri 9625 6847 9677 6899 se
rect 9677 6847 10985 6899
rect 11037 6847 11111 6899
rect 11163 6847 11164 6899
tri 9611 6833 9625 6847 se
rect 9625 6833 11164 6847
rect 9099 6804 9112 6830
rect 3440 6783 5591 6795
rect 3440 6731 3446 6783
rect 3498 6731 3511 6783
rect 3563 6731 3576 6783
rect 3628 6731 3641 6783
rect 3693 6731 3706 6783
rect 3758 6731 3771 6783
rect 3823 6731 3836 6783
rect 3888 6731 3901 6783
rect 3953 6731 3966 6783
rect 4018 6731 4031 6783
rect 4083 6731 4096 6783
rect 4148 6731 4161 6783
rect 4213 6731 4226 6783
rect 4278 6731 4291 6783
rect 4343 6731 4356 6783
rect 4408 6731 4421 6783
rect 4473 6731 4486 6783
rect 4538 6731 4551 6783
rect 4603 6731 4616 6783
rect 4668 6731 4681 6783
rect 4733 6731 4746 6783
rect 4798 6731 4811 6783
rect 4863 6731 4876 6783
rect 4928 6731 4941 6783
rect 4993 6731 5006 6783
rect 5058 6731 5071 6783
rect 5123 6731 5136 6783
rect 5188 6731 5201 6783
rect 5253 6731 5266 6783
rect 5318 6731 5331 6783
rect 5383 6731 5396 6783
rect 5448 6731 5461 6783
rect 5513 6731 5526 6783
rect 5578 6731 5591 6783
rect 9103 6748 9112 6804
tri 9559 6781 9611 6833 se
rect 9611 6781 10985 6833
rect 11037 6781 11111 6833
rect 11163 6781 11164 6833
tri 9545 6767 9559 6781 se
rect 9559 6767 11164 6781
rect 3440 6719 5591 6731
rect 9099 6722 9112 6748
rect 3440 6667 3446 6719
rect 3498 6667 3511 6719
rect 3563 6667 3576 6719
rect 3628 6667 3641 6719
rect 3693 6667 3706 6719
rect 3758 6667 3771 6719
rect 3823 6667 3836 6719
rect 3888 6667 3901 6719
rect 3953 6667 3966 6719
rect 4018 6667 4031 6719
rect 4083 6667 4096 6719
rect 4148 6667 4161 6719
rect 4213 6667 4226 6719
rect 4278 6667 4291 6719
rect 4343 6667 4356 6719
rect 4408 6667 4421 6719
rect 4473 6667 4486 6719
rect 4538 6667 4551 6719
rect 4603 6667 4616 6719
rect 4668 6667 4681 6719
rect 4733 6667 4746 6719
rect 4798 6667 4811 6719
rect 4863 6667 4876 6719
rect 4928 6667 4941 6719
rect 4993 6667 5006 6719
rect 5058 6667 5071 6719
rect 5123 6667 5136 6719
rect 5188 6667 5201 6719
rect 5253 6667 5266 6719
rect 5318 6667 5331 6719
rect 5383 6667 5396 6719
rect 5448 6667 5461 6719
rect 5513 6667 5526 6719
rect 5578 6667 5591 6719
rect 3440 6666 7588 6667
rect 7644 6666 7670 6667
rect 7726 6666 7751 6667
rect 7807 6666 7832 6667
rect 7888 6666 7913 6667
rect 7969 6666 7994 6667
rect 8050 6666 8075 6667
rect 8131 6666 8156 6667
rect 8212 6666 8237 6667
rect 8293 6666 8318 6667
rect 8374 6666 8399 6667
rect 8455 6666 8480 6667
rect 8536 6666 8561 6667
rect 8617 6666 8642 6667
rect 8698 6666 8723 6667
rect 8779 6666 8804 6667
rect 8860 6666 8885 6667
rect 8941 6666 8966 6667
rect 9022 6666 9047 6667
rect 9103 6666 9112 6722
tri 9493 6715 9545 6767 se
rect 9545 6715 10985 6767
rect 11037 6715 11111 6767
rect 11163 6715 11164 6767
tri 9479 6701 9493 6715 se
rect 9493 6701 11164 6715
rect 3440 6665 9112 6666
tri 9443 6665 9479 6701 se
rect 9479 6665 10985 6701
tri 9427 6649 9443 6665 se
rect 9443 6649 10985 6665
rect 11037 6649 11111 6701
rect 11163 6649 11164 6701
rect 187 6634 3041 6646
tri 9413 6635 9427 6649 se
rect 9427 6635 11164 6649
rect 187 6582 631 6634
rect 683 6633 3041 6634
rect 683 6582 749 6633
rect 187 6581 749 6582
rect 801 6581 3041 6633
tri 9362 6584 9413 6635 se
rect 9413 6584 10985 6635
rect 187 6570 3041 6581
rect 187 6518 631 6570
rect 683 6568 3041 6570
rect 683 6518 749 6568
rect 187 6516 749 6518
rect 801 6516 3041 6568
rect 187 6506 3041 6516
rect 187 6454 631 6506
rect 683 6503 3041 6506
rect 683 6454 749 6503
rect 187 6451 749 6454
rect 801 6451 3041 6503
rect 187 6442 3041 6451
rect 187 6390 631 6442
rect 683 6438 3041 6442
rect 683 6390 749 6438
rect 187 6386 749 6390
rect 801 6386 3041 6438
rect 187 6378 3041 6386
rect 187 6326 631 6378
rect 683 6373 3041 6378
rect 683 6326 749 6373
rect 187 6321 749 6326
rect 801 6321 3041 6373
rect 187 6314 3041 6321
rect 187 6262 631 6314
rect 683 6308 3041 6314
rect 683 6262 749 6308
rect 187 6256 749 6262
rect 801 6256 3041 6308
rect 187 6250 3041 6256
rect 187 6198 631 6250
rect 683 6243 3041 6250
rect 683 6198 749 6243
rect 187 6191 749 6198
rect 801 6191 3041 6243
rect 187 6186 3041 6191
rect 187 6134 631 6186
rect 683 6178 3041 6186
rect 683 6134 749 6178
rect 187 6126 749 6134
rect 801 6126 3041 6178
rect 187 6122 3041 6126
rect 187 6070 631 6122
rect 683 6113 3041 6122
rect 683 6070 749 6113
rect 187 6061 749 6070
rect 801 6061 3041 6113
rect 187 6058 3041 6061
rect 187 6006 631 6058
rect 683 6048 3041 6058
rect 683 6006 749 6048
rect 187 5996 749 6006
rect 801 5996 3041 6048
rect 187 5994 3041 5996
rect 187 5942 631 5994
rect 683 5983 3041 5994
rect 683 5942 749 5983
rect 187 5931 749 5942
rect 801 5931 3041 5983
rect 187 5929 3041 5931
rect 187 5877 631 5929
rect 683 5918 3041 5929
rect 683 5877 749 5918
rect 187 5866 749 5877
rect 801 5866 3041 5918
rect 187 5864 3041 5866
rect 187 5812 631 5864
rect 683 5853 3041 5864
rect 3848 6570 4040 6584
rect 3848 6518 3857 6570
rect 3909 6518 3981 6570
rect 4033 6518 4040 6570
rect 3848 6500 4040 6518
rect 3848 6448 3857 6500
rect 3909 6448 3981 6500
rect 4033 6448 4040 6500
rect 3848 6430 4040 6448
rect 3848 6378 3857 6430
rect 3909 6378 3981 6430
rect 4033 6378 4040 6430
rect 3848 6359 4040 6378
rect 3848 6307 3857 6359
rect 3909 6307 3981 6359
rect 4033 6307 4040 6359
rect 3848 6288 4040 6307
rect 3848 6236 3857 6288
rect 3909 6236 3981 6288
rect 4033 6236 4040 6288
rect 3848 6217 4040 6236
rect 3848 6165 3857 6217
rect 3909 6165 3981 6217
rect 4033 6165 4040 6217
rect 3848 6146 4040 6165
rect 3848 6094 3857 6146
rect 3909 6094 3981 6146
rect 4033 6094 4040 6146
rect 3848 6075 4040 6094
rect 3848 6023 3857 6075
rect 3909 6023 3981 6075
rect 4033 6023 4040 6075
rect 3848 6004 4040 6023
rect 3848 5952 3857 6004
rect 3909 5952 3981 6004
rect 4033 5952 4040 6004
rect 683 5812 749 5853
rect 187 5801 749 5812
rect 801 5801 3041 5853
rect 187 5799 3041 5801
rect 187 5747 631 5799
rect 683 5788 3041 5799
rect 683 5747 749 5788
rect 187 5736 749 5747
rect 801 5736 3041 5788
rect 187 5734 3041 5736
rect 187 5682 631 5734
rect 683 5723 3041 5734
rect 683 5682 749 5723
rect 187 5671 749 5682
rect 801 5671 3041 5723
rect 187 5669 3041 5671
rect 187 5617 631 5669
rect 683 5658 3041 5669
rect 683 5617 749 5658
rect 187 5606 749 5617
rect 801 5606 3041 5658
rect 187 5604 3041 5606
rect 187 5552 631 5604
rect 683 5593 3041 5604
rect 683 5552 749 5593
rect 187 5541 749 5552
rect 801 5541 813 5593
rect 865 5541 877 5593
rect 929 5541 941 5593
rect 993 5541 1005 5593
rect 1057 5541 1069 5593
rect 1121 5541 1133 5593
rect 1185 5541 1197 5593
rect 1249 5541 1261 5593
rect 1313 5541 1325 5593
rect 1377 5541 1389 5593
rect 1441 5541 1453 5593
rect 1505 5541 1517 5593
rect 1569 5541 1581 5593
rect 1633 5541 1646 5593
rect 1698 5541 1711 5593
rect 1763 5541 1776 5593
rect 1828 5541 1841 5593
rect 1893 5541 1906 5593
rect 1958 5541 1971 5593
rect 2023 5541 2036 5593
rect 2088 5541 2101 5593
rect 2153 5541 2166 5593
rect 2218 5541 3041 5593
rect 187 5539 3041 5541
rect 187 5487 631 5539
rect 683 5487 3041 5539
rect 187 5475 3041 5487
rect 187 5423 697 5475
rect 749 5423 763 5475
rect 815 5423 829 5475
rect 881 5423 895 5475
rect 947 5423 961 5475
rect 1013 5423 1027 5475
rect 1079 5423 1094 5475
rect 1146 5423 1161 5475
rect 1213 5423 1228 5475
rect 1280 5423 1295 5475
rect 1347 5423 1362 5475
rect 1414 5423 1429 5475
rect 1481 5423 1496 5475
rect 1548 5423 1563 5475
rect 1615 5423 1630 5475
rect 1682 5423 1697 5475
rect 1749 5423 1764 5475
rect 1816 5423 1831 5475
rect 1883 5423 1898 5475
rect 1950 5423 1965 5475
rect 2017 5423 2032 5475
rect 2084 5423 2099 5475
rect 2151 5423 2166 5475
rect 2218 5423 3041 5475
rect 187 5140 3041 5423
tri 3041 5140 3764 5863 sw
rect 3848 5365 4040 5952
rect 8941 6583 10985 6584
rect 11037 6583 11111 6635
rect 11163 6583 11164 6635
rect 8941 6578 11164 6583
rect 8993 6526 9011 6578
rect 9063 6569 11164 6578
rect 9063 6526 10985 6569
rect 8941 6517 10985 6526
rect 11037 6517 11111 6569
rect 11163 6517 11164 6569
rect 8941 6514 11164 6517
rect 8993 6462 9011 6514
rect 9063 6511 11164 6514
rect 9063 6462 9709 6511
rect 8941 6450 9709 6462
rect 8993 6398 9011 6450
rect 9063 6398 9709 6450
rect 8941 6386 9709 6398
rect 8993 6334 9011 6386
rect 9063 6334 9709 6386
rect 8941 6322 9709 6334
rect 8993 6270 9011 6322
rect 9063 6270 9709 6322
rect 8941 6258 9709 6270
rect 8993 6206 9011 6258
rect 9063 6206 9709 6258
rect 8941 6194 9709 6206
rect 8993 6142 9011 6194
rect 9063 6142 9709 6194
rect 8941 6130 9709 6142
rect 8993 6078 9011 6130
rect 9063 6078 9709 6130
rect 8941 6065 9709 6078
rect 8993 6013 9011 6065
rect 9063 6013 9709 6065
rect 8941 6000 9709 6013
rect 8993 5948 9011 6000
rect 9063 5948 9709 6000
rect 8941 5942 9709 5948
tri 9709 5942 10278 6511 nw
rect 3848 5313 3854 5365
rect 3906 5313 3918 5365
rect 3970 5313 3982 5365
rect 4034 5313 4040 5365
rect 3848 5299 4040 5313
rect 187 5101 7379 5140
tri 11163 5132 12222 6191 se
rect 12222 5132 14858 9016
rect 187 5045 5191 5101
rect 5247 5045 5273 5101
rect 5329 5045 5355 5101
rect 5411 5045 5437 5101
rect 5493 5045 5519 5101
rect 5575 5045 5601 5101
rect 5657 5045 5683 5101
rect 5739 5045 5765 5101
rect 5821 5045 5847 5101
rect 5903 5045 5929 5101
rect 5985 5045 6011 5101
rect 6067 5045 6093 5101
rect 6149 5045 6175 5101
rect 6231 5045 6257 5101
rect 6313 5045 6339 5101
rect 6395 5045 6421 5101
rect 6477 5045 6503 5101
rect 6559 5045 6585 5101
rect 6641 5045 6666 5101
rect 6722 5045 6747 5101
rect 6803 5045 6828 5101
rect 6884 5045 6909 5101
rect 6965 5045 6990 5101
rect 7046 5045 7071 5101
rect 7127 5045 7152 5101
rect 7208 5045 7233 5101
rect 7289 5045 7314 5101
rect 7370 5045 7379 5101
rect 187 5021 7379 5045
rect 187 4965 5191 5021
rect 5247 4965 5273 5021
rect 5329 4965 5355 5021
rect 5411 4965 5437 5021
rect 5493 4965 5519 5021
rect 5575 4965 5601 5021
rect 5657 4965 5683 5021
rect 5739 4965 5765 5021
rect 5821 4965 5847 5021
rect 5903 4965 5929 5021
rect 5985 4965 6011 5021
rect 6067 4965 6093 5021
rect 6149 4965 6175 5021
rect 6231 4965 6257 5021
rect 6313 4965 6339 5021
rect 6395 4965 6421 5021
rect 6477 4965 6503 5021
rect 6559 4965 6585 5021
rect 6641 4965 6666 5021
rect 6722 4965 6747 5021
rect 6803 4965 6828 5021
rect 6884 4965 6909 5021
rect 6965 4965 6990 5021
rect 7046 4965 7071 5021
rect 7127 4965 7152 5021
rect 7208 4965 7233 5021
rect 7289 4965 7314 5021
rect 7370 4965 7379 5021
rect 187 4941 7379 4965
rect 187 4885 5191 4941
rect 5247 4885 5273 4941
rect 5329 4885 5355 4941
rect 5411 4885 5437 4941
rect 5493 4885 5519 4941
rect 5575 4885 5601 4941
rect 5657 4885 5683 4941
rect 5739 4885 5765 4941
rect 5821 4885 5847 4941
rect 5903 4885 5929 4941
rect 5985 4885 6011 4941
rect 6067 4885 6093 4941
rect 6149 4885 6175 4941
rect 6231 4885 6257 4941
rect 6313 4885 6339 4941
rect 6395 4885 6421 4941
rect 6477 4885 6503 4941
rect 6559 4885 6585 4941
rect 6641 4885 6666 4941
rect 6722 4885 6747 4941
rect 6803 4885 6828 4941
rect 6884 4885 6909 4941
rect 6965 4885 6990 4941
rect 7046 4885 7071 4941
rect 7127 4885 7152 4941
rect 7208 4885 7233 4941
rect 7289 4885 7314 4941
rect 7370 4885 7379 4941
rect 187 4861 7379 4885
rect 187 4805 5191 4861
rect 5247 4805 5273 4861
rect 5329 4805 5355 4861
rect 5411 4805 5437 4861
rect 5493 4805 5519 4861
rect 5575 4805 5601 4861
rect 5657 4805 5683 4861
rect 5739 4805 5765 4861
rect 5821 4805 5847 4861
rect 5903 4805 5929 4861
rect 5985 4805 6011 4861
rect 6067 4805 6093 4861
rect 6149 4805 6175 4861
rect 6231 4805 6257 4861
rect 6313 4805 6339 4861
rect 6395 4805 6421 4861
rect 6477 4805 6503 4861
rect 6559 4805 6585 4861
rect 6641 4805 6666 4861
rect 6722 4805 6747 4861
rect 6803 4805 6828 4861
rect 6884 4805 6909 4861
rect 6965 4805 6990 4861
rect 7046 4805 7071 4861
rect 7127 4805 7152 4861
rect 7208 4805 7233 4861
rect 7289 4805 7314 4861
rect 7370 4805 7379 4861
rect 187 4781 7379 4805
rect 187 4725 5191 4781
rect 5247 4725 5273 4781
rect 5329 4725 5355 4781
rect 5411 4725 5437 4781
rect 5493 4725 5519 4781
rect 5575 4725 5601 4781
rect 5657 4725 5683 4781
rect 5739 4725 5765 4781
rect 5821 4725 5847 4781
rect 5903 4725 5929 4781
rect 5985 4725 6011 4781
rect 6067 4725 6093 4781
rect 6149 4725 6175 4781
rect 6231 4725 6257 4781
rect 6313 4725 6339 4781
rect 6395 4725 6421 4781
rect 6477 4725 6503 4781
rect 6559 4725 6585 4781
rect 6641 4725 6666 4781
rect 6722 4725 6747 4781
rect 6803 4725 6828 4781
rect 6884 4725 6909 4781
rect 6965 4725 6990 4781
rect 7046 4725 7071 4781
rect 7127 4725 7152 4781
rect 7208 4725 7233 4781
rect 7289 4725 7314 4781
rect 7370 4725 7379 4781
rect 187 4701 7379 4725
rect 187 4645 5191 4701
rect 5247 4645 5273 4701
rect 5329 4645 5355 4701
rect 5411 4645 5437 4701
rect 5493 4645 5519 4701
rect 5575 4645 5601 4701
rect 5657 4645 5683 4701
rect 5739 4645 5765 4701
rect 5821 4645 5847 4701
rect 5903 4645 5929 4701
rect 5985 4645 6011 4701
rect 6067 4645 6093 4701
rect 6149 4645 6175 4701
rect 6231 4645 6257 4701
rect 6313 4645 6339 4701
rect 6395 4645 6421 4701
rect 6477 4645 6503 4701
rect 6559 4645 6585 4701
rect 6641 4645 6666 4701
rect 6722 4645 6747 4701
rect 6803 4645 6828 4701
rect 6884 4645 6909 4701
rect 6965 4645 6990 4701
rect 7046 4645 7071 4701
rect 7127 4645 7152 4701
rect 7208 4645 7233 4701
rect 7289 4645 7314 4701
rect 7370 4645 7379 4701
rect 187 4621 7379 4645
rect 187 4565 5191 4621
rect 5247 4565 5273 4621
rect 5329 4565 5355 4621
rect 5411 4565 5437 4621
rect 5493 4565 5519 4621
rect 5575 4565 5601 4621
rect 5657 4565 5683 4621
rect 5739 4565 5765 4621
rect 5821 4565 5847 4621
rect 5903 4565 5929 4621
rect 5985 4565 6011 4621
rect 6067 4565 6093 4621
rect 6149 4565 6175 4621
rect 6231 4565 6257 4621
rect 6313 4565 6339 4621
rect 6395 4565 6421 4621
rect 6477 4565 6503 4621
rect 6559 4565 6585 4621
rect 6641 4565 6666 4621
rect 6722 4565 6747 4621
rect 6803 4565 6828 4621
rect 6884 4565 6909 4621
rect 6965 4565 6990 4621
rect 7046 4565 7071 4621
rect 7127 4565 7152 4621
rect 7208 4565 7233 4621
rect 7289 4565 7314 4621
rect 7370 4565 7379 4621
rect 187 4541 7379 4565
rect 187 4485 5191 4541
rect 5247 4485 5273 4541
rect 5329 4485 5355 4541
rect 5411 4485 5437 4541
rect 5493 4485 5519 4541
rect 5575 4485 5601 4541
rect 5657 4485 5683 4541
rect 5739 4485 5765 4541
rect 5821 4485 5847 4541
rect 5903 4485 5929 4541
rect 5985 4485 6011 4541
rect 6067 4485 6093 4541
rect 6149 4485 6175 4541
rect 6231 4485 6257 4541
rect 6313 4485 6339 4541
rect 6395 4485 6421 4541
rect 6477 4485 6503 4541
rect 6559 4485 6585 4541
rect 6641 4485 6666 4541
rect 6722 4485 6747 4541
rect 6803 4485 6828 4541
rect 6884 4485 6909 4541
rect 6965 4485 6990 4541
rect 7046 4485 7071 4541
rect 7127 4485 7152 4541
rect 7208 4485 7233 4541
rect 7289 4485 7314 4541
rect 7370 4485 7379 4541
rect 187 4461 7379 4485
rect 187 4405 5191 4461
rect 5247 4405 5273 4461
rect 5329 4405 5355 4461
rect 5411 4405 5437 4461
rect 5493 4405 5519 4461
rect 5575 4405 5601 4461
rect 5657 4405 5683 4461
rect 5739 4405 5765 4461
rect 5821 4405 5847 4461
rect 5903 4405 5929 4461
rect 5985 4405 6011 4461
rect 6067 4405 6093 4461
rect 6149 4405 6175 4461
rect 6231 4405 6257 4461
rect 6313 4405 6339 4461
rect 6395 4405 6421 4461
rect 6477 4405 6503 4461
rect 6559 4405 6585 4461
rect 6641 4405 6666 4461
rect 6722 4405 6747 4461
rect 6803 4405 6828 4461
rect 6884 4405 6909 4461
rect 6965 4405 6990 4461
rect 7046 4405 7071 4461
rect 7127 4405 7152 4461
rect 7208 4405 7233 4461
rect 7289 4405 7314 4461
rect 7370 4405 7379 4461
rect 187 4381 7379 4405
rect 187 4325 5191 4381
rect 5247 4325 5273 4381
rect 5329 4325 5355 4381
rect 5411 4325 5437 4381
rect 5493 4325 5519 4381
rect 5575 4325 5601 4381
rect 5657 4325 5683 4381
rect 5739 4325 5765 4381
rect 5821 4325 5847 4381
rect 5903 4325 5929 4381
rect 5985 4325 6011 4381
rect 6067 4325 6093 4381
rect 6149 4325 6175 4381
rect 6231 4325 6257 4381
rect 6313 4325 6339 4381
rect 6395 4325 6421 4381
rect 6477 4325 6503 4381
rect 6559 4325 6585 4381
rect 6641 4325 6666 4381
rect 6722 4325 6747 4381
rect 6803 4325 6828 4381
rect 6884 4325 6909 4381
rect 6965 4325 6990 4381
rect 7046 4325 7071 4381
rect 7127 4325 7152 4381
rect 7208 4325 7233 4381
rect 7289 4325 7314 4381
rect 7370 4325 7379 4381
rect 187 4301 7379 4325
rect 187 4245 5191 4301
rect 5247 4245 5273 4301
rect 5329 4245 5355 4301
rect 5411 4245 5437 4301
rect 5493 4245 5519 4301
rect 5575 4245 5601 4301
rect 5657 4245 5683 4301
rect 5739 4245 5765 4301
rect 5821 4245 5847 4301
rect 5903 4245 5929 4301
rect 5985 4245 6011 4301
rect 6067 4245 6093 4301
rect 6149 4245 6175 4301
rect 6231 4245 6257 4301
rect 6313 4245 6339 4301
rect 6395 4245 6421 4301
rect 6477 4245 6503 4301
rect 6559 4245 6585 4301
rect 6641 4245 6666 4301
rect 6722 4245 6747 4301
rect 6803 4245 6828 4301
rect 6884 4245 6909 4301
rect 6965 4245 6990 4301
rect 7046 4245 7071 4301
rect 7127 4245 7152 4301
rect 7208 4245 7233 4301
rect 7289 4245 7314 4301
rect 7370 4245 7379 4301
rect 187 4221 7379 4245
rect 187 4165 5191 4221
rect 5247 4165 5273 4221
rect 5329 4165 5355 4221
rect 5411 4165 5437 4221
rect 5493 4165 5519 4221
rect 5575 4165 5601 4221
rect 5657 4165 5683 4221
rect 5739 4165 5765 4221
rect 5821 4165 5847 4221
rect 5903 4165 5929 4221
rect 5985 4165 6011 4221
rect 6067 4165 6093 4221
rect 6149 4165 6175 4221
rect 6231 4165 6257 4221
rect 6313 4165 6339 4221
rect 6395 4165 6421 4221
rect 6477 4165 6503 4221
rect 6559 4165 6585 4221
rect 6641 4165 6666 4221
rect 6722 4165 6747 4221
rect 6803 4165 6828 4221
rect 6884 4165 6909 4221
rect 6965 4165 6990 4221
rect 7046 4165 7071 4221
rect 7127 4165 7152 4221
rect 7208 4165 7233 4221
rect 7289 4165 7314 4221
rect 7370 4165 7379 4221
rect 187 4141 7379 4165
rect 187 4085 5191 4141
rect 5247 4085 5273 4141
rect 5329 4085 5355 4141
rect 5411 4085 5437 4141
rect 5493 4085 5519 4141
rect 5575 4085 5601 4141
rect 5657 4085 5683 4141
rect 5739 4085 5765 4141
rect 5821 4085 5847 4141
rect 5903 4085 5929 4141
rect 5985 4085 6011 4141
rect 6067 4085 6093 4141
rect 6149 4085 6175 4141
rect 6231 4085 6257 4141
rect 6313 4085 6339 4141
rect 6395 4085 6421 4141
rect 6477 4085 6503 4141
rect 6559 4085 6585 4141
rect 6641 4085 6666 4141
rect 6722 4085 6747 4141
rect 6803 4085 6828 4141
rect 6884 4085 6909 4141
rect 6965 4085 6990 4141
rect 7046 4085 7071 4141
rect 7127 4085 7152 4141
rect 7208 4085 7233 4141
rect 7289 4085 7314 4141
rect 7370 4085 7379 4141
rect 187 4061 7379 4085
rect 187 4005 5191 4061
rect 5247 4005 5273 4061
rect 5329 4005 5355 4061
rect 5411 4005 5437 4061
rect 5493 4005 5519 4061
rect 5575 4005 5601 4061
rect 5657 4005 5683 4061
rect 5739 4005 5765 4061
rect 5821 4005 5847 4061
rect 5903 4005 5929 4061
rect 5985 4005 6011 4061
rect 6067 4005 6093 4061
rect 6149 4005 6175 4061
rect 6231 4005 6257 4061
rect 6313 4005 6339 4061
rect 6395 4005 6421 4061
rect 6477 4005 6503 4061
rect 6559 4005 6585 4061
rect 6641 4005 6666 4061
rect 6722 4005 6747 4061
rect 6803 4005 6828 4061
rect 6884 4005 6909 4061
rect 6965 4005 6990 4061
rect 7046 4005 7071 4061
rect 7127 4005 7152 4061
rect 7208 4005 7233 4061
rect 7289 4005 7314 4061
rect 7370 4005 7379 4061
rect 187 4004 7379 4005
rect 187 3952 2771 4004
rect 2823 3952 2838 4004
rect 2890 3952 2905 4004
rect 2957 3952 2972 4004
rect 3024 3952 3039 4004
rect 3091 3952 3106 4004
rect 3158 3952 3173 4004
rect 3225 3952 3240 4004
rect 3292 3952 3307 4004
rect 3359 3952 3374 4004
rect 3426 3952 3441 4004
rect 3493 3952 3508 4004
rect 3560 3952 3575 4004
rect 3627 3952 3642 4004
rect 3694 3952 3708 4004
rect 3760 3952 3774 4004
rect 3826 3981 7379 4004
rect 3826 3952 5191 3981
rect 187 3936 5191 3952
rect 187 3884 2771 3936
rect 2823 3884 2838 3936
rect 2890 3884 2905 3936
rect 2957 3884 2972 3936
rect 3024 3884 3039 3936
rect 3091 3884 3106 3936
rect 3158 3884 3173 3936
rect 3225 3884 3240 3936
rect 3292 3884 3307 3936
rect 3359 3884 3374 3936
rect 3426 3884 3441 3936
rect 3493 3884 3508 3936
rect 3560 3884 3575 3936
rect 3627 3884 3642 3936
rect 3694 3884 3708 3936
rect 3760 3884 3774 3936
rect 3826 3925 5191 3936
rect 5247 3925 5273 3981
rect 5329 3925 5355 3981
rect 5411 3925 5437 3981
rect 5493 3925 5519 3981
rect 5575 3925 5601 3981
rect 5657 3925 5683 3981
rect 5739 3925 5765 3981
rect 5821 3925 5847 3981
rect 5903 3925 5929 3981
rect 5985 3925 6011 3981
rect 6067 3925 6093 3981
rect 6149 3925 6175 3981
rect 6231 3925 6257 3981
rect 6313 3925 6339 3981
rect 6395 3925 6421 3981
rect 6477 3925 6503 3981
rect 6559 3925 6585 3981
rect 6641 3925 6666 3981
rect 6722 3925 6747 3981
rect 6803 3925 6828 3981
rect 6884 3925 6909 3981
rect 6965 3925 6990 3981
rect 7046 3925 7071 3981
rect 7127 3925 7152 3981
rect 7208 3925 7233 3981
rect 7289 3925 7314 3981
rect 7370 3925 7379 3981
rect 3826 3901 7379 3925
rect 3826 3884 5191 3901
rect 187 3868 5191 3884
rect 187 3816 2771 3868
rect 2823 3816 2838 3868
rect 2890 3816 2905 3868
rect 2957 3816 2972 3868
rect 3024 3816 3039 3868
rect 3091 3816 3106 3868
rect 3158 3816 3173 3868
rect 3225 3816 3240 3868
rect 3292 3816 3307 3868
rect 3359 3816 3374 3868
rect 3426 3816 3441 3868
rect 3493 3816 3508 3868
rect 3560 3816 3575 3868
rect 3627 3816 3642 3868
rect 3694 3816 3708 3868
rect 3760 3816 3774 3868
rect 3826 3845 5191 3868
rect 5247 3845 5273 3901
rect 5329 3845 5355 3901
rect 5411 3845 5437 3901
rect 5493 3845 5519 3901
rect 5575 3845 5601 3901
rect 5657 3845 5683 3901
rect 5739 3845 5765 3901
rect 5821 3845 5847 3901
rect 5903 3845 5929 3901
rect 5985 3845 6011 3901
rect 6067 3845 6093 3901
rect 6149 3845 6175 3901
rect 6231 3845 6257 3901
rect 6313 3845 6339 3901
rect 6395 3845 6421 3901
rect 6477 3845 6503 3901
rect 6559 3845 6585 3901
rect 6641 3845 6666 3901
rect 6722 3845 6747 3901
rect 6803 3845 6828 3901
rect 6884 3845 6909 3901
rect 6965 3845 6990 3901
rect 7046 3845 7071 3901
rect 7127 3845 7152 3901
rect 7208 3845 7233 3901
rect 7289 3845 7314 3901
rect 7370 3845 7379 3901
rect 3826 3821 7379 3845
rect 3826 3816 5191 3821
rect 187 3800 5191 3816
rect 187 3748 2771 3800
rect 2823 3748 2838 3800
rect 2890 3748 2905 3800
rect 2957 3748 2972 3800
rect 3024 3748 3039 3800
rect 3091 3748 3106 3800
rect 3158 3748 3173 3800
rect 3225 3748 3240 3800
rect 3292 3748 3307 3800
rect 3359 3748 3374 3800
rect 3426 3748 3441 3800
rect 3493 3748 3508 3800
rect 3560 3748 3575 3800
rect 3627 3748 3642 3800
rect 3694 3748 3708 3800
rect 3760 3748 3774 3800
rect 3826 3765 5191 3800
rect 5247 3765 5273 3821
rect 5329 3765 5355 3821
rect 5411 3765 5437 3821
rect 5493 3765 5519 3821
rect 5575 3765 5601 3821
rect 5657 3765 5683 3821
rect 5739 3765 5765 3821
rect 5821 3765 5847 3821
rect 5903 3765 5929 3821
rect 5985 3765 6011 3821
rect 6067 3765 6093 3821
rect 6149 3765 6175 3821
rect 6231 3765 6257 3821
rect 6313 3765 6339 3821
rect 6395 3765 6421 3821
rect 6477 3765 6503 3821
rect 6559 3765 6585 3821
rect 6641 3765 6666 3821
rect 6722 3765 6747 3821
rect 6803 3765 6828 3821
rect 6884 3765 6909 3821
rect 6965 3765 6990 3821
rect 7046 3765 7071 3821
rect 7127 3765 7152 3821
rect 7208 3765 7233 3821
rect 7289 3765 7314 3821
rect 7370 3765 7379 3821
rect 3826 3748 7379 3765
rect 187 3741 7379 3748
rect 187 3732 5191 3741
rect 187 3680 2771 3732
rect 2823 3680 2838 3732
rect 2890 3680 2905 3732
rect 2957 3680 2972 3732
rect 3024 3680 3039 3732
rect 3091 3680 3106 3732
rect 3158 3680 3173 3732
rect 3225 3680 3240 3732
rect 3292 3680 3307 3732
rect 3359 3680 3374 3732
rect 3426 3680 3441 3732
rect 3493 3680 3508 3732
rect 3560 3680 3575 3732
rect 3627 3680 3642 3732
rect 3694 3680 3708 3732
rect 3760 3680 3774 3732
rect 3826 3685 5191 3732
rect 5247 3685 5273 3741
rect 5329 3685 5355 3741
rect 5411 3685 5437 3741
rect 5493 3685 5519 3741
rect 5575 3685 5601 3741
rect 5657 3685 5683 3741
rect 5739 3685 5765 3741
rect 5821 3685 5847 3741
rect 5903 3685 5929 3741
rect 5985 3685 6011 3741
rect 6067 3685 6093 3741
rect 6149 3685 6175 3741
rect 6231 3685 6257 3741
rect 6313 3685 6339 3741
rect 6395 3685 6421 3741
rect 6477 3685 6503 3741
rect 6559 3685 6585 3741
rect 6641 3685 6666 3741
rect 6722 3685 6747 3741
rect 6803 3685 6828 3741
rect 6884 3685 6909 3741
rect 6965 3685 6990 3741
rect 7046 3685 7071 3741
rect 7127 3685 7152 3741
rect 7208 3685 7233 3741
rect 7289 3685 7314 3741
rect 7370 3685 7379 3741
rect 3826 3680 7379 3685
rect 187 3664 7379 3680
rect 187 3612 2771 3664
rect 2823 3612 2838 3664
rect 2890 3612 2905 3664
rect 2957 3612 2972 3664
rect 3024 3612 3039 3664
rect 3091 3612 3106 3664
rect 3158 3612 3173 3664
rect 3225 3612 3240 3664
rect 3292 3612 3307 3664
rect 3359 3612 3374 3664
rect 3426 3612 3441 3664
rect 3493 3612 3508 3664
rect 3560 3612 3575 3664
rect 3627 3612 3642 3664
rect 3694 3612 3708 3664
rect 3760 3612 3774 3664
rect 3826 3661 7379 3664
rect 3826 3612 5191 3661
rect 187 3605 5191 3612
rect 5247 3605 5273 3661
rect 5329 3605 5355 3661
rect 5411 3605 5437 3661
rect 5493 3605 5519 3661
rect 5575 3605 5601 3661
rect 5657 3605 5683 3661
rect 5739 3605 5765 3661
rect 5821 3605 5847 3661
rect 5903 3605 5929 3661
rect 5985 3605 6011 3661
rect 6067 3605 6093 3661
rect 6149 3605 6175 3661
rect 6231 3605 6257 3661
rect 6313 3605 6339 3661
rect 6395 3605 6421 3661
rect 6477 3605 6503 3661
rect 6559 3605 6585 3661
rect 6641 3605 6666 3661
rect 6722 3605 6747 3661
rect 6803 3605 6828 3661
rect 6884 3605 6909 3661
rect 6965 3605 6990 3661
rect 7046 3605 7071 3661
rect 7127 3605 7152 3661
rect 7208 3605 7233 3661
rect 7289 3605 7314 3661
rect 7370 3605 7379 3661
rect 187 3596 7379 3605
rect 187 3544 2771 3596
rect 2823 3544 2838 3596
rect 2890 3544 2905 3596
rect 2957 3544 2972 3596
rect 3024 3544 3039 3596
rect 3091 3544 3106 3596
rect 3158 3544 3173 3596
rect 3225 3544 3240 3596
rect 3292 3544 3307 3596
rect 3359 3544 3374 3596
rect 3426 3544 3441 3596
rect 3493 3544 3508 3596
rect 3560 3544 3575 3596
rect 3627 3544 3642 3596
rect 3694 3544 3708 3596
rect 3760 3544 3774 3596
rect 3826 3581 7379 3596
rect 3826 3544 5191 3581
rect 187 3528 5191 3544
rect 187 3476 2771 3528
rect 2823 3476 2838 3528
rect 2890 3476 2905 3528
rect 2957 3476 2972 3528
rect 3024 3476 3039 3528
rect 3091 3476 3106 3528
rect 3158 3476 3173 3528
rect 3225 3476 3240 3528
rect 3292 3476 3307 3528
rect 3359 3476 3374 3528
rect 3426 3476 3441 3528
rect 3493 3476 3508 3528
rect 3560 3476 3575 3528
rect 3627 3476 3642 3528
rect 3694 3476 3708 3528
rect 3760 3476 3774 3528
rect 3826 3525 5191 3528
rect 5247 3525 5273 3581
rect 5329 3525 5355 3581
rect 5411 3525 5437 3581
rect 5493 3525 5519 3581
rect 5575 3525 5601 3581
rect 5657 3525 5683 3581
rect 5739 3525 5765 3581
rect 5821 3525 5847 3581
rect 5903 3525 5929 3581
rect 5985 3525 6011 3581
rect 6067 3525 6093 3581
rect 6149 3525 6175 3581
rect 6231 3525 6257 3581
rect 6313 3525 6339 3581
rect 6395 3525 6421 3581
rect 6477 3525 6503 3581
rect 6559 3525 6585 3581
rect 6641 3525 6666 3581
rect 6722 3525 6747 3581
rect 6803 3525 6828 3581
rect 6884 3525 6909 3581
rect 6965 3525 6990 3581
rect 7046 3525 7071 3581
rect 7127 3525 7152 3581
rect 7208 3525 7233 3581
rect 7289 3525 7314 3581
rect 7370 3525 7379 3581
rect 3826 3501 7379 3525
rect 3826 3476 5191 3501
rect 187 3445 5191 3476
rect 5247 3445 5273 3501
rect 5329 3445 5355 3501
rect 5411 3445 5437 3501
rect 5493 3445 5519 3501
rect 5575 3445 5601 3501
rect 5657 3445 5683 3501
rect 5739 3445 5765 3501
rect 5821 3445 5847 3501
rect 5903 3445 5929 3501
rect 5985 3445 6011 3501
rect 6067 3445 6093 3501
rect 6149 3445 6175 3501
rect 6231 3445 6257 3501
rect 6313 3445 6339 3501
rect 6395 3445 6421 3501
rect 6477 3445 6503 3501
rect 6559 3445 6585 3501
rect 6641 3445 6666 3501
rect 6722 3445 6747 3501
rect 6803 3445 6828 3501
rect 6884 3445 6909 3501
rect 6965 3445 6990 3501
rect 7046 3445 7071 3501
rect 7127 3445 7152 3501
rect 7208 3445 7233 3501
rect 7289 3445 7314 3501
rect 7370 3445 7379 3501
rect 187 3421 7379 3445
rect 187 3365 5191 3421
rect 5247 3365 5273 3421
rect 5329 3365 5355 3421
rect 5411 3365 5437 3421
rect 5493 3365 5519 3421
rect 5575 3365 5601 3421
rect 5657 3365 5683 3421
rect 5739 3365 5765 3421
rect 5821 3365 5847 3421
rect 5903 3365 5929 3421
rect 5985 3365 6011 3421
rect 6067 3365 6093 3421
rect 6149 3365 6175 3421
rect 6231 3365 6257 3421
rect 6313 3365 6339 3421
rect 6395 3365 6421 3421
rect 6477 3365 6503 3421
rect 6559 3365 6585 3421
rect 6641 3365 6666 3421
rect 6722 3365 6747 3421
rect 6803 3365 6828 3421
rect 6884 3365 6909 3421
rect 6965 3365 6990 3421
rect 7046 3365 7071 3421
rect 7127 3365 7152 3421
rect 7208 3365 7233 3421
rect 7289 3365 7314 3421
rect 7370 3365 7379 3421
rect 187 3341 7379 3365
rect 187 3285 5191 3341
rect 5247 3285 5273 3341
rect 5329 3285 5355 3341
rect 5411 3285 5437 3341
rect 5493 3285 5519 3341
rect 5575 3285 5601 3341
rect 5657 3285 5683 3341
rect 5739 3285 5765 3341
rect 5821 3285 5847 3341
rect 5903 3285 5929 3341
rect 5985 3285 6011 3341
rect 6067 3285 6093 3341
rect 6149 3285 6175 3341
rect 6231 3285 6257 3341
rect 6313 3285 6339 3341
rect 6395 3285 6421 3341
rect 6477 3285 6503 3341
rect 6559 3285 6585 3341
rect 6641 3285 6666 3341
rect 6722 3285 6747 3341
rect 6803 3285 6828 3341
rect 6884 3285 6909 3341
rect 6965 3285 6990 3341
rect 7046 3285 7071 3341
rect 7127 3285 7152 3341
rect 7208 3285 7233 3341
rect 7289 3285 7314 3341
rect 7370 3285 7379 3341
rect 187 3261 7379 3285
rect 187 3205 5191 3261
rect 5247 3205 5273 3261
rect 5329 3205 5355 3261
rect 5411 3205 5437 3261
rect 5493 3205 5519 3261
rect 5575 3205 5601 3261
rect 5657 3205 5683 3261
rect 5739 3205 5765 3261
rect 5821 3205 5847 3261
rect 5903 3205 5929 3261
rect 5985 3205 6011 3261
rect 6067 3205 6093 3261
rect 6149 3205 6175 3261
rect 6231 3205 6257 3261
rect 6313 3205 6339 3261
rect 6395 3205 6421 3261
rect 6477 3205 6503 3261
rect 6559 3205 6585 3261
rect 6641 3205 6666 3261
rect 6722 3205 6747 3261
rect 6803 3205 6828 3261
rect 6884 3205 6909 3261
rect 6965 3205 6990 3261
rect 7046 3205 7071 3261
rect 7127 3205 7152 3261
rect 7208 3205 7233 3261
rect 7289 3205 7314 3261
rect 7370 3205 7379 3261
rect 187 3181 7379 3205
rect 187 3125 5191 3181
rect 5247 3125 5273 3181
rect 5329 3125 5355 3181
rect 5411 3125 5437 3181
rect 5493 3125 5519 3181
rect 5575 3125 5601 3181
rect 5657 3125 5683 3181
rect 5739 3125 5765 3181
rect 5821 3125 5847 3181
rect 5903 3125 5929 3181
rect 5985 3125 6011 3181
rect 6067 3125 6093 3181
rect 6149 3125 6175 3181
rect 6231 3125 6257 3181
rect 6313 3125 6339 3181
rect 6395 3125 6421 3181
rect 6477 3125 6503 3181
rect 6559 3125 6585 3181
rect 6641 3125 6666 3181
rect 6722 3125 6747 3181
rect 6803 3125 6828 3181
rect 6884 3125 6909 3181
rect 6965 3125 6990 3181
rect 7046 3125 7071 3181
rect 7127 3125 7152 3181
rect 7208 3125 7233 3181
rect 7289 3125 7314 3181
rect 7370 3125 7379 3181
rect 187 3101 7379 3125
rect 187 3045 5191 3101
rect 5247 3045 5273 3101
rect 5329 3045 5355 3101
rect 5411 3045 5437 3101
rect 5493 3045 5519 3101
rect 5575 3045 5601 3101
rect 5657 3045 5683 3101
rect 5739 3045 5765 3101
rect 5821 3045 5847 3101
rect 5903 3045 5929 3101
rect 5985 3045 6011 3101
rect 6067 3045 6093 3101
rect 6149 3045 6175 3101
rect 6231 3045 6257 3101
rect 6313 3045 6339 3101
rect 6395 3045 6421 3101
rect 6477 3045 6503 3101
rect 6559 3045 6585 3101
rect 6641 3045 6666 3101
rect 6722 3045 6747 3101
rect 6803 3045 6828 3101
rect 6884 3045 6909 3101
rect 6965 3045 6990 3101
rect 7046 3045 7071 3101
rect 7127 3045 7152 3101
rect 7208 3045 7233 3101
rect 7289 3045 7314 3101
rect 7370 3045 7379 3101
rect 187 3021 7379 3045
rect 187 2965 5191 3021
rect 5247 2965 5273 3021
rect 5329 2965 5355 3021
rect 5411 2965 5437 3021
rect 5493 2965 5519 3021
rect 5575 2965 5601 3021
rect 5657 2965 5683 3021
rect 5739 2965 5765 3021
rect 5821 2965 5847 3021
rect 5903 2965 5929 3021
rect 5985 2965 6011 3021
rect 6067 2965 6093 3021
rect 6149 2965 6175 3021
rect 6231 2965 6257 3021
rect 6313 2965 6339 3021
rect 6395 2965 6421 3021
rect 6477 2965 6503 3021
rect 6559 2965 6585 3021
rect 6641 2965 6666 3021
rect 6722 2965 6747 3021
rect 6803 2965 6828 3021
rect 6884 2965 6909 3021
rect 6965 2965 6990 3021
rect 7046 2965 7071 3021
rect 7127 2965 7152 3021
rect 7208 2965 7233 3021
rect 7289 2965 7314 3021
rect 7370 2965 7379 3021
rect 187 2941 7379 2965
rect 187 2885 5191 2941
rect 5247 2885 5273 2941
rect 5329 2885 5355 2941
rect 5411 2885 5437 2941
rect 5493 2885 5519 2941
rect 5575 2885 5601 2941
rect 5657 2885 5683 2941
rect 5739 2885 5765 2941
rect 5821 2885 5847 2941
rect 5903 2885 5929 2941
rect 5985 2885 6011 2941
rect 6067 2885 6093 2941
rect 6149 2885 6175 2941
rect 6231 2885 6257 2941
rect 6313 2885 6339 2941
rect 6395 2885 6421 2941
rect 6477 2885 6503 2941
rect 6559 2885 6585 2941
rect 6641 2885 6666 2941
rect 6722 2885 6747 2941
rect 6803 2885 6828 2941
rect 6884 2885 6909 2941
rect 6965 2885 6990 2941
rect 7046 2885 7071 2941
rect 7127 2885 7152 2941
rect 7208 2885 7233 2941
rect 7289 2885 7314 2941
rect 7370 2885 7379 2941
rect 187 2861 7379 2885
rect 187 2805 5191 2861
rect 5247 2805 5273 2861
rect 5329 2805 5355 2861
rect 5411 2805 5437 2861
rect 5493 2805 5519 2861
rect 5575 2805 5601 2861
rect 5657 2805 5683 2861
rect 5739 2805 5765 2861
rect 5821 2805 5847 2861
rect 5903 2805 5929 2861
rect 5985 2805 6011 2861
rect 6067 2805 6093 2861
rect 6149 2805 6175 2861
rect 6231 2805 6257 2861
rect 6313 2805 6339 2861
rect 6395 2805 6421 2861
rect 6477 2805 6503 2861
rect 6559 2805 6585 2861
rect 6641 2805 6666 2861
rect 6722 2805 6747 2861
rect 6803 2805 6828 2861
rect 6884 2805 6909 2861
rect 6965 2805 6990 2861
rect 7046 2805 7071 2861
rect 7127 2805 7152 2861
rect 7208 2805 7233 2861
rect 7289 2805 7314 2861
rect 7370 2805 7379 2861
rect 187 2792 7379 2805
rect 187 2740 2766 2792
rect 2818 2740 2831 2792
rect 2883 2740 2896 2792
rect 2948 2740 2961 2792
rect 3013 2740 3026 2792
rect 3078 2740 3091 2792
rect 3143 2740 3156 2792
rect 3208 2740 3221 2792
rect 3273 2740 3285 2792
rect 3337 2740 3349 2792
rect 3401 2740 3413 2792
rect 3465 2740 3477 2792
rect 3529 2740 3541 2792
rect 3593 2740 3605 2792
rect 3657 2740 3669 2792
rect 3721 2740 3733 2792
rect 3785 2740 3797 2792
rect 3849 2740 3861 2792
rect 3913 2740 3925 2792
rect 3977 2740 3989 2792
rect 4041 2740 4053 2792
rect 4105 2740 4117 2792
rect 4169 2740 4181 2792
rect 4233 2740 4245 2792
rect 4297 2740 4309 2792
rect 4361 2740 4373 2792
rect 4425 2740 4437 2792
rect 4489 2740 4501 2792
rect 4553 2740 4565 2792
rect 4617 2740 4629 2792
rect 4681 2740 4693 2792
rect 4745 2740 4757 2792
rect 4809 2740 4821 2792
rect 4873 2781 7379 2792
rect 4873 2740 5191 2781
rect 187 2726 5191 2740
rect 187 2674 2766 2726
rect 2818 2674 2831 2726
rect 2883 2674 2896 2726
rect 2948 2674 2961 2726
rect 3013 2674 3026 2726
rect 3078 2674 3091 2726
rect 3143 2674 3156 2726
rect 3208 2674 3221 2726
rect 3273 2674 3285 2726
rect 3337 2674 3349 2726
rect 3401 2674 3413 2726
rect 3465 2674 3477 2726
rect 3529 2674 3541 2726
rect 3593 2674 3605 2726
rect 3657 2674 3669 2726
rect 3721 2674 3733 2726
rect 3785 2674 3797 2726
rect 3849 2674 3861 2726
rect 3913 2674 3925 2726
rect 3977 2674 3989 2726
rect 4041 2674 4053 2726
rect 4105 2674 4117 2726
rect 4169 2674 4181 2726
rect 4233 2674 4245 2726
rect 4297 2674 4309 2726
rect 4361 2674 4373 2726
rect 4425 2674 4437 2726
rect 4489 2674 4501 2726
rect 4553 2674 4565 2726
rect 4617 2674 4629 2726
rect 4681 2674 4693 2726
rect 4745 2674 4757 2726
rect 4809 2674 4821 2726
rect 4873 2725 5191 2726
rect 5247 2725 5273 2781
rect 5329 2725 5355 2781
rect 5411 2725 5437 2781
rect 5493 2725 5519 2781
rect 5575 2725 5601 2781
rect 5657 2725 5683 2781
rect 5739 2725 5765 2781
rect 5821 2725 5847 2781
rect 5903 2725 5929 2781
rect 5985 2725 6011 2781
rect 6067 2725 6093 2781
rect 6149 2725 6175 2781
rect 6231 2725 6257 2781
rect 6313 2725 6339 2781
rect 6395 2725 6421 2781
rect 6477 2725 6503 2781
rect 6559 2725 6585 2781
rect 6641 2725 6666 2781
rect 6722 2725 6747 2781
rect 6803 2725 6828 2781
rect 6884 2725 6909 2781
rect 6965 2725 6990 2781
rect 7046 2725 7071 2781
rect 7127 2725 7152 2781
rect 7208 2725 7233 2781
rect 7289 2725 7314 2781
rect 7370 2725 7379 2781
rect 4873 2701 7379 2725
rect 4873 2674 5191 2701
rect 187 2660 5191 2674
rect 187 2608 2766 2660
rect 2818 2608 2831 2660
rect 2883 2608 2896 2660
rect 2948 2608 2961 2660
rect 3013 2608 3026 2660
rect 3078 2608 3091 2660
rect 3143 2608 3156 2660
rect 3208 2608 3221 2660
rect 3273 2608 3285 2660
rect 3337 2608 3349 2660
rect 3401 2608 3413 2660
rect 3465 2608 3477 2660
rect 3529 2608 3541 2660
rect 3593 2608 3605 2660
rect 3657 2608 3669 2660
rect 3721 2608 3733 2660
rect 3785 2608 3797 2660
rect 3849 2608 3861 2660
rect 3913 2608 3925 2660
rect 3977 2608 3989 2660
rect 4041 2608 4053 2660
rect 4105 2608 4117 2660
rect 4169 2608 4181 2660
rect 4233 2608 4245 2660
rect 4297 2608 4309 2660
rect 4361 2608 4373 2660
rect 4425 2608 4437 2660
rect 4489 2608 4501 2660
rect 4553 2608 4565 2660
rect 4617 2608 4629 2660
rect 4681 2608 4693 2660
rect 4745 2608 4757 2660
rect 4809 2608 4821 2660
rect 4873 2645 5191 2660
rect 5247 2645 5273 2701
rect 5329 2645 5355 2701
rect 5411 2645 5437 2701
rect 5493 2645 5519 2701
rect 5575 2645 5601 2701
rect 5657 2645 5683 2701
rect 5739 2645 5765 2701
rect 5821 2645 5847 2701
rect 5903 2645 5929 2701
rect 5985 2645 6011 2701
rect 6067 2645 6093 2701
rect 6149 2645 6175 2701
rect 6231 2645 6257 2701
rect 6313 2645 6339 2701
rect 6395 2645 6421 2701
rect 6477 2645 6503 2701
rect 6559 2645 6585 2701
rect 6641 2645 6666 2701
rect 6722 2645 6747 2701
rect 6803 2645 6828 2701
rect 6884 2645 6909 2701
rect 6965 2645 6990 2701
rect 7046 2645 7071 2701
rect 7127 2645 7152 2701
rect 7208 2645 7233 2701
rect 7289 2645 7314 2701
rect 7370 2645 7379 2701
rect 4873 2621 7379 2645
rect 4873 2608 5191 2621
rect 187 2594 5191 2608
rect 187 2542 2766 2594
rect 2818 2542 2831 2594
rect 2883 2542 2896 2594
rect 2948 2542 2961 2594
rect 3013 2542 3026 2594
rect 3078 2542 3091 2594
rect 3143 2542 3156 2594
rect 3208 2542 3221 2594
rect 3273 2542 3285 2594
rect 3337 2542 3349 2594
rect 3401 2542 3413 2594
rect 3465 2542 3477 2594
rect 3529 2542 3541 2594
rect 3593 2542 3605 2594
rect 3657 2542 3669 2594
rect 3721 2542 3733 2594
rect 3785 2542 3797 2594
rect 3849 2542 3861 2594
rect 3913 2542 3925 2594
rect 3977 2542 3989 2594
rect 4041 2542 4053 2594
rect 4105 2542 4117 2594
rect 4169 2542 4181 2594
rect 4233 2542 4245 2594
rect 4297 2542 4309 2594
rect 4361 2542 4373 2594
rect 4425 2542 4437 2594
rect 4489 2542 4501 2594
rect 4553 2542 4565 2594
rect 4617 2542 4629 2594
rect 4681 2542 4693 2594
rect 4745 2542 4757 2594
rect 4809 2542 4821 2594
rect 4873 2565 5191 2594
rect 5247 2565 5273 2621
rect 5329 2565 5355 2621
rect 5411 2565 5437 2621
rect 5493 2565 5519 2621
rect 5575 2565 5601 2621
rect 5657 2565 5683 2621
rect 5739 2565 5765 2621
rect 5821 2565 5847 2621
rect 5903 2565 5929 2621
rect 5985 2565 6011 2621
rect 6067 2565 6093 2621
rect 6149 2565 6175 2621
rect 6231 2565 6257 2621
rect 6313 2565 6339 2621
rect 6395 2565 6421 2621
rect 6477 2565 6503 2621
rect 6559 2565 6585 2621
rect 6641 2565 6666 2621
rect 6722 2565 6747 2621
rect 6803 2565 6828 2621
rect 6884 2565 6909 2621
rect 6965 2565 6990 2621
rect 7046 2565 7071 2621
rect 7127 2565 7152 2621
rect 7208 2565 7233 2621
rect 7289 2565 7314 2621
rect 7370 2565 7379 2621
rect 4873 2542 7379 2565
rect 187 2541 7379 2542
rect 187 2528 5191 2541
rect 187 2476 2766 2528
rect 2818 2476 2831 2528
rect 2883 2476 2896 2528
rect 2948 2476 2961 2528
rect 3013 2476 3026 2528
rect 3078 2476 3091 2528
rect 3143 2476 3156 2528
rect 3208 2476 3221 2528
rect 3273 2476 3285 2528
rect 3337 2476 3349 2528
rect 3401 2476 3413 2528
rect 3465 2476 3477 2528
rect 3529 2476 3541 2528
rect 3593 2476 3605 2528
rect 3657 2476 3669 2528
rect 3721 2476 3733 2528
rect 3785 2476 3797 2528
rect 3849 2476 3861 2528
rect 3913 2476 3925 2528
rect 3977 2476 3989 2528
rect 4041 2476 4053 2528
rect 4105 2476 4117 2528
rect 4169 2476 4181 2528
rect 4233 2476 4245 2528
rect 4297 2476 4309 2528
rect 4361 2476 4373 2528
rect 4425 2476 4437 2528
rect 4489 2476 4501 2528
rect 4553 2476 4565 2528
rect 4617 2476 4629 2528
rect 4681 2476 4693 2528
rect 4745 2476 4757 2528
rect 4809 2476 4821 2528
rect 4873 2485 5191 2528
rect 5247 2485 5273 2541
rect 5329 2485 5355 2541
rect 5411 2485 5437 2541
rect 5493 2485 5519 2541
rect 5575 2485 5601 2541
rect 5657 2485 5683 2541
rect 5739 2485 5765 2541
rect 5821 2485 5847 2541
rect 5903 2485 5929 2541
rect 5985 2485 6011 2541
rect 6067 2485 6093 2541
rect 6149 2485 6175 2541
rect 6231 2485 6257 2541
rect 6313 2485 6339 2541
rect 6395 2485 6421 2541
rect 6477 2485 6503 2541
rect 6559 2485 6585 2541
rect 6641 2485 6666 2541
rect 6722 2485 6747 2541
rect 6803 2485 6828 2541
rect 6884 2485 6909 2541
rect 6965 2485 6990 2541
rect 7046 2485 7071 2541
rect 7127 2485 7152 2541
rect 7208 2485 7233 2541
rect 7289 2485 7314 2541
rect 7370 2485 7379 2541
rect 4873 2480 7379 2485
rect 7578 5092 14858 5132
rect 7578 5036 7587 5092
rect 7643 5036 7669 5092
rect 7725 5036 7751 5092
rect 7807 5036 7833 5092
rect 7889 5036 7915 5092
rect 7971 5036 7997 5092
rect 8053 5036 8079 5092
rect 8135 5036 8161 5092
rect 8217 5036 8243 5092
rect 8299 5036 8325 5092
rect 8381 5036 8407 5092
rect 8463 5036 8489 5092
rect 8545 5036 8571 5092
rect 8627 5036 8653 5092
rect 8709 5036 8735 5092
rect 8791 5036 8817 5092
rect 8873 5036 8899 5092
rect 8955 5036 8981 5092
rect 9037 5036 9063 5092
rect 9119 5036 9145 5092
rect 9201 5036 9227 5092
rect 9283 5036 9308 5092
rect 9364 5036 9389 5092
rect 9445 5036 9470 5092
rect 9526 5036 9551 5092
rect 9607 5036 9632 5092
rect 9688 5036 9713 5092
rect 9769 5036 14858 5092
rect 7578 5012 14858 5036
rect 7578 4956 7587 5012
rect 7643 4956 7669 5012
rect 7725 4956 7751 5012
rect 7807 4956 7833 5012
rect 7889 4956 7915 5012
rect 7971 4956 7997 5012
rect 8053 4956 8079 5012
rect 8135 4956 8161 5012
rect 8217 4956 8243 5012
rect 8299 4956 8325 5012
rect 8381 4956 8407 5012
rect 8463 4956 8489 5012
rect 8545 4956 8571 5012
rect 8627 4956 8653 5012
rect 8709 4956 8735 5012
rect 8791 4956 8817 5012
rect 8873 4956 8899 5012
rect 8955 4956 8981 5012
rect 9037 4956 9063 5012
rect 9119 4956 9145 5012
rect 9201 4956 9227 5012
rect 9283 4956 9308 5012
rect 9364 4956 9389 5012
rect 9445 4956 9470 5012
rect 9526 4956 9551 5012
rect 9607 4956 9632 5012
rect 9688 4956 9713 5012
rect 9769 4956 14858 5012
rect 7578 4932 14858 4956
rect 7578 4876 7587 4932
rect 7643 4876 7669 4932
rect 7725 4876 7751 4932
rect 7807 4876 7833 4932
rect 7889 4876 7915 4932
rect 7971 4876 7997 4932
rect 8053 4876 8079 4932
rect 8135 4876 8161 4932
rect 8217 4876 8243 4932
rect 8299 4876 8325 4932
rect 8381 4876 8407 4932
rect 8463 4876 8489 4932
rect 8545 4876 8571 4932
rect 8627 4876 8653 4932
rect 8709 4876 8735 4932
rect 8791 4876 8817 4932
rect 8873 4876 8899 4932
rect 8955 4876 8981 4932
rect 9037 4876 9063 4932
rect 9119 4876 9145 4932
rect 9201 4876 9227 4932
rect 9283 4876 9308 4932
rect 9364 4876 9389 4932
rect 9445 4876 9470 4932
rect 9526 4876 9551 4932
rect 9607 4876 9632 4932
rect 9688 4876 9713 4932
rect 9769 4876 14858 4932
rect 7578 4852 14858 4876
rect 7578 4796 7587 4852
rect 7643 4796 7669 4852
rect 7725 4796 7751 4852
rect 7807 4796 7833 4852
rect 7889 4796 7915 4852
rect 7971 4796 7997 4852
rect 8053 4796 8079 4852
rect 8135 4796 8161 4852
rect 8217 4796 8243 4852
rect 8299 4796 8325 4852
rect 8381 4796 8407 4852
rect 8463 4796 8489 4852
rect 8545 4796 8571 4852
rect 8627 4796 8653 4852
rect 8709 4796 8735 4852
rect 8791 4796 8817 4852
rect 8873 4796 8899 4852
rect 8955 4796 8981 4852
rect 9037 4796 9063 4852
rect 9119 4796 9145 4852
rect 9201 4796 9227 4852
rect 9283 4796 9308 4852
rect 9364 4796 9389 4852
rect 9445 4796 9470 4852
rect 9526 4796 9551 4852
rect 9607 4796 9632 4852
rect 9688 4796 9713 4852
rect 9769 4796 14858 4852
rect 7578 4772 14858 4796
rect 7578 4716 7587 4772
rect 7643 4716 7669 4772
rect 7725 4716 7751 4772
rect 7807 4716 7833 4772
rect 7889 4716 7915 4772
rect 7971 4716 7997 4772
rect 8053 4716 8079 4772
rect 8135 4716 8161 4772
rect 8217 4716 8243 4772
rect 8299 4716 8325 4772
rect 8381 4716 8407 4772
rect 8463 4716 8489 4772
rect 8545 4716 8571 4772
rect 8627 4716 8653 4772
rect 8709 4716 8735 4772
rect 8791 4716 8817 4772
rect 8873 4716 8899 4772
rect 8955 4716 8981 4772
rect 9037 4716 9063 4772
rect 9119 4716 9145 4772
rect 9201 4716 9227 4772
rect 9283 4716 9308 4772
rect 9364 4716 9389 4772
rect 9445 4716 9470 4772
rect 9526 4716 9551 4772
rect 9607 4716 9632 4772
rect 9688 4716 9713 4772
rect 9769 4716 14858 4772
rect 7578 4692 14858 4716
rect 7578 4636 7587 4692
rect 7643 4636 7669 4692
rect 7725 4636 7751 4692
rect 7807 4636 7833 4692
rect 7889 4636 7915 4692
rect 7971 4636 7997 4692
rect 8053 4636 8079 4692
rect 8135 4636 8161 4692
rect 8217 4636 8243 4692
rect 8299 4636 8325 4692
rect 8381 4636 8407 4692
rect 8463 4636 8489 4692
rect 8545 4636 8571 4692
rect 8627 4636 8653 4692
rect 8709 4636 8735 4692
rect 8791 4636 8817 4692
rect 8873 4636 8899 4692
rect 8955 4636 8981 4692
rect 9037 4636 9063 4692
rect 9119 4636 9145 4692
rect 9201 4636 9227 4692
rect 9283 4636 9308 4692
rect 9364 4636 9389 4692
rect 9445 4636 9470 4692
rect 9526 4636 9551 4692
rect 9607 4636 9632 4692
rect 9688 4636 9713 4692
rect 9769 4636 14858 4692
rect 7578 4612 14858 4636
rect 7578 4556 7587 4612
rect 7643 4556 7669 4612
rect 7725 4556 7751 4612
rect 7807 4556 7833 4612
rect 7889 4556 7915 4612
rect 7971 4556 7997 4612
rect 8053 4556 8079 4612
rect 8135 4556 8161 4612
rect 8217 4556 8243 4612
rect 8299 4556 8325 4612
rect 8381 4556 8407 4612
rect 8463 4556 8489 4612
rect 8545 4556 8571 4612
rect 8627 4556 8653 4612
rect 8709 4556 8735 4612
rect 8791 4556 8817 4612
rect 8873 4556 8899 4612
rect 8955 4556 8981 4612
rect 9037 4556 9063 4612
rect 9119 4556 9145 4612
rect 9201 4556 9227 4612
rect 9283 4556 9308 4612
rect 9364 4556 9389 4612
rect 9445 4556 9470 4612
rect 9526 4556 9551 4612
rect 9607 4556 9632 4612
rect 9688 4556 9713 4612
rect 9769 4556 14858 4612
rect 7578 4532 14858 4556
rect 7578 4476 7587 4532
rect 7643 4476 7669 4532
rect 7725 4476 7751 4532
rect 7807 4476 7833 4532
rect 7889 4476 7915 4532
rect 7971 4476 7997 4532
rect 8053 4476 8079 4532
rect 8135 4476 8161 4532
rect 8217 4476 8243 4532
rect 8299 4476 8325 4532
rect 8381 4476 8407 4532
rect 8463 4476 8489 4532
rect 8545 4476 8571 4532
rect 8627 4476 8653 4532
rect 8709 4476 8735 4532
rect 8791 4476 8817 4532
rect 8873 4476 8899 4532
rect 8955 4476 8981 4532
rect 9037 4476 9063 4532
rect 9119 4476 9145 4532
rect 9201 4476 9227 4532
rect 9283 4476 9308 4532
rect 9364 4476 9389 4532
rect 9445 4476 9470 4532
rect 9526 4476 9551 4532
rect 9607 4476 9632 4532
rect 9688 4476 9713 4532
rect 9769 4476 14858 4532
rect 7578 4452 14858 4476
rect 7578 4396 7587 4452
rect 7643 4396 7669 4452
rect 7725 4396 7751 4452
rect 7807 4396 7833 4452
rect 7889 4396 7915 4452
rect 7971 4396 7997 4452
rect 8053 4396 8079 4452
rect 8135 4396 8161 4452
rect 8217 4396 8243 4452
rect 8299 4396 8325 4452
rect 8381 4396 8407 4452
rect 8463 4396 8489 4452
rect 8545 4396 8571 4452
rect 8627 4396 8653 4452
rect 8709 4396 8735 4452
rect 8791 4396 8817 4452
rect 8873 4396 8899 4452
rect 8955 4396 8981 4452
rect 9037 4396 9063 4452
rect 9119 4396 9145 4452
rect 9201 4396 9227 4452
rect 9283 4396 9308 4452
rect 9364 4396 9389 4452
rect 9445 4396 9470 4452
rect 9526 4396 9551 4452
rect 9607 4396 9632 4452
rect 9688 4396 9713 4452
rect 9769 4396 14858 4452
rect 7578 4372 14858 4396
rect 7578 4316 7587 4372
rect 7643 4316 7669 4372
rect 7725 4316 7751 4372
rect 7807 4316 7833 4372
rect 7889 4316 7915 4372
rect 7971 4316 7997 4372
rect 8053 4316 8079 4372
rect 8135 4316 8161 4372
rect 8217 4316 8243 4372
rect 8299 4316 8325 4372
rect 8381 4316 8407 4372
rect 8463 4316 8489 4372
rect 8545 4316 8571 4372
rect 8627 4316 8653 4372
rect 8709 4316 8735 4372
rect 8791 4316 8817 4372
rect 8873 4316 8899 4372
rect 8955 4316 8981 4372
rect 9037 4316 9063 4372
rect 9119 4316 9145 4372
rect 9201 4316 9227 4372
rect 9283 4316 9308 4372
rect 9364 4316 9389 4372
rect 9445 4316 9470 4372
rect 9526 4316 9551 4372
rect 9607 4316 9632 4372
rect 9688 4316 9713 4372
rect 9769 4316 14858 4372
rect 7578 4292 14858 4316
rect 7578 4236 7587 4292
rect 7643 4236 7669 4292
rect 7725 4236 7751 4292
rect 7807 4236 7833 4292
rect 7889 4236 7915 4292
rect 7971 4236 7997 4292
rect 8053 4236 8079 4292
rect 8135 4236 8161 4292
rect 8217 4236 8243 4292
rect 8299 4236 8325 4292
rect 8381 4236 8407 4292
rect 8463 4236 8489 4292
rect 8545 4236 8571 4292
rect 8627 4236 8653 4292
rect 8709 4236 8735 4292
rect 8791 4236 8817 4292
rect 8873 4236 8899 4292
rect 8955 4236 8981 4292
rect 9037 4236 9063 4292
rect 9119 4236 9145 4292
rect 9201 4236 9227 4292
rect 9283 4236 9308 4292
rect 9364 4236 9389 4292
rect 9445 4236 9470 4292
rect 9526 4236 9551 4292
rect 9607 4236 9632 4292
rect 9688 4236 9713 4292
rect 9769 4236 14858 4292
rect 7578 4212 14858 4236
rect 7578 4156 7587 4212
rect 7643 4156 7669 4212
rect 7725 4156 7751 4212
rect 7807 4156 7833 4212
rect 7889 4156 7915 4212
rect 7971 4156 7997 4212
rect 8053 4156 8079 4212
rect 8135 4156 8161 4212
rect 8217 4156 8243 4212
rect 8299 4156 8325 4212
rect 8381 4156 8407 4212
rect 8463 4156 8489 4212
rect 8545 4156 8571 4212
rect 8627 4156 8653 4212
rect 8709 4156 8735 4212
rect 8791 4156 8817 4212
rect 8873 4156 8899 4212
rect 8955 4156 8981 4212
rect 9037 4156 9063 4212
rect 9119 4156 9145 4212
rect 9201 4156 9227 4212
rect 9283 4156 9308 4212
rect 9364 4156 9389 4212
rect 9445 4156 9470 4212
rect 9526 4156 9551 4212
rect 9607 4156 9632 4212
rect 9688 4156 9713 4212
rect 9769 4156 14858 4212
rect 7578 4132 14858 4156
rect 7578 4076 7587 4132
rect 7643 4076 7669 4132
rect 7725 4076 7751 4132
rect 7807 4076 7833 4132
rect 7889 4076 7915 4132
rect 7971 4076 7997 4132
rect 8053 4076 8079 4132
rect 8135 4076 8161 4132
rect 8217 4076 8243 4132
rect 8299 4076 8325 4132
rect 8381 4076 8407 4132
rect 8463 4076 8489 4132
rect 8545 4076 8571 4132
rect 8627 4076 8653 4132
rect 8709 4076 8735 4132
rect 8791 4076 8817 4132
rect 8873 4076 8899 4132
rect 8955 4076 8981 4132
rect 9037 4076 9063 4132
rect 9119 4076 9145 4132
rect 9201 4076 9227 4132
rect 9283 4076 9308 4132
rect 9364 4076 9389 4132
rect 9445 4076 9470 4132
rect 9526 4076 9551 4132
rect 9607 4076 9632 4132
rect 9688 4076 9713 4132
rect 9769 4076 14858 4132
rect 7578 4052 14858 4076
rect 7578 3996 7587 4052
rect 7643 3996 7669 4052
rect 7725 3996 7751 4052
rect 7807 3996 7833 4052
rect 7889 3996 7915 4052
rect 7971 3996 7997 4052
rect 8053 3996 8079 4052
rect 8135 3996 8161 4052
rect 8217 3996 8243 4052
rect 8299 3996 8325 4052
rect 8381 3996 8407 4052
rect 8463 3996 8489 4052
rect 8545 3996 8571 4052
rect 8627 3996 8653 4052
rect 8709 3996 8735 4052
rect 8791 3996 8817 4052
rect 8873 3996 8899 4052
rect 8955 3996 8981 4052
rect 9037 3996 9063 4052
rect 9119 3996 9145 4052
rect 9201 3996 9227 4052
rect 9283 3996 9308 4052
rect 9364 3996 9389 4052
rect 9445 3996 9470 4052
rect 9526 3996 9551 4052
rect 9607 3996 9632 4052
rect 9688 3996 9713 4052
rect 9769 3996 14858 4052
rect 7578 3972 14858 3996
rect 7578 3916 7587 3972
rect 7643 3916 7669 3972
rect 7725 3916 7751 3972
rect 7807 3916 7833 3972
rect 7889 3916 7915 3972
rect 7971 3916 7997 3972
rect 8053 3916 8079 3972
rect 8135 3916 8161 3972
rect 8217 3916 8243 3972
rect 8299 3916 8325 3972
rect 8381 3916 8407 3972
rect 8463 3916 8489 3972
rect 8545 3916 8571 3972
rect 8627 3916 8653 3972
rect 8709 3916 8735 3972
rect 8791 3916 8817 3972
rect 8873 3916 8899 3972
rect 8955 3916 8981 3972
rect 9037 3916 9063 3972
rect 9119 3916 9145 3972
rect 9201 3916 9227 3972
rect 9283 3916 9308 3972
rect 9364 3916 9389 3972
rect 9445 3916 9470 3972
rect 9526 3916 9551 3972
rect 9607 3916 9632 3972
rect 9688 3916 9713 3972
rect 9769 3916 14858 3972
rect 7578 3892 14858 3916
rect 7578 3836 7587 3892
rect 7643 3836 7669 3892
rect 7725 3836 7751 3892
rect 7807 3836 7833 3892
rect 7889 3836 7915 3892
rect 7971 3836 7997 3892
rect 8053 3836 8079 3892
rect 8135 3836 8161 3892
rect 8217 3836 8243 3892
rect 8299 3836 8325 3892
rect 8381 3836 8407 3892
rect 8463 3836 8489 3892
rect 8545 3836 8571 3892
rect 8627 3836 8653 3892
rect 8709 3836 8735 3892
rect 8791 3836 8817 3892
rect 8873 3836 8899 3892
rect 8955 3836 8981 3892
rect 9037 3836 9063 3892
rect 9119 3836 9145 3892
rect 9201 3836 9227 3892
rect 9283 3836 9308 3892
rect 9364 3836 9389 3892
rect 9445 3836 9470 3892
rect 9526 3836 9551 3892
rect 9607 3836 9632 3892
rect 9688 3836 9713 3892
rect 9769 3836 14858 3892
rect 7578 3812 14858 3836
rect 7578 3756 7587 3812
rect 7643 3756 7669 3812
rect 7725 3756 7751 3812
rect 7807 3756 7833 3812
rect 7889 3756 7915 3812
rect 7971 3756 7997 3812
rect 8053 3756 8079 3812
rect 8135 3756 8161 3812
rect 8217 3756 8243 3812
rect 8299 3756 8325 3812
rect 8381 3756 8407 3812
rect 8463 3756 8489 3812
rect 8545 3756 8571 3812
rect 8627 3756 8653 3812
rect 8709 3756 8735 3812
rect 8791 3756 8817 3812
rect 8873 3756 8899 3812
rect 8955 3756 8981 3812
rect 9037 3756 9063 3812
rect 9119 3756 9145 3812
rect 9201 3756 9227 3812
rect 9283 3756 9308 3812
rect 9364 3756 9389 3812
rect 9445 3756 9470 3812
rect 9526 3756 9551 3812
rect 9607 3756 9632 3812
rect 9688 3756 9713 3812
rect 9769 3756 14858 3812
rect 7578 3732 14858 3756
rect 7578 3676 7587 3732
rect 7643 3676 7669 3732
rect 7725 3676 7751 3732
rect 7807 3676 7833 3732
rect 7889 3676 7915 3732
rect 7971 3676 7997 3732
rect 8053 3676 8079 3732
rect 8135 3676 8161 3732
rect 8217 3676 8243 3732
rect 8299 3676 8325 3732
rect 8381 3676 8407 3732
rect 8463 3676 8489 3732
rect 8545 3676 8571 3732
rect 8627 3676 8653 3732
rect 8709 3676 8735 3732
rect 8791 3676 8817 3732
rect 8873 3676 8899 3732
rect 8955 3676 8981 3732
rect 9037 3676 9063 3732
rect 9119 3676 9145 3732
rect 9201 3676 9227 3732
rect 9283 3676 9308 3732
rect 9364 3676 9389 3732
rect 9445 3676 9470 3732
rect 9526 3676 9551 3732
rect 9607 3676 9632 3732
rect 9688 3676 9713 3732
rect 9769 3676 14858 3732
rect 7578 3652 14858 3676
rect 7578 3596 7587 3652
rect 7643 3596 7669 3652
rect 7725 3596 7751 3652
rect 7807 3596 7833 3652
rect 7889 3596 7915 3652
rect 7971 3596 7997 3652
rect 8053 3596 8079 3652
rect 8135 3596 8161 3652
rect 8217 3596 8243 3652
rect 8299 3596 8325 3652
rect 8381 3596 8407 3652
rect 8463 3596 8489 3652
rect 8545 3596 8571 3652
rect 8627 3596 8653 3652
rect 8709 3596 8735 3652
rect 8791 3596 8817 3652
rect 8873 3596 8899 3652
rect 8955 3596 8981 3652
rect 9037 3596 9063 3652
rect 9119 3596 9145 3652
rect 9201 3596 9227 3652
rect 9283 3596 9308 3652
rect 9364 3596 9389 3652
rect 9445 3596 9470 3652
rect 9526 3596 9551 3652
rect 9607 3596 9632 3652
rect 9688 3596 9713 3652
rect 9769 3596 14858 3652
rect 7578 3572 14858 3596
rect 7578 3516 7587 3572
rect 7643 3516 7669 3572
rect 7725 3516 7751 3572
rect 7807 3516 7833 3572
rect 7889 3516 7915 3572
rect 7971 3516 7997 3572
rect 8053 3516 8079 3572
rect 8135 3516 8161 3572
rect 8217 3516 8243 3572
rect 8299 3516 8325 3572
rect 8381 3516 8407 3572
rect 8463 3516 8489 3572
rect 8545 3516 8571 3572
rect 8627 3516 8653 3572
rect 8709 3516 8735 3572
rect 8791 3516 8817 3572
rect 8873 3516 8899 3572
rect 8955 3516 8981 3572
rect 9037 3516 9063 3572
rect 9119 3516 9145 3572
rect 9201 3516 9227 3572
rect 9283 3516 9308 3572
rect 9364 3516 9389 3572
rect 9445 3516 9470 3572
rect 9526 3516 9551 3572
rect 9607 3516 9632 3572
rect 9688 3516 9713 3572
rect 9769 3516 14858 3572
rect 7578 3492 14858 3516
rect 7578 3436 7587 3492
rect 7643 3436 7669 3492
rect 7725 3436 7751 3492
rect 7807 3436 7833 3492
rect 7889 3436 7915 3492
rect 7971 3436 7997 3492
rect 8053 3436 8079 3492
rect 8135 3436 8161 3492
rect 8217 3436 8243 3492
rect 8299 3436 8325 3492
rect 8381 3436 8407 3492
rect 8463 3436 8489 3492
rect 8545 3436 8571 3492
rect 8627 3436 8653 3492
rect 8709 3436 8735 3492
rect 8791 3436 8817 3492
rect 8873 3436 8899 3492
rect 8955 3436 8981 3492
rect 9037 3436 9063 3492
rect 9119 3436 9145 3492
rect 9201 3436 9227 3492
rect 9283 3436 9308 3492
rect 9364 3436 9389 3492
rect 9445 3436 9470 3492
rect 9526 3436 9551 3492
rect 9607 3436 9632 3492
rect 9688 3436 9713 3492
rect 9769 3436 14858 3492
rect 7578 3412 14858 3436
rect 7578 3356 7587 3412
rect 7643 3356 7669 3412
rect 7725 3356 7751 3412
rect 7807 3356 7833 3412
rect 7889 3356 7915 3412
rect 7971 3356 7997 3412
rect 8053 3356 8079 3412
rect 8135 3356 8161 3412
rect 8217 3356 8243 3412
rect 8299 3356 8325 3412
rect 8381 3356 8407 3412
rect 8463 3356 8489 3412
rect 8545 3356 8571 3412
rect 8627 3356 8653 3412
rect 8709 3356 8735 3412
rect 8791 3356 8817 3412
rect 8873 3356 8899 3412
rect 8955 3356 8981 3412
rect 9037 3356 9063 3412
rect 9119 3356 9145 3412
rect 9201 3356 9227 3412
rect 9283 3356 9308 3412
rect 9364 3356 9389 3412
rect 9445 3356 9470 3412
rect 9526 3356 9551 3412
rect 9607 3356 9632 3412
rect 9688 3356 9713 3412
rect 9769 3356 14858 3412
rect 7578 3332 14858 3356
rect 7578 3276 7587 3332
rect 7643 3276 7669 3332
rect 7725 3276 7751 3332
rect 7807 3276 7833 3332
rect 7889 3276 7915 3332
rect 7971 3276 7997 3332
rect 8053 3276 8079 3332
rect 8135 3276 8161 3332
rect 8217 3276 8243 3332
rect 8299 3276 8325 3332
rect 8381 3276 8407 3332
rect 8463 3276 8489 3332
rect 8545 3276 8571 3332
rect 8627 3276 8653 3332
rect 8709 3276 8735 3332
rect 8791 3276 8817 3332
rect 8873 3276 8899 3332
rect 8955 3276 8981 3332
rect 9037 3276 9063 3332
rect 9119 3276 9145 3332
rect 9201 3276 9227 3332
rect 9283 3276 9308 3332
rect 9364 3276 9389 3332
rect 9445 3276 9470 3332
rect 9526 3276 9551 3332
rect 9607 3276 9632 3332
rect 9688 3276 9713 3332
rect 9769 3276 14858 3332
rect 7578 3252 14858 3276
rect 7578 3196 7587 3252
rect 7643 3196 7669 3252
rect 7725 3196 7751 3252
rect 7807 3196 7833 3252
rect 7889 3196 7915 3252
rect 7971 3196 7997 3252
rect 8053 3196 8079 3252
rect 8135 3196 8161 3252
rect 8217 3196 8243 3252
rect 8299 3196 8325 3252
rect 8381 3196 8407 3252
rect 8463 3196 8489 3252
rect 8545 3196 8571 3252
rect 8627 3196 8653 3252
rect 8709 3196 8735 3252
rect 8791 3196 8817 3252
rect 8873 3196 8899 3252
rect 8955 3196 8981 3252
rect 9037 3196 9063 3252
rect 9119 3196 9145 3252
rect 9201 3196 9227 3252
rect 9283 3196 9308 3252
rect 9364 3196 9389 3252
rect 9445 3196 9470 3252
rect 9526 3196 9551 3252
rect 9607 3196 9632 3252
rect 9688 3196 9713 3252
rect 9769 3196 14858 3252
rect 7578 3172 14858 3196
rect 7578 3116 7587 3172
rect 7643 3116 7669 3172
rect 7725 3116 7751 3172
rect 7807 3116 7833 3172
rect 7889 3116 7915 3172
rect 7971 3116 7997 3172
rect 8053 3116 8079 3172
rect 8135 3116 8161 3172
rect 8217 3116 8243 3172
rect 8299 3116 8325 3172
rect 8381 3116 8407 3172
rect 8463 3116 8489 3172
rect 8545 3116 8571 3172
rect 8627 3116 8653 3172
rect 8709 3116 8735 3172
rect 8791 3116 8817 3172
rect 8873 3116 8899 3172
rect 8955 3116 8981 3172
rect 9037 3116 9063 3172
rect 9119 3116 9145 3172
rect 9201 3116 9227 3172
rect 9283 3116 9308 3172
rect 9364 3116 9389 3172
rect 9445 3116 9470 3172
rect 9526 3116 9551 3172
rect 9607 3116 9632 3172
rect 9688 3116 9713 3172
rect 9769 3116 14858 3172
rect 7578 3092 14858 3116
rect 7578 3036 7587 3092
rect 7643 3036 7669 3092
rect 7725 3036 7751 3092
rect 7807 3036 7833 3092
rect 7889 3036 7915 3092
rect 7971 3036 7997 3092
rect 8053 3036 8079 3092
rect 8135 3036 8161 3092
rect 8217 3036 8243 3092
rect 8299 3036 8325 3092
rect 8381 3036 8407 3092
rect 8463 3036 8489 3092
rect 8545 3036 8571 3092
rect 8627 3036 8653 3092
rect 8709 3036 8735 3092
rect 8791 3036 8817 3092
rect 8873 3036 8899 3092
rect 8955 3036 8981 3092
rect 9037 3036 9063 3092
rect 9119 3036 9145 3092
rect 9201 3036 9227 3092
rect 9283 3036 9308 3092
rect 9364 3036 9389 3092
rect 9445 3036 9470 3092
rect 9526 3036 9551 3092
rect 9607 3036 9632 3092
rect 9688 3036 9713 3092
rect 9769 3036 14858 3092
rect 7578 3012 14858 3036
rect 7578 2956 7587 3012
rect 7643 2956 7669 3012
rect 7725 2956 7751 3012
rect 7807 2956 7833 3012
rect 7889 2956 7915 3012
rect 7971 2956 7997 3012
rect 8053 2956 8079 3012
rect 8135 2956 8161 3012
rect 8217 2956 8243 3012
rect 8299 2956 8325 3012
rect 8381 2956 8407 3012
rect 8463 2956 8489 3012
rect 8545 2956 8571 3012
rect 8627 2956 8653 3012
rect 8709 2956 8735 3012
rect 8791 2956 8817 3012
rect 8873 2956 8899 3012
rect 8955 2956 8981 3012
rect 9037 2956 9063 3012
rect 9119 2956 9145 3012
rect 9201 2956 9227 3012
rect 9283 2956 9308 3012
rect 9364 2956 9389 3012
rect 9445 2956 9470 3012
rect 9526 2956 9551 3012
rect 9607 2956 9632 3012
rect 9688 2956 9713 3012
rect 9769 2956 14858 3012
rect 7578 2932 14858 2956
rect 7578 2876 7587 2932
rect 7643 2876 7669 2932
rect 7725 2876 7751 2932
rect 7807 2876 7833 2932
rect 7889 2876 7915 2932
rect 7971 2876 7997 2932
rect 8053 2876 8079 2932
rect 8135 2876 8161 2932
rect 8217 2876 8243 2932
rect 8299 2876 8325 2932
rect 8381 2876 8407 2932
rect 8463 2876 8489 2932
rect 8545 2876 8571 2932
rect 8627 2876 8653 2932
rect 8709 2876 8735 2932
rect 8791 2876 8817 2932
rect 8873 2876 8899 2932
rect 8955 2876 8981 2932
rect 9037 2876 9063 2932
rect 9119 2876 9145 2932
rect 9201 2876 9227 2932
rect 9283 2876 9308 2932
rect 9364 2876 9389 2932
rect 9445 2876 9470 2932
rect 9526 2876 9551 2932
rect 9607 2876 9632 2932
rect 9688 2876 9713 2932
rect 9769 2876 14858 2932
rect 7578 2852 14858 2876
rect 7578 2796 7587 2852
rect 7643 2796 7669 2852
rect 7725 2796 7751 2852
rect 7807 2796 7833 2852
rect 7889 2796 7915 2852
rect 7971 2796 7997 2852
rect 8053 2796 8079 2852
rect 8135 2796 8161 2852
rect 8217 2796 8243 2852
rect 8299 2796 8325 2852
rect 8381 2796 8407 2852
rect 8463 2796 8489 2852
rect 8545 2796 8571 2852
rect 8627 2796 8653 2852
rect 8709 2796 8735 2852
rect 8791 2796 8817 2852
rect 8873 2796 8899 2852
rect 8955 2796 8981 2852
rect 9037 2796 9063 2852
rect 9119 2796 9145 2852
rect 9201 2796 9227 2852
rect 9283 2796 9308 2852
rect 9364 2796 9389 2852
rect 9445 2796 9470 2852
rect 9526 2796 9551 2852
rect 9607 2796 9632 2852
rect 9688 2796 9713 2852
rect 9769 2796 14858 2852
rect 7578 2772 14858 2796
rect 7578 2716 7587 2772
rect 7643 2716 7669 2772
rect 7725 2716 7751 2772
rect 7807 2716 7833 2772
rect 7889 2716 7915 2772
rect 7971 2716 7997 2772
rect 8053 2716 8079 2772
rect 8135 2716 8161 2772
rect 8217 2716 8243 2772
rect 8299 2716 8325 2772
rect 8381 2716 8407 2772
rect 8463 2716 8489 2772
rect 8545 2716 8571 2772
rect 8627 2716 8653 2772
rect 8709 2716 8735 2772
rect 8791 2716 8817 2772
rect 8873 2716 8899 2772
rect 8955 2716 8981 2772
rect 9037 2716 9063 2772
rect 9119 2716 9145 2772
rect 9201 2716 9227 2772
rect 9283 2716 9308 2772
rect 9364 2716 9389 2772
rect 9445 2716 9470 2772
rect 9526 2716 9551 2772
rect 9607 2716 9632 2772
rect 9688 2716 9713 2772
rect 9769 2716 14858 2772
rect 7578 2692 14858 2716
rect 7578 2636 7587 2692
rect 7643 2636 7669 2692
rect 7725 2636 7751 2692
rect 7807 2636 7833 2692
rect 7889 2636 7915 2692
rect 7971 2636 7997 2692
rect 8053 2636 8079 2692
rect 8135 2636 8161 2692
rect 8217 2636 8243 2692
rect 8299 2636 8325 2692
rect 8381 2636 8407 2692
rect 8463 2636 8489 2692
rect 8545 2636 8571 2692
rect 8627 2636 8653 2692
rect 8709 2636 8735 2692
rect 8791 2636 8817 2692
rect 8873 2636 8899 2692
rect 8955 2636 8981 2692
rect 9037 2636 9063 2692
rect 9119 2636 9145 2692
rect 9201 2636 9227 2692
rect 9283 2636 9308 2692
rect 9364 2636 9389 2692
rect 9445 2636 9470 2692
rect 9526 2636 9551 2692
rect 9607 2636 9632 2692
rect 9688 2636 9713 2692
rect 9769 2636 14858 2692
rect 7578 2612 14858 2636
rect 7578 2556 7587 2612
rect 7643 2556 7669 2612
rect 7725 2556 7751 2612
rect 7807 2556 7833 2612
rect 7889 2556 7915 2612
rect 7971 2556 7997 2612
rect 8053 2556 8079 2612
rect 8135 2556 8161 2612
rect 8217 2556 8243 2612
rect 8299 2556 8325 2612
rect 8381 2556 8407 2612
rect 8463 2556 8489 2612
rect 8545 2556 8571 2612
rect 8627 2556 8653 2612
rect 8709 2556 8735 2612
rect 8791 2556 8817 2612
rect 8873 2556 8899 2612
rect 8955 2556 8981 2612
rect 9037 2556 9063 2612
rect 9119 2556 9145 2612
rect 9201 2556 9227 2612
rect 9283 2556 9308 2612
rect 9364 2556 9389 2612
rect 9445 2556 9470 2612
rect 9526 2556 9551 2612
rect 9607 2556 9632 2612
rect 9688 2556 9713 2612
rect 9769 2556 14858 2612
rect 7578 2532 14858 2556
rect 4873 2476 4879 2480
rect 187 2462 4879 2476
rect 187 2410 2766 2462
rect 2818 2410 2831 2462
rect 2883 2410 2896 2462
rect 2948 2410 2961 2462
rect 3013 2410 3026 2462
rect 3078 2410 3091 2462
rect 3143 2410 3156 2462
rect 3208 2410 3221 2462
rect 3273 2410 3285 2462
rect 3337 2410 3349 2462
rect 3401 2410 3413 2462
rect 3465 2410 3477 2462
rect 3529 2410 3541 2462
rect 3593 2410 3605 2462
rect 3657 2410 3669 2462
rect 3721 2410 3733 2462
rect 3785 2410 3797 2462
rect 3849 2410 3861 2462
rect 3913 2410 3925 2462
rect 3977 2410 3989 2462
rect 4041 2410 4053 2462
rect 4105 2410 4117 2462
rect 4169 2410 4181 2462
rect 4233 2410 4245 2462
rect 4297 2410 4309 2462
rect 4361 2410 4373 2462
rect 4425 2410 4437 2462
rect 4489 2410 4501 2462
rect 4553 2410 4565 2462
rect 4617 2410 4629 2462
rect 4681 2410 4693 2462
rect 4745 2410 4757 2462
rect 4809 2410 4821 2462
rect 4873 2410 4879 2462
rect 187 2396 4879 2410
rect 187 2344 2766 2396
rect 2818 2344 2831 2396
rect 2883 2344 2896 2396
rect 2948 2344 2961 2396
rect 3013 2344 3026 2396
rect 3078 2344 3091 2396
rect 3143 2344 3156 2396
rect 3208 2344 3221 2396
rect 3273 2344 3285 2396
rect 3337 2344 3349 2396
rect 3401 2344 3413 2396
rect 3465 2344 3477 2396
rect 3529 2344 3541 2396
rect 3593 2344 3605 2396
rect 3657 2344 3669 2396
rect 3721 2344 3733 2396
rect 3785 2344 3797 2396
rect 3849 2344 3861 2396
rect 3913 2344 3925 2396
rect 3977 2344 3989 2396
rect 4041 2344 4053 2396
rect 4105 2344 4117 2396
rect 4169 2344 4181 2396
rect 4233 2344 4245 2396
rect 4297 2344 4309 2396
rect 4361 2344 4373 2396
rect 4425 2344 4437 2396
rect 4489 2344 4501 2396
rect 4553 2344 4565 2396
rect 4617 2344 4629 2396
rect 4681 2344 4693 2396
rect 4745 2344 4757 2396
rect 4809 2344 4821 2396
rect 4873 2344 4879 2396
rect 187 2330 4879 2344
rect 187 2278 2766 2330
rect 2818 2278 2831 2330
rect 2883 2278 2896 2330
rect 2948 2278 2961 2330
rect 3013 2278 3026 2330
rect 3078 2278 3091 2330
rect 3143 2278 3156 2330
rect 3208 2278 3221 2330
rect 3273 2278 3285 2330
rect 3337 2278 3349 2330
rect 3401 2278 3413 2330
rect 3465 2278 3477 2330
rect 3529 2278 3541 2330
rect 3593 2278 3605 2330
rect 3657 2278 3669 2330
rect 3721 2278 3733 2330
rect 3785 2278 3797 2330
rect 3849 2278 3861 2330
rect 3913 2278 3925 2330
rect 3977 2278 3989 2330
rect 4041 2278 4053 2330
rect 4105 2278 4117 2330
rect 4169 2278 4181 2330
rect 4233 2278 4245 2330
rect 4297 2278 4309 2330
rect 4361 2278 4373 2330
rect 4425 2278 4437 2330
rect 4489 2278 4501 2330
rect 4553 2278 4565 2330
rect 4617 2278 4629 2330
rect 4681 2278 4693 2330
rect 4745 2278 4757 2330
rect 4809 2278 4821 2330
rect 4873 2278 4879 2330
rect 187 2264 4879 2278
rect 187 2212 2766 2264
rect 2818 2212 2831 2264
rect 2883 2212 2896 2264
rect 2948 2212 2961 2264
rect 3013 2212 3026 2264
rect 3078 2212 3091 2264
rect 3143 2212 3156 2264
rect 3208 2212 3221 2264
rect 3273 2212 3285 2264
rect 3337 2212 3349 2264
rect 3401 2212 3413 2264
rect 3465 2212 3477 2264
rect 3529 2212 3541 2264
rect 3593 2212 3605 2264
rect 3657 2212 3669 2264
rect 3721 2212 3733 2264
rect 3785 2212 3797 2264
rect 3849 2212 3861 2264
rect 3913 2212 3925 2264
rect 3977 2212 3989 2264
rect 4041 2212 4053 2264
rect 4105 2212 4117 2264
rect 4169 2212 4181 2264
rect 4233 2212 4245 2264
rect 4297 2212 4309 2264
rect 4361 2212 4373 2264
rect 4425 2212 4437 2264
rect 4489 2212 4501 2264
rect 4553 2212 4565 2264
rect 4617 2212 4629 2264
rect 4681 2212 4693 2264
rect 4745 2212 4757 2264
rect 4809 2212 4821 2264
rect 4873 2212 4879 2264
rect 187 1513 4879 2212
tri 4879 1719 5640 2480 nw
rect 7578 2476 7587 2532
rect 7643 2476 7669 2532
rect 7725 2476 7751 2532
rect 7807 2476 7833 2532
rect 7889 2476 7915 2532
rect 7971 2476 7997 2532
rect 8053 2476 8079 2532
rect 8135 2476 8161 2532
rect 8217 2476 8243 2532
rect 8299 2476 8325 2532
rect 8381 2476 8407 2532
rect 8463 2476 8489 2532
rect 8545 2476 8571 2532
rect 8627 2476 8653 2532
rect 8709 2476 8735 2532
rect 8791 2476 8817 2532
rect 8873 2476 8899 2532
rect 8955 2476 8981 2532
rect 9037 2476 9063 2532
rect 9119 2476 9145 2532
rect 9201 2476 9227 2532
rect 9283 2476 9308 2532
rect 9364 2476 9389 2532
rect 9445 2476 9470 2532
rect 9526 2476 9551 2532
rect 9607 2476 9632 2532
rect 9688 2476 9713 2532
rect 9769 2476 14858 2532
rect 7578 2459 14858 2476
tri 9344 1725 10078 2459 ne
rect 187 1461 2776 1513
rect 2828 1461 2842 1513
rect 2894 1461 2908 1513
rect 2960 1461 2974 1513
rect 3026 1461 3040 1513
rect 3092 1461 3106 1513
rect 3158 1461 3172 1513
rect 3224 1461 3238 1513
rect 3290 1461 3304 1513
rect 3356 1461 3370 1513
rect 3422 1461 3436 1513
rect 3488 1461 3502 1513
rect 3554 1461 3568 1513
rect 3620 1461 3634 1513
rect 3686 1461 3700 1513
rect 3752 1461 3766 1513
rect 3818 1461 3832 1513
rect 3884 1461 3898 1513
rect 3950 1461 3964 1513
rect 4016 1461 4030 1513
rect 4082 1461 4096 1513
rect 4148 1461 4162 1513
rect 4214 1461 4228 1513
rect 4280 1461 4294 1513
rect 4346 1461 4360 1513
rect 4412 1461 4426 1513
rect 4478 1461 4492 1513
rect 4544 1461 4558 1513
rect 4610 1461 4624 1513
rect 4676 1461 4690 1513
rect 4742 1461 4756 1513
rect 4808 1461 4821 1513
rect 4873 1461 4879 1513
rect 187 1445 4879 1461
rect 187 1393 2776 1445
rect 2828 1393 2842 1445
rect 2894 1393 2908 1445
rect 2960 1393 2974 1445
rect 3026 1393 3040 1445
rect 3092 1393 3106 1445
rect 3158 1393 3172 1445
rect 3224 1393 3238 1445
rect 3290 1393 3304 1445
rect 3356 1393 3370 1445
rect 3422 1393 3436 1445
rect 3488 1393 3502 1445
rect 3554 1393 3568 1445
rect 3620 1393 3634 1445
rect 3686 1393 3700 1445
rect 3752 1393 3766 1445
rect 3818 1393 3832 1445
rect 3884 1393 3898 1445
rect 3950 1393 3964 1445
rect 4016 1393 4030 1445
rect 4082 1393 4096 1445
rect 4148 1393 4162 1445
rect 4214 1393 4228 1445
rect 4280 1393 4294 1445
rect 4346 1393 4360 1445
rect 4412 1393 4426 1445
rect 4478 1393 4492 1445
rect 4544 1393 4558 1445
rect 4610 1393 4624 1445
rect 4676 1393 4690 1445
rect 4742 1393 4756 1445
rect 4808 1393 4821 1445
rect 4873 1393 4879 1445
rect 187 1377 4879 1393
rect 187 1325 2776 1377
rect 2828 1325 2842 1377
rect 2894 1325 2908 1377
rect 2960 1325 2974 1377
rect 3026 1325 3040 1377
rect 3092 1325 3106 1377
rect 3158 1325 3172 1377
rect 3224 1325 3238 1377
rect 3290 1325 3304 1377
rect 3356 1325 3370 1377
rect 3422 1325 3436 1377
rect 3488 1325 3502 1377
rect 3554 1325 3568 1377
rect 3620 1325 3634 1377
rect 3686 1325 3700 1377
rect 3752 1325 3766 1377
rect 3818 1325 3832 1377
rect 3884 1325 3898 1377
rect 3950 1325 3964 1377
rect 4016 1325 4030 1377
rect 4082 1325 4096 1377
rect 4148 1325 4162 1377
rect 4214 1325 4228 1377
rect 4280 1325 4294 1377
rect 4346 1325 4360 1377
rect 4412 1325 4426 1377
rect 4478 1325 4492 1377
rect 4544 1325 4558 1377
rect 4610 1325 4624 1377
rect 4676 1325 4690 1377
rect 4742 1325 4756 1377
rect 4808 1325 4821 1377
rect 4873 1325 4879 1377
rect 187 1309 4879 1325
rect 187 1257 2776 1309
rect 2828 1257 2842 1309
rect 2894 1257 2908 1309
rect 2960 1257 2974 1309
rect 3026 1257 3040 1309
rect 3092 1257 3106 1309
rect 3158 1257 3172 1309
rect 3224 1257 3238 1309
rect 3290 1257 3304 1309
rect 3356 1257 3370 1309
rect 3422 1257 3436 1309
rect 3488 1257 3502 1309
rect 3554 1257 3568 1309
rect 3620 1257 3634 1309
rect 3686 1257 3700 1309
rect 3752 1257 3766 1309
rect 3818 1257 3832 1309
rect 3884 1257 3898 1309
rect 3950 1257 3964 1309
rect 4016 1257 4030 1309
rect 4082 1257 4096 1309
rect 4148 1257 4162 1309
rect 4214 1257 4228 1309
rect 4280 1257 4294 1309
rect 4346 1257 4360 1309
rect 4412 1257 4426 1309
rect 4478 1257 4492 1309
rect 4544 1257 4558 1309
rect 4610 1257 4624 1309
rect 4676 1257 4690 1309
rect 4742 1257 4756 1309
rect 4808 1257 4821 1309
rect 4873 1257 4879 1309
rect 187 1241 4879 1257
rect 187 1189 2776 1241
rect 2828 1189 2842 1241
rect 2894 1189 2908 1241
rect 2960 1189 2974 1241
rect 3026 1189 3040 1241
rect 3092 1189 3106 1241
rect 3158 1189 3172 1241
rect 3224 1189 3238 1241
rect 3290 1189 3304 1241
rect 3356 1189 3370 1241
rect 3422 1189 3436 1241
rect 3488 1189 3502 1241
rect 3554 1189 3568 1241
rect 3620 1189 3634 1241
rect 3686 1189 3700 1241
rect 3752 1189 3766 1241
rect 3818 1189 3832 1241
rect 3884 1189 3898 1241
rect 3950 1189 3964 1241
rect 4016 1189 4030 1241
rect 4082 1189 4096 1241
rect 4148 1189 4162 1241
rect 4214 1189 4228 1241
rect 4280 1189 4294 1241
rect 4346 1189 4360 1241
rect 4412 1189 4426 1241
rect 4478 1189 4492 1241
rect 4544 1189 4558 1241
rect 4610 1189 4624 1241
rect 4676 1189 4690 1241
rect 4742 1189 4756 1241
rect 4808 1189 4821 1241
rect 4873 1189 4879 1241
rect 187 1173 4879 1189
rect 187 1121 2776 1173
rect 2828 1121 2842 1173
rect 2894 1121 2908 1173
rect 2960 1121 2974 1173
rect 3026 1121 3040 1173
rect 3092 1121 3106 1173
rect 3158 1121 3172 1173
rect 3224 1121 3238 1173
rect 3290 1121 3304 1173
rect 3356 1121 3370 1173
rect 3422 1121 3436 1173
rect 3488 1121 3502 1173
rect 3554 1121 3568 1173
rect 3620 1121 3634 1173
rect 3686 1121 3700 1173
rect 3752 1121 3766 1173
rect 3818 1121 3832 1173
rect 3884 1121 3898 1173
rect 3950 1121 3964 1173
rect 4016 1121 4030 1173
rect 4082 1121 4096 1173
rect 4148 1121 4162 1173
rect 4214 1121 4228 1173
rect 4280 1121 4294 1173
rect 4346 1121 4360 1173
rect 4412 1121 4426 1173
rect 4478 1121 4492 1173
rect 4544 1121 4558 1173
rect 4610 1121 4624 1173
rect 4676 1121 4690 1173
rect 4742 1121 4756 1173
rect 4808 1121 4821 1173
rect 4873 1121 4879 1173
rect 187 1105 4879 1121
rect 187 1053 2776 1105
rect 2828 1053 2842 1105
rect 2894 1053 2908 1105
rect 2960 1053 2974 1105
rect 3026 1053 3040 1105
rect 3092 1053 3106 1105
rect 3158 1053 3172 1105
rect 3224 1053 3238 1105
rect 3290 1053 3304 1105
rect 3356 1053 3370 1105
rect 3422 1053 3436 1105
rect 3488 1053 3502 1105
rect 3554 1053 3568 1105
rect 3620 1053 3634 1105
rect 3686 1053 3700 1105
rect 3752 1053 3766 1105
rect 3818 1053 3832 1105
rect 3884 1053 3898 1105
rect 3950 1053 3964 1105
rect 4016 1053 4030 1105
rect 4082 1053 4096 1105
rect 4148 1053 4162 1105
rect 4214 1053 4228 1105
rect 4280 1053 4294 1105
rect 4346 1053 4360 1105
rect 4412 1053 4426 1105
rect 4478 1053 4492 1105
rect 4544 1053 4558 1105
rect 4610 1053 4624 1105
rect 4676 1053 4690 1105
rect 4742 1053 4756 1105
rect 4808 1053 4821 1105
rect 4873 1053 4879 1105
rect 187 1037 4879 1053
rect 187 985 2776 1037
rect 2828 985 2842 1037
rect 2894 985 2908 1037
rect 2960 985 2974 1037
rect 3026 985 3040 1037
rect 3092 985 3106 1037
rect 3158 985 3172 1037
rect 3224 985 3238 1037
rect 3290 985 3304 1037
rect 3356 985 3370 1037
rect 3422 985 3436 1037
rect 3488 985 3502 1037
rect 3554 985 3568 1037
rect 3620 985 3634 1037
rect 3686 985 3700 1037
rect 3752 985 3766 1037
rect 3818 985 3832 1037
rect 3884 985 3898 1037
rect 3950 985 3964 1037
rect 4016 985 4030 1037
rect 4082 985 4096 1037
rect 4148 985 4162 1037
rect 4214 985 4228 1037
rect 4280 985 4294 1037
rect 4346 985 4360 1037
rect 4412 985 4426 1037
rect 4478 985 4492 1037
rect 4544 985 4558 1037
rect 4610 985 4624 1037
rect 4676 985 4690 1037
rect 4742 985 4756 1037
rect 4808 985 4821 1037
rect 4873 985 4879 1037
tri 99 411 187 499 se
rect 187 411 4879 985
rect 6749 1106 6801 1112
rect 6749 1022 6801 1054
tri 6715 567 6749 601 se
rect 6749 567 6801 970
rect 8703 1106 8755 1112
rect 8703 1022 8755 1054
tri 6801 567 6835 601 sw
tri 8669 567 8703 601 se
rect 8703 567 8755 970
tri 8755 567 8789 601 sw
rect 6701 515 6707 567
rect 6759 515 6791 567
rect 6843 515 6849 567
rect 8655 515 8661 567
rect 8713 515 8745 567
rect 8797 515 8803 567
rect 99 0 4879 411
rect 5179 377 5579 384
rect 5179 325 5190 377
rect 5242 325 5256 377
rect 5308 325 5322 377
rect 5374 325 5388 377
rect 5440 325 5453 377
rect 5505 325 5518 377
rect 5570 325 5579 377
rect 5179 313 5579 325
rect 5179 261 5190 313
rect 5242 261 5256 313
rect 5308 261 5322 313
rect 5374 261 5388 313
rect 5440 261 5453 313
rect 5505 261 5518 313
rect 5570 261 5579 313
rect 5179 249 5579 261
rect 5179 197 5190 249
rect 5242 197 5256 249
rect 5308 197 5322 249
rect 5374 197 5388 249
rect 5440 197 5453 249
rect 5505 197 5518 249
rect 5570 197 5579 249
rect 5179 0 5579 197
rect 10078 0 14858 2459
<< via2 >>
rect 2534 38953 2590 39009
rect 2617 38953 2673 39009
rect 2700 38953 2756 39009
rect 2783 38953 2839 39009
rect 2866 38957 2872 39009
rect 2872 38957 2922 39009
rect 2949 38957 2992 39009
rect 2992 38957 3005 39009
rect 3032 38957 3060 39009
rect 3060 38957 3088 39009
rect 2866 38953 2922 38957
rect 2949 38953 3005 38957
rect 3032 38953 3088 38957
rect 3115 38953 3171 39009
rect 3198 38953 3254 39009
rect 3281 38953 3337 39009
rect 3364 38953 3420 39009
rect 3447 38953 3503 39009
rect 3530 38953 3586 39009
rect 3613 38953 3669 39009
rect 3696 38953 3752 39009
rect 3779 38957 3792 39009
rect 3792 38957 3835 39009
rect 3862 38957 3912 39009
rect 3912 38957 3918 39009
rect 3945 38957 3980 39009
rect 3980 38957 4001 39009
rect 3779 38953 3835 38957
rect 3862 38953 3918 38957
rect 3945 38953 4001 38957
rect 4028 38953 4084 39009
rect 4111 38953 4167 39009
rect 4194 38953 4250 39009
rect 4276 38953 4332 39009
rect 4358 38953 4414 39009
rect 4440 38953 4496 39009
rect 4522 38953 4578 39009
rect 4604 38953 4660 39009
rect 4686 38957 4712 39009
rect 4712 38957 4742 39009
rect 4768 38957 4780 39009
rect 4780 38957 4824 39009
rect 4850 38957 4900 39009
rect 4900 38957 4906 39009
rect 4686 38953 4742 38957
rect 4768 38953 4824 38957
rect 4850 38953 4906 38957
rect 4932 38953 4988 39009
rect 5195 38953 5251 39009
rect 5276 38953 5332 39009
rect 5357 38953 5413 39009
rect 5438 38953 5494 39009
rect 5519 38953 5575 39009
rect 5600 38957 5632 39009
rect 5632 38957 5656 39009
rect 5681 38957 5684 39009
rect 5684 38957 5700 39009
rect 5700 38957 5737 39009
rect 5762 38957 5768 39009
rect 5768 38957 5818 39009
rect 5600 38953 5656 38957
rect 5681 38953 5737 38957
rect 5762 38953 5818 38957
rect 5843 38953 5899 39009
rect 5924 38953 5980 39009
rect 6005 38953 6061 39009
rect 6086 38953 6142 39009
rect 6167 38953 6223 39009
rect 6248 38953 6304 39009
rect 6329 38953 6385 39009
rect 6410 38953 6466 39009
rect 6491 38953 6547 39009
rect 6572 38957 6604 39009
rect 6604 38957 6620 39009
rect 6620 38957 6628 39009
rect 6653 38957 6672 39009
rect 6672 38957 6688 39009
rect 6688 38957 6709 39009
rect 6734 38957 6740 39009
rect 6740 38957 6790 39009
rect 6572 38953 6628 38957
rect 6653 38953 6709 38957
rect 6734 38953 6790 38957
rect 6815 38953 6871 39009
rect 6896 38953 6952 39009
rect 6977 38953 7033 39009
rect 7058 38953 7114 39009
rect 7139 38953 7195 39009
rect 7221 38953 7277 39009
rect 7303 38953 7359 39009
rect 2534 38869 2590 38925
rect 2617 38869 2673 38925
rect 2700 38869 2756 38925
rect 2783 38869 2839 38925
rect 2866 38892 2872 38925
rect 2872 38892 2922 38925
rect 2949 38892 2992 38925
rect 2992 38892 3005 38925
rect 3032 38892 3060 38925
rect 3060 38892 3088 38925
rect 2866 38879 2922 38892
rect 2949 38879 3005 38892
rect 3032 38879 3088 38892
rect 2866 38869 2872 38879
rect 2872 38869 2922 38879
rect 2534 38785 2590 38841
rect 2617 38785 2673 38841
rect 2700 38785 2756 38841
rect 2783 38785 2839 38841
rect 2866 38827 2872 38841
rect 2872 38827 2922 38841
rect 2949 38869 2992 38879
rect 2992 38869 3005 38879
rect 3032 38869 3060 38879
rect 3060 38869 3088 38879
rect 3115 38869 3171 38925
rect 3198 38869 3254 38925
rect 3281 38869 3337 38925
rect 3364 38869 3420 38925
rect 3447 38869 3503 38925
rect 3530 38869 3586 38925
rect 3613 38869 3669 38925
rect 3696 38869 3752 38925
rect 3779 38892 3792 38925
rect 3792 38892 3835 38925
rect 3862 38892 3912 38925
rect 3912 38892 3918 38925
rect 3945 38892 3980 38925
rect 3980 38892 4001 38925
rect 3779 38879 3835 38892
rect 3862 38879 3918 38892
rect 3945 38879 4001 38892
rect 3779 38869 3792 38879
rect 3792 38869 3835 38879
rect 2949 38827 2992 38841
rect 2992 38827 3005 38841
rect 3032 38827 3060 38841
rect 3060 38827 3088 38841
rect 2866 38814 2922 38827
rect 2949 38814 3005 38827
rect 3032 38814 3088 38827
rect 2866 38785 2872 38814
rect 2872 38785 2922 38814
rect 2949 38785 2992 38814
rect 2992 38785 3005 38814
rect 3032 38785 3060 38814
rect 3060 38785 3088 38814
rect 3115 38785 3171 38841
rect 3198 38785 3254 38841
rect 3281 38785 3337 38841
rect 3364 38785 3420 38841
rect 3447 38785 3503 38841
rect 3530 38785 3586 38841
rect 3613 38785 3669 38841
rect 3696 38785 3752 38841
rect 3779 38827 3792 38841
rect 3792 38827 3835 38841
rect 3862 38869 3912 38879
rect 3912 38869 3918 38879
rect 3945 38869 3980 38879
rect 3980 38869 4001 38879
rect 4028 38869 4084 38925
rect 4111 38869 4167 38925
rect 4194 38869 4250 38925
rect 4276 38869 4332 38925
rect 4358 38869 4414 38925
rect 4440 38869 4496 38925
rect 4522 38869 4578 38925
rect 4604 38869 4660 38925
rect 4686 38892 4712 38925
rect 4712 38892 4742 38925
rect 4768 38892 4780 38925
rect 4780 38892 4824 38925
rect 4850 38892 4900 38925
rect 4900 38892 4906 38925
rect 4686 38879 4742 38892
rect 4768 38879 4824 38892
rect 4850 38879 4906 38892
rect 4686 38869 4712 38879
rect 4712 38869 4742 38879
rect 4768 38869 4780 38879
rect 4780 38869 4824 38879
rect 3862 38827 3912 38841
rect 3912 38827 3918 38841
rect 3945 38827 3980 38841
rect 3980 38827 4001 38841
rect 3779 38814 3835 38827
rect 3862 38814 3918 38827
rect 3945 38814 4001 38827
rect 3779 38785 3792 38814
rect 3792 38785 3835 38814
rect 3862 38785 3912 38814
rect 3912 38785 3918 38814
rect 3945 38785 3980 38814
rect 3980 38785 4001 38814
rect 4028 38785 4084 38841
rect 4111 38785 4167 38841
rect 4194 38785 4250 38841
rect 4276 38785 4332 38841
rect 4358 38785 4414 38841
rect 4440 38785 4496 38841
rect 4522 38785 4578 38841
rect 4604 38785 4660 38841
rect 4686 38827 4712 38841
rect 4712 38827 4742 38841
rect 4768 38827 4780 38841
rect 4780 38827 4824 38841
rect 4850 38869 4900 38879
rect 4900 38869 4906 38879
rect 4932 38869 4988 38925
rect 5195 38869 5251 38925
rect 5276 38869 5332 38925
rect 5357 38869 5413 38925
rect 5438 38869 5494 38925
rect 5519 38869 5575 38925
rect 5600 38892 5632 38925
rect 5632 38892 5656 38925
rect 5681 38892 5684 38925
rect 5684 38892 5700 38925
rect 5700 38892 5737 38925
rect 5762 38892 5768 38925
rect 5768 38892 5818 38925
rect 5600 38879 5656 38892
rect 5681 38879 5737 38892
rect 5762 38879 5818 38892
rect 5600 38869 5632 38879
rect 5632 38869 5656 38879
rect 5681 38869 5684 38879
rect 5684 38869 5700 38879
rect 5700 38869 5737 38879
rect 5762 38869 5768 38879
rect 5768 38869 5818 38879
rect 5843 38869 5899 38925
rect 5924 38869 5980 38925
rect 6005 38869 6061 38925
rect 6086 38869 6142 38925
rect 6167 38869 6223 38925
rect 6248 38869 6304 38925
rect 6329 38869 6385 38925
rect 6410 38869 6466 38925
rect 6491 38869 6547 38925
rect 6572 38892 6604 38925
rect 6604 38892 6620 38925
rect 6620 38892 6628 38925
rect 6653 38892 6672 38925
rect 6672 38892 6688 38925
rect 6688 38892 6709 38925
rect 6734 38892 6740 38925
rect 6740 38892 6790 38925
rect 6572 38879 6628 38892
rect 6653 38879 6709 38892
rect 6734 38879 6790 38892
rect 6572 38869 6604 38879
rect 6604 38869 6620 38879
rect 6620 38869 6628 38879
rect 6653 38869 6672 38879
rect 6672 38869 6688 38879
rect 6688 38869 6709 38879
rect 6734 38869 6740 38879
rect 6740 38869 6790 38879
rect 6815 38869 6871 38925
rect 6896 38869 6952 38925
rect 6977 38869 7033 38925
rect 7058 38869 7114 38925
rect 7139 38869 7195 38925
rect 7221 38869 7277 38925
rect 7303 38869 7359 38925
rect 4850 38827 4900 38841
rect 4900 38827 4906 38841
rect 4686 38814 4742 38827
rect 4768 38814 4824 38827
rect 4850 38814 4906 38827
rect 4686 38785 4712 38814
rect 4712 38785 4742 38814
rect 4768 38785 4780 38814
rect 4780 38785 4824 38814
rect 4850 38785 4900 38814
rect 4900 38785 4906 38814
rect 4932 38785 4988 38841
rect 5195 38785 5251 38841
rect 5276 38785 5332 38841
rect 5357 38785 5413 38841
rect 5438 38785 5494 38841
rect 5519 38785 5575 38841
rect 5600 38827 5632 38841
rect 5632 38827 5656 38841
rect 5681 38827 5684 38841
rect 5684 38827 5700 38841
rect 5700 38827 5737 38841
rect 5762 38827 5768 38841
rect 5768 38827 5818 38841
rect 5600 38814 5656 38827
rect 5681 38814 5737 38827
rect 5762 38814 5818 38827
rect 5600 38785 5632 38814
rect 5632 38785 5656 38814
rect 5681 38785 5684 38814
rect 5684 38785 5700 38814
rect 5700 38785 5737 38814
rect 5762 38785 5768 38814
rect 5768 38785 5818 38814
rect 5843 38785 5899 38841
rect 5924 38785 5980 38841
rect 6005 38785 6061 38841
rect 6086 38785 6142 38841
rect 6167 38785 6223 38841
rect 6248 38785 6304 38841
rect 6329 38785 6385 38841
rect 6410 38785 6466 38841
rect 6491 38785 6547 38841
rect 6572 38827 6604 38841
rect 6604 38827 6620 38841
rect 6620 38827 6628 38841
rect 6653 38827 6672 38841
rect 6672 38827 6688 38841
rect 6688 38827 6709 38841
rect 6734 38827 6740 38841
rect 6740 38827 6790 38841
rect 6572 38814 6628 38827
rect 6653 38814 6709 38827
rect 6734 38814 6790 38827
rect 6572 38785 6604 38814
rect 6604 38785 6620 38814
rect 6620 38785 6628 38814
rect 6653 38785 6672 38814
rect 6672 38785 6688 38814
rect 6688 38785 6709 38814
rect 6734 38785 6740 38814
rect 6740 38785 6790 38814
rect 6815 38785 6871 38841
rect 6896 38785 6952 38841
rect 6977 38785 7033 38841
rect 7058 38785 7114 38841
rect 7139 38785 7195 38841
rect 7221 38785 7277 38841
rect 7303 38785 7359 38841
rect 2534 38701 2590 38757
rect 2617 38701 2673 38757
rect 2700 38701 2756 38757
rect 2783 38701 2839 38757
rect 2866 38749 2922 38757
rect 2949 38749 3005 38757
rect 3032 38749 3088 38757
rect 2866 38701 2872 38749
rect 2872 38701 2922 38749
rect 2949 38701 2992 38749
rect 2992 38701 3005 38749
rect 3032 38701 3060 38749
rect 3060 38701 3088 38749
rect 3115 38701 3171 38757
rect 3198 38701 3254 38757
rect 3281 38701 3337 38757
rect 3364 38701 3420 38757
rect 3447 38701 3503 38757
rect 3530 38701 3586 38757
rect 3613 38701 3669 38757
rect 3696 38701 3752 38757
rect 3779 38749 3835 38757
rect 3862 38749 3918 38757
rect 3945 38749 4001 38757
rect 3779 38701 3792 38749
rect 3792 38701 3835 38749
rect 3862 38701 3912 38749
rect 3912 38701 3918 38749
rect 3945 38701 3980 38749
rect 3980 38701 4001 38749
rect 4028 38701 4084 38757
rect 4111 38701 4167 38757
rect 4194 38701 4250 38757
rect 4276 38701 4332 38757
rect 4358 38701 4414 38757
rect 4440 38701 4496 38757
rect 4522 38701 4578 38757
rect 4604 38701 4660 38757
rect 4686 38749 4742 38757
rect 4768 38749 4824 38757
rect 4850 38749 4906 38757
rect 4686 38701 4712 38749
rect 4712 38701 4742 38749
rect 4768 38701 4780 38749
rect 4780 38701 4824 38749
rect 4850 38701 4900 38749
rect 4900 38701 4906 38749
rect 4932 38701 4988 38757
rect 5195 38701 5251 38757
rect 5276 38701 5332 38757
rect 5357 38701 5413 38757
rect 5438 38701 5494 38757
rect 5519 38701 5575 38757
rect 5600 38749 5656 38757
rect 5681 38749 5737 38757
rect 5762 38749 5818 38757
rect 5600 38701 5632 38749
rect 5632 38701 5656 38749
rect 5681 38701 5684 38749
rect 5684 38701 5700 38749
rect 5700 38701 5737 38749
rect 5762 38701 5768 38749
rect 5768 38701 5818 38749
rect 5843 38701 5899 38757
rect 5924 38701 5980 38757
rect 6005 38701 6061 38757
rect 6086 38701 6142 38757
rect 6167 38701 6223 38757
rect 6248 38701 6304 38757
rect 6329 38701 6385 38757
rect 6410 38701 6466 38757
rect 6491 38701 6547 38757
rect 6572 38749 6628 38757
rect 6653 38749 6709 38757
rect 6734 38749 6790 38757
rect 6572 38701 6604 38749
rect 6604 38701 6620 38749
rect 6620 38701 6628 38749
rect 6653 38701 6672 38749
rect 6672 38701 6688 38749
rect 6688 38701 6709 38749
rect 6734 38701 6740 38749
rect 6740 38701 6790 38749
rect 6815 38701 6871 38757
rect 6896 38701 6952 38757
rect 6977 38701 7033 38757
rect 7058 38701 7114 38757
rect 7139 38701 7195 38757
rect 7221 38701 7277 38757
rect 7303 38701 7359 38757
rect 2534 38617 2590 38673
rect 2617 38617 2673 38673
rect 2700 38617 2756 38673
rect 2783 38617 2839 38673
rect 2866 38632 2872 38673
rect 2872 38632 2922 38673
rect 2949 38632 2992 38673
rect 2992 38632 3005 38673
rect 3032 38632 3060 38673
rect 3060 38632 3088 38673
rect 2866 38619 2922 38632
rect 2949 38619 3005 38632
rect 3032 38619 3088 38632
rect 2866 38617 2872 38619
rect 2872 38617 2922 38619
rect 2534 38533 2590 38589
rect 2617 38533 2673 38589
rect 2700 38533 2756 38589
rect 2783 38533 2839 38589
rect 2866 38567 2872 38589
rect 2872 38567 2922 38589
rect 2949 38617 2992 38619
rect 2992 38617 3005 38619
rect 3032 38617 3060 38619
rect 3060 38617 3088 38619
rect 3115 38617 3171 38673
rect 3198 38617 3254 38673
rect 3281 38617 3337 38673
rect 3364 38617 3420 38673
rect 3447 38617 3503 38673
rect 3530 38617 3586 38673
rect 3613 38617 3669 38673
rect 3696 38617 3752 38673
rect 3779 38632 3792 38673
rect 3792 38632 3835 38673
rect 3862 38632 3912 38673
rect 3912 38632 3918 38673
rect 3945 38632 3980 38673
rect 3980 38632 4001 38673
rect 3779 38619 3835 38632
rect 3862 38619 3918 38632
rect 3945 38619 4001 38632
rect 3779 38617 3792 38619
rect 3792 38617 3835 38619
rect 2949 38567 2992 38589
rect 2992 38567 3005 38589
rect 3032 38567 3060 38589
rect 3060 38567 3088 38589
rect 2866 38554 2922 38567
rect 2949 38554 3005 38567
rect 3032 38554 3088 38567
rect 2866 38533 2872 38554
rect 2872 38533 2922 38554
rect 2534 38449 2590 38505
rect 2617 38449 2673 38505
rect 2700 38449 2756 38505
rect 2783 38449 2839 38505
rect 2866 38502 2872 38505
rect 2872 38502 2922 38505
rect 2949 38533 2992 38554
rect 2992 38533 3005 38554
rect 3032 38533 3060 38554
rect 3060 38533 3088 38554
rect 3115 38533 3171 38589
rect 3198 38533 3254 38589
rect 3281 38533 3337 38589
rect 3364 38533 3420 38589
rect 3447 38533 3503 38589
rect 3530 38533 3586 38589
rect 3613 38533 3669 38589
rect 3696 38533 3752 38589
rect 3779 38567 3792 38589
rect 3792 38567 3835 38589
rect 3862 38617 3912 38619
rect 3912 38617 3918 38619
rect 3945 38617 3980 38619
rect 3980 38617 4001 38619
rect 4028 38617 4084 38673
rect 4111 38617 4167 38673
rect 4194 38617 4250 38673
rect 4276 38617 4332 38673
rect 4358 38617 4414 38673
rect 4440 38617 4496 38673
rect 4522 38617 4578 38673
rect 4604 38617 4660 38673
rect 4686 38632 4712 38673
rect 4712 38632 4742 38673
rect 4768 38632 4780 38673
rect 4780 38632 4824 38673
rect 4850 38632 4900 38673
rect 4900 38632 4906 38673
rect 4686 38619 4742 38632
rect 4768 38619 4824 38632
rect 4850 38619 4906 38632
rect 4686 38617 4712 38619
rect 4712 38617 4742 38619
rect 4768 38617 4780 38619
rect 4780 38617 4824 38619
rect 3862 38567 3912 38589
rect 3912 38567 3918 38589
rect 3945 38567 3980 38589
rect 3980 38567 4001 38589
rect 3779 38554 3835 38567
rect 3862 38554 3918 38567
rect 3945 38554 4001 38567
rect 3779 38533 3792 38554
rect 3792 38533 3835 38554
rect 2949 38502 2992 38505
rect 2992 38502 3005 38505
rect 3032 38502 3060 38505
rect 3060 38502 3088 38505
rect 2866 38490 2922 38502
rect 2949 38490 3005 38502
rect 3032 38490 3088 38502
rect 2866 38449 2872 38490
rect 2872 38449 2922 38490
rect 2949 38449 2992 38490
rect 2992 38449 3005 38490
rect 3032 38449 3060 38490
rect 3060 38449 3088 38490
rect 3115 38449 3171 38505
rect 3198 38449 3254 38505
rect 3281 38449 3337 38505
rect 3364 38449 3420 38505
rect 3447 38449 3503 38505
rect 3530 38449 3586 38505
rect 3613 38449 3669 38505
rect 3696 38449 3752 38505
rect 3779 38502 3792 38505
rect 3792 38502 3835 38505
rect 3862 38533 3912 38554
rect 3912 38533 3918 38554
rect 3945 38533 3980 38554
rect 3980 38533 4001 38554
rect 4028 38533 4084 38589
rect 4111 38533 4167 38589
rect 4194 38533 4250 38589
rect 4276 38533 4332 38589
rect 4358 38533 4414 38589
rect 4440 38533 4496 38589
rect 4522 38533 4578 38589
rect 4604 38533 4660 38589
rect 4686 38567 4712 38589
rect 4712 38567 4742 38589
rect 4768 38567 4780 38589
rect 4780 38567 4824 38589
rect 4850 38617 4900 38619
rect 4900 38617 4906 38619
rect 4932 38617 4988 38673
rect 5195 38617 5251 38673
rect 5276 38617 5332 38673
rect 5357 38617 5413 38673
rect 5438 38617 5494 38673
rect 5519 38617 5575 38673
rect 5600 38632 5632 38673
rect 5632 38632 5656 38673
rect 5681 38632 5684 38673
rect 5684 38632 5700 38673
rect 5700 38632 5737 38673
rect 5762 38632 5768 38673
rect 5768 38632 5818 38673
rect 5600 38619 5656 38632
rect 5681 38619 5737 38632
rect 5762 38619 5818 38632
rect 5600 38617 5632 38619
rect 5632 38617 5656 38619
rect 5681 38617 5684 38619
rect 5684 38617 5700 38619
rect 5700 38617 5737 38619
rect 5762 38617 5768 38619
rect 5768 38617 5818 38619
rect 5843 38617 5899 38673
rect 5924 38617 5980 38673
rect 6005 38617 6061 38673
rect 6086 38617 6142 38673
rect 6167 38617 6223 38673
rect 6248 38617 6304 38673
rect 6329 38617 6385 38673
rect 6410 38617 6466 38673
rect 6491 38617 6547 38673
rect 6572 38632 6604 38673
rect 6604 38632 6620 38673
rect 6620 38632 6628 38673
rect 6653 38632 6672 38673
rect 6672 38632 6688 38673
rect 6688 38632 6709 38673
rect 6734 38632 6740 38673
rect 6740 38632 6790 38673
rect 6572 38619 6628 38632
rect 6653 38619 6709 38632
rect 6734 38619 6790 38632
rect 6572 38617 6604 38619
rect 6604 38617 6620 38619
rect 6620 38617 6628 38619
rect 6653 38617 6672 38619
rect 6672 38617 6688 38619
rect 6688 38617 6709 38619
rect 6734 38617 6740 38619
rect 6740 38617 6790 38619
rect 6815 38617 6871 38673
rect 6896 38617 6952 38673
rect 6977 38617 7033 38673
rect 7058 38617 7114 38673
rect 7139 38617 7195 38673
rect 7221 38617 7277 38673
rect 7303 38617 7359 38673
rect 4850 38567 4900 38589
rect 4900 38567 4906 38589
rect 4686 38554 4742 38567
rect 4768 38554 4824 38567
rect 4850 38554 4906 38567
rect 4686 38533 4712 38554
rect 4712 38533 4742 38554
rect 4768 38533 4780 38554
rect 4780 38533 4824 38554
rect 3862 38502 3912 38505
rect 3912 38502 3918 38505
rect 3945 38502 3980 38505
rect 3980 38502 4001 38505
rect 3779 38490 3835 38502
rect 3862 38490 3918 38502
rect 3945 38490 4001 38502
rect 3779 38449 3792 38490
rect 3792 38449 3835 38490
rect 3862 38449 3912 38490
rect 3912 38449 3918 38490
rect 3945 38449 3980 38490
rect 3980 38449 4001 38490
rect 4028 38449 4084 38505
rect 4111 38449 4167 38505
rect 4194 38449 4250 38505
rect 4276 38449 4332 38505
rect 4358 38449 4414 38505
rect 4440 38449 4496 38505
rect 4522 38449 4578 38505
rect 4604 38449 4660 38505
rect 4686 38502 4712 38505
rect 4712 38502 4742 38505
rect 4768 38502 4780 38505
rect 4780 38502 4824 38505
rect 4850 38533 4900 38554
rect 4900 38533 4906 38554
rect 4932 38533 4988 38589
rect 5195 38533 5251 38589
rect 5276 38533 5332 38589
rect 5357 38533 5413 38589
rect 5438 38533 5494 38589
rect 5519 38533 5575 38589
rect 5600 38567 5632 38589
rect 5632 38567 5656 38589
rect 5681 38567 5684 38589
rect 5684 38567 5700 38589
rect 5700 38567 5737 38589
rect 5762 38567 5768 38589
rect 5768 38567 5818 38589
rect 5600 38554 5656 38567
rect 5681 38554 5737 38567
rect 5762 38554 5818 38567
rect 5600 38533 5632 38554
rect 5632 38533 5656 38554
rect 5681 38533 5684 38554
rect 5684 38533 5700 38554
rect 5700 38533 5737 38554
rect 5762 38533 5768 38554
rect 5768 38533 5818 38554
rect 5843 38533 5899 38589
rect 5924 38533 5980 38589
rect 6005 38533 6061 38589
rect 6086 38533 6142 38589
rect 6167 38533 6223 38589
rect 6248 38533 6304 38589
rect 6329 38533 6385 38589
rect 6410 38533 6466 38589
rect 6491 38533 6547 38589
rect 6572 38567 6604 38589
rect 6604 38567 6620 38589
rect 6620 38567 6628 38589
rect 6653 38567 6672 38589
rect 6672 38567 6688 38589
rect 6688 38567 6709 38589
rect 6734 38567 6740 38589
rect 6740 38567 6790 38589
rect 6572 38554 6628 38567
rect 6653 38554 6709 38567
rect 6734 38554 6790 38567
rect 6572 38533 6604 38554
rect 6604 38533 6620 38554
rect 6620 38533 6628 38554
rect 6653 38533 6672 38554
rect 6672 38533 6688 38554
rect 6688 38533 6709 38554
rect 6734 38533 6740 38554
rect 6740 38533 6790 38554
rect 6815 38533 6871 38589
rect 6896 38533 6952 38589
rect 6977 38533 7033 38589
rect 7058 38533 7114 38589
rect 7139 38533 7195 38589
rect 7221 38533 7277 38589
rect 7303 38533 7359 38589
rect 4850 38502 4900 38505
rect 4900 38502 4906 38505
rect 4686 38490 4742 38502
rect 4768 38490 4824 38502
rect 4850 38490 4906 38502
rect 4686 38449 4712 38490
rect 4712 38449 4742 38490
rect 4768 38449 4780 38490
rect 4780 38449 4824 38490
rect 4850 38449 4900 38490
rect 4900 38449 4906 38490
rect 4932 38449 4988 38505
rect 5195 38449 5251 38505
rect 5276 38449 5332 38505
rect 5357 38449 5413 38505
rect 5438 38449 5494 38505
rect 5519 38449 5575 38505
rect 5600 38502 5632 38505
rect 5632 38502 5656 38505
rect 5681 38502 5684 38505
rect 5684 38502 5700 38505
rect 5700 38502 5737 38505
rect 5762 38502 5768 38505
rect 5768 38502 5818 38505
rect 5600 38490 5656 38502
rect 5681 38490 5737 38502
rect 5762 38490 5818 38502
rect 5600 38449 5632 38490
rect 5632 38449 5656 38490
rect 5681 38449 5684 38490
rect 5684 38449 5700 38490
rect 5700 38449 5737 38490
rect 5762 38449 5768 38490
rect 5768 38449 5818 38490
rect 5843 38449 5899 38505
rect 5924 38449 5980 38505
rect 6005 38449 6061 38505
rect 6086 38449 6142 38505
rect 6167 38449 6223 38505
rect 6248 38449 6304 38505
rect 6329 38449 6385 38505
rect 6410 38449 6466 38505
rect 6491 38449 6547 38505
rect 6572 38502 6604 38505
rect 6604 38502 6620 38505
rect 6620 38502 6628 38505
rect 6653 38502 6672 38505
rect 6672 38502 6688 38505
rect 6688 38502 6709 38505
rect 6734 38502 6740 38505
rect 6740 38502 6790 38505
rect 6572 38490 6628 38502
rect 6653 38490 6709 38502
rect 6734 38490 6790 38502
rect 6572 38449 6604 38490
rect 6604 38449 6620 38490
rect 6620 38449 6628 38490
rect 6653 38449 6672 38490
rect 6672 38449 6688 38490
rect 6688 38449 6709 38490
rect 6734 38449 6740 38490
rect 6740 38449 6790 38490
rect 6815 38449 6871 38505
rect 6896 38449 6952 38505
rect 6977 38449 7033 38505
rect 7058 38449 7114 38505
rect 7139 38449 7195 38505
rect 7221 38449 7277 38505
rect 7303 38449 7359 38505
rect 2534 38365 2590 38421
rect 2617 38365 2673 38421
rect 2700 38365 2756 38421
rect 2783 38365 2839 38421
rect 2866 38374 2872 38421
rect 2872 38374 2922 38421
rect 2949 38374 2992 38421
rect 2992 38374 3005 38421
rect 3032 38374 3060 38421
rect 3060 38374 3088 38421
rect 2866 38365 2922 38374
rect 2949 38365 3005 38374
rect 3032 38365 3088 38374
rect 3115 38365 3171 38421
rect 3198 38365 3254 38421
rect 3281 38365 3337 38421
rect 3364 38365 3420 38421
rect 3447 38365 3503 38421
rect 3530 38365 3586 38421
rect 3613 38365 3669 38421
rect 3696 38365 3752 38421
rect 3779 38374 3792 38421
rect 3792 38374 3835 38421
rect 3862 38374 3912 38421
rect 3912 38374 3918 38421
rect 3945 38374 3980 38421
rect 3980 38374 4001 38421
rect 3779 38365 3835 38374
rect 3862 38365 3918 38374
rect 3945 38365 4001 38374
rect 4028 38365 4084 38421
rect 4111 38365 4167 38421
rect 4194 38365 4250 38421
rect 4276 38365 4332 38421
rect 4358 38365 4414 38421
rect 4440 38365 4496 38421
rect 4522 38365 4578 38421
rect 4604 38365 4660 38421
rect 4686 38374 4712 38421
rect 4712 38374 4742 38421
rect 4768 38374 4780 38421
rect 4780 38374 4824 38421
rect 4850 38374 4900 38421
rect 4900 38374 4906 38421
rect 4686 38365 4742 38374
rect 4768 38365 4824 38374
rect 4850 38365 4906 38374
rect 4932 38365 4988 38421
rect 5195 38365 5251 38421
rect 5276 38365 5332 38421
rect 5357 38365 5413 38421
rect 5438 38365 5494 38421
rect 5519 38365 5575 38421
rect 5600 38374 5632 38421
rect 5632 38374 5656 38421
rect 5681 38374 5684 38421
rect 5684 38374 5700 38421
rect 5700 38374 5737 38421
rect 5762 38374 5768 38421
rect 5768 38374 5818 38421
rect 5600 38365 5656 38374
rect 5681 38365 5737 38374
rect 5762 38365 5818 38374
rect 5843 38365 5899 38421
rect 5924 38365 5980 38421
rect 6005 38365 6061 38421
rect 6086 38365 6142 38421
rect 6167 38365 6223 38421
rect 6248 38365 6304 38421
rect 6329 38365 6385 38421
rect 6410 38365 6466 38421
rect 6491 38365 6547 38421
rect 6572 38374 6604 38421
rect 6604 38374 6620 38421
rect 6620 38374 6628 38421
rect 6653 38374 6672 38421
rect 6672 38374 6688 38421
rect 6688 38374 6709 38421
rect 6734 38374 6740 38421
rect 6740 38374 6790 38421
rect 6572 38365 6628 38374
rect 6653 38365 6709 38374
rect 6734 38365 6790 38374
rect 6815 38365 6871 38421
rect 6896 38365 6952 38421
rect 6977 38365 7033 38421
rect 7058 38365 7114 38421
rect 7139 38365 7195 38421
rect 7221 38365 7277 38421
rect 7303 38365 7359 38421
rect 2534 38281 2590 38337
rect 2617 38281 2673 38337
rect 2700 38281 2756 38337
rect 2783 38281 2839 38337
rect 2866 38310 2872 38337
rect 2872 38310 2922 38337
rect 2949 38310 2992 38337
rect 2992 38310 3005 38337
rect 3032 38310 3060 38337
rect 3060 38310 3088 38337
rect 2866 38298 2922 38310
rect 2949 38298 3005 38310
rect 3032 38298 3088 38310
rect 2866 38281 2872 38298
rect 2872 38281 2922 38298
rect 2534 38197 2590 38253
rect 2617 38197 2673 38253
rect 2700 38197 2756 38253
rect 2783 38197 2839 38253
rect 2866 38246 2872 38253
rect 2872 38246 2922 38253
rect 2949 38281 2992 38298
rect 2992 38281 3005 38298
rect 3032 38281 3060 38298
rect 3060 38281 3088 38298
rect 3115 38281 3171 38337
rect 3198 38281 3254 38337
rect 3281 38281 3337 38337
rect 3364 38281 3420 38337
rect 3447 38281 3503 38337
rect 3530 38281 3586 38337
rect 3613 38281 3669 38337
rect 3696 38281 3752 38337
rect 3779 38310 3792 38337
rect 3792 38310 3835 38337
rect 3862 38310 3912 38337
rect 3912 38310 3918 38337
rect 3945 38310 3980 38337
rect 3980 38310 4001 38337
rect 3779 38298 3835 38310
rect 3862 38298 3918 38310
rect 3945 38298 4001 38310
rect 3779 38281 3792 38298
rect 3792 38281 3835 38298
rect 2949 38246 2992 38253
rect 2992 38246 3005 38253
rect 3032 38246 3060 38253
rect 3060 38246 3088 38253
rect 2866 38234 2922 38246
rect 2949 38234 3005 38246
rect 3032 38234 3088 38246
rect 2866 38197 2872 38234
rect 2872 38197 2922 38234
rect 2949 38197 2992 38234
rect 2992 38197 3005 38234
rect 3032 38197 3060 38234
rect 3060 38197 3088 38234
rect 3115 38197 3171 38253
rect 3198 38197 3254 38253
rect 3281 38197 3337 38253
rect 3364 38197 3420 38253
rect 3447 38197 3503 38253
rect 3530 38197 3586 38253
rect 3613 38197 3669 38253
rect 3696 38197 3752 38253
rect 3779 38246 3792 38253
rect 3792 38246 3835 38253
rect 3862 38281 3912 38298
rect 3912 38281 3918 38298
rect 3945 38281 3980 38298
rect 3980 38281 4001 38298
rect 4028 38281 4084 38337
rect 4111 38281 4167 38337
rect 4194 38281 4250 38337
rect 4276 38281 4332 38337
rect 4358 38281 4414 38337
rect 4440 38281 4496 38337
rect 4522 38281 4578 38337
rect 4604 38281 4660 38337
rect 4686 38310 4712 38337
rect 4712 38310 4742 38337
rect 4768 38310 4780 38337
rect 4780 38310 4824 38337
rect 4850 38310 4900 38337
rect 4900 38310 4906 38337
rect 4686 38298 4742 38310
rect 4768 38298 4824 38310
rect 4850 38298 4906 38310
rect 4686 38281 4712 38298
rect 4712 38281 4742 38298
rect 4768 38281 4780 38298
rect 4780 38281 4824 38298
rect 3862 38246 3912 38253
rect 3912 38246 3918 38253
rect 3945 38246 3980 38253
rect 3980 38246 4001 38253
rect 3779 38234 3835 38246
rect 3862 38234 3918 38246
rect 3945 38234 4001 38246
rect 3779 38197 3792 38234
rect 3792 38197 3835 38234
rect 3862 38197 3912 38234
rect 3912 38197 3918 38234
rect 3945 38197 3980 38234
rect 3980 38197 4001 38234
rect 4028 38197 4084 38253
rect 4111 38197 4167 38253
rect 4194 38197 4250 38253
rect 4276 38197 4332 38253
rect 4358 38197 4414 38253
rect 4440 38197 4496 38253
rect 4522 38197 4578 38253
rect 4604 38197 4660 38253
rect 4686 38246 4712 38253
rect 4712 38246 4742 38253
rect 4768 38246 4780 38253
rect 4780 38246 4824 38253
rect 4850 38281 4900 38298
rect 4900 38281 4906 38298
rect 4932 38281 4988 38337
rect 5195 38281 5251 38337
rect 5276 38281 5332 38337
rect 5357 38281 5413 38337
rect 5438 38281 5494 38337
rect 5519 38281 5575 38337
rect 5600 38310 5632 38337
rect 5632 38310 5656 38337
rect 5681 38310 5684 38337
rect 5684 38310 5700 38337
rect 5700 38310 5737 38337
rect 5762 38310 5768 38337
rect 5768 38310 5818 38337
rect 5600 38298 5656 38310
rect 5681 38298 5737 38310
rect 5762 38298 5818 38310
rect 5600 38281 5632 38298
rect 5632 38281 5656 38298
rect 5681 38281 5684 38298
rect 5684 38281 5700 38298
rect 5700 38281 5737 38298
rect 5762 38281 5768 38298
rect 5768 38281 5818 38298
rect 5843 38281 5899 38337
rect 5924 38281 5980 38337
rect 6005 38281 6061 38337
rect 6086 38281 6142 38337
rect 6167 38281 6223 38337
rect 6248 38281 6304 38337
rect 6329 38281 6385 38337
rect 6410 38281 6466 38337
rect 6491 38281 6547 38337
rect 6572 38310 6604 38337
rect 6604 38310 6620 38337
rect 6620 38310 6628 38337
rect 6653 38310 6672 38337
rect 6672 38310 6688 38337
rect 6688 38310 6709 38337
rect 6734 38310 6740 38337
rect 6740 38310 6790 38337
rect 6572 38298 6628 38310
rect 6653 38298 6709 38310
rect 6734 38298 6790 38310
rect 6572 38281 6604 38298
rect 6604 38281 6620 38298
rect 6620 38281 6628 38298
rect 6653 38281 6672 38298
rect 6672 38281 6688 38298
rect 6688 38281 6709 38298
rect 6734 38281 6740 38298
rect 6740 38281 6790 38298
rect 6815 38281 6871 38337
rect 6896 38281 6952 38337
rect 6977 38281 7033 38337
rect 7058 38281 7114 38337
rect 7139 38281 7195 38337
rect 7221 38281 7277 38337
rect 7303 38281 7359 38337
rect 4850 38246 4900 38253
rect 4900 38246 4906 38253
rect 4686 38234 4742 38246
rect 4768 38234 4824 38246
rect 4850 38234 4906 38246
rect 4686 38197 4712 38234
rect 4712 38197 4742 38234
rect 4768 38197 4780 38234
rect 4780 38197 4824 38234
rect 4850 38197 4900 38234
rect 4900 38197 4906 38234
rect 4932 38197 4988 38253
rect 5195 38197 5251 38253
rect 5276 38197 5332 38253
rect 5357 38197 5413 38253
rect 5438 38197 5494 38253
rect 5519 38197 5575 38253
rect 5600 38246 5632 38253
rect 5632 38246 5656 38253
rect 5681 38246 5684 38253
rect 5684 38246 5700 38253
rect 5700 38246 5737 38253
rect 5762 38246 5768 38253
rect 5768 38246 5818 38253
rect 5600 38234 5656 38246
rect 5681 38234 5737 38246
rect 5762 38234 5818 38246
rect 5600 38197 5632 38234
rect 5632 38197 5656 38234
rect 5681 38197 5684 38234
rect 5684 38197 5700 38234
rect 5700 38197 5737 38234
rect 5762 38197 5768 38234
rect 5768 38197 5818 38234
rect 5843 38197 5899 38253
rect 5924 38197 5980 38253
rect 6005 38197 6061 38253
rect 6086 38197 6142 38253
rect 6167 38197 6223 38253
rect 6248 38197 6304 38253
rect 6329 38197 6385 38253
rect 6410 38197 6466 38253
rect 6491 38197 6547 38253
rect 6572 38246 6604 38253
rect 6604 38246 6620 38253
rect 6620 38246 6628 38253
rect 6653 38246 6672 38253
rect 6672 38246 6688 38253
rect 6688 38246 6709 38253
rect 6734 38246 6740 38253
rect 6740 38246 6790 38253
rect 6572 38234 6628 38246
rect 6653 38234 6709 38246
rect 6734 38234 6790 38246
rect 6572 38197 6604 38234
rect 6604 38197 6620 38234
rect 6620 38197 6628 38234
rect 6653 38197 6672 38234
rect 6672 38197 6688 38234
rect 6688 38197 6709 38234
rect 6734 38197 6740 38234
rect 6740 38197 6790 38234
rect 6815 38197 6871 38253
rect 6896 38197 6952 38253
rect 6977 38197 7033 38253
rect 7058 38197 7114 38253
rect 7139 38197 7195 38253
rect 7221 38197 7277 38253
rect 7303 38197 7359 38253
rect 2534 38113 2590 38169
rect 2617 38113 2673 38169
rect 2700 38113 2756 38169
rect 2783 38113 2839 38169
rect 2866 38118 2872 38169
rect 2872 38118 2922 38169
rect 2949 38118 2992 38169
rect 2992 38118 3005 38169
rect 3032 38118 3060 38169
rect 3060 38118 3088 38169
rect 2866 38113 2922 38118
rect 2949 38113 3005 38118
rect 3032 38113 3088 38118
rect 3115 38113 3171 38169
rect 3198 38113 3254 38169
rect 3281 38113 3337 38169
rect 3364 38113 3420 38169
rect 3447 38113 3503 38169
rect 3530 38113 3586 38169
rect 3613 38113 3669 38169
rect 3696 38113 3752 38169
rect 3779 38118 3792 38169
rect 3792 38118 3835 38169
rect 3862 38118 3912 38169
rect 3912 38118 3918 38169
rect 3945 38118 3980 38169
rect 3980 38118 4001 38169
rect 3779 38113 3835 38118
rect 3862 38113 3918 38118
rect 3945 38113 4001 38118
rect 4028 38113 4084 38169
rect 4111 38113 4167 38169
rect 4194 38113 4250 38169
rect 4276 38113 4332 38169
rect 4358 38113 4414 38169
rect 4440 38113 4496 38169
rect 4522 38113 4578 38169
rect 4604 38113 4660 38169
rect 4686 38118 4712 38169
rect 4712 38118 4742 38169
rect 4768 38118 4780 38169
rect 4780 38118 4824 38169
rect 4850 38118 4900 38169
rect 4900 38118 4906 38169
rect 4686 38113 4742 38118
rect 4768 38113 4824 38118
rect 4850 38113 4906 38118
rect 4932 38113 4988 38169
rect 5195 38113 5251 38169
rect 5276 38113 5332 38169
rect 5357 38113 5413 38169
rect 5438 38113 5494 38169
rect 5519 38113 5575 38169
rect 5600 38118 5632 38169
rect 5632 38118 5656 38169
rect 5681 38118 5684 38169
rect 5684 38118 5700 38169
rect 5700 38118 5737 38169
rect 5762 38118 5768 38169
rect 5768 38118 5818 38169
rect 5600 38113 5656 38118
rect 5681 38113 5737 38118
rect 5762 38113 5818 38118
rect 5843 38113 5899 38169
rect 5924 38113 5980 38169
rect 6005 38113 6061 38169
rect 6086 38113 6142 38169
rect 6167 38113 6223 38169
rect 6248 38113 6304 38169
rect 6329 38113 6385 38169
rect 6410 38113 6466 38169
rect 6491 38113 6547 38169
rect 6572 38118 6604 38169
rect 6604 38118 6620 38169
rect 6620 38118 6628 38169
rect 6653 38118 6672 38169
rect 6672 38118 6688 38169
rect 6688 38118 6709 38169
rect 6734 38118 6740 38169
rect 6740 38118 6790 38169
rect 6572 38113 6628 38118
rect 6653 38113 6709 38118
rect 6734 38113 6790 38118
rect 6815 38113 6871 38169
rect 6896 38113 6952 38169
rect 6977 38113 7033 38169
rect 7058 38113 7114 38169
rect 7139 38113 7195 38169
rect 7221 38113 7277 38169
rect 7303 38113 7359 38169
rect 2531 38017 2587 38073
rect 2649 38017 2705 38073
rect 2767 38017 2823 38073
rect 2531 37932 2587 37988
rect 2649 37932 2705 37988
rect 2767 37932 2823 37988
rect 2531 37847 2587 37903
rect 2649 37847 2705 37903
rect 2767 37847 2823 37903
rect 2531 37762 2587 37818
rect 2649 37762 2705 37818
rect 2767 37762 2823 37818
rect 2531 37677 2587 37733
rect 2649 37677 2705 37733
rect 2767 37677 2823 37733
rect 2531 37592 2587 37648
rect 2649 37592 2705 37648
rect 2767 37592 2823 37648
rect 2531 37507 2587 37563
rect 2649 37507 2705 37563
rect 2767 37507 2823 37563
rect 2531 37422 2587 37478
rect 2649 37422 2705 37478
rect 2767 37422 2823 37478
rect 2531 37337 2587 37393
rect 2649 37337 2705 37393
rect 2767 37337 2823 37393
rect 2531 37252 2587 37308
rect 2649 37252 2705 37308
rect 2767 37252 2823 37308
rect 2531 37166 2587 37222
rect 2649 37166 2705 37222
rect 2767 37166 2823 37222
rect 2531 37080 2587 37136
rect 2649 37080 2705 37136
rect 2767 37080 2823 37136
rect 2531 36994 2587 37050
rect 2649 36994 2705 37050
rect 2767 36994 2823 37050
rect 2531 36908 2587 36964
rect 2649 36908 2705 36964
rect 2767 36908 2823 36964
rect 2531 36822 2587 36878
rect 2649 36822 2705 36878
rect 2767 36822 2823 36878
rect 2538 36716 2594 36772
rect 2632 36716 2688 36772
rect 2726 36716 2782 36772
rect 2820 36716 2876 36772
rect 2914 36716 2970 36772
rect 3008 36716 3064 36772
rect 2538 36636 2594 36692
rect 2632 36636 2688 36692
rect 2726 36636 2782 36692
rect 2820 36636 2876 36692
rect 2914 36636 2970 36692
rect 3008 36636 3064 36692
rect 2538 36556 2594 36612
rect 2632 36556 2688 36612
rect 2726 36556 2782 36612
rect 2820 36556 2876 36612
rect 2914 36556 2970 36612
rect 3008 36556 3064 36612
rect 3099 36594 3155 36650
rect 2538 36476 2594 36532
rect 2632 36476 2688 36532
rect 2726 36476 2782 36532
rect 2820 36476 2876 36532
rect 2914 36476 2970 36532
rect 3008 36476 3064 36532
rect 3112 36506 3168 36562
rect 3206 36506 3262 36562
rect 2538 36396 2594 36452
rect 2632 36396 2688 36452
rect 2726 36396 2782 36452
rect 2820 36396 2876 36452
rect 2914 36396 2970 36452
rect 3008 36396 3064 36452
rect 3112 36420 3168 36476
rect 3206 36420 3262 36476
rect 2538 36316 2594 36372
rect 2632 36316 2688 36372
rect 2726 36316 2782 36372
rect 2820 36368 2876 36372
rect 2914 36368 2970 36372
rect 3008 36368 3064 36372
rect 2820 36316 2872 36368
rect 2872 36316 2876 36368
rect 2914 36316 2924 36368
rect 2924 36316 2940 36368
rect 2940 36316 2970 36368
rect 3008 36316 3060 36368
rect 3060 36316 3064 36368
rect 3112 36334 3168 36390
rect 3206 36334 3262 36390
rect 3321 36359 3377 36415
rect 2538 36236 2594 36292
rect 2632 36236 2688 36292
rect 2726 36236 2782 36292
rect 2820 36252 2872 36292
rect 2872 36252 2876 36292
rect 2914 36252 2924 36292
rect 2924 36252 2940 36292
rect 2940 36252 2970 36292
rect 3008 36252 3060 36292
rect 3060 36252 3064 36292
rect 2820 36239 2876 36252
rect 2914 36239 2970 36252
rect 3008 36239 3064 36252
rect 2820 36236 2872 36239
rect 2872 36236 2876 36239
rect 2914 36236 2924 36239
rect 2924 36236 2940 36239
rect 2940 36236 2970 36239
rect 2538 36156 2594 36212
rect 2632 36156 2688 36212
rect 2726 36156 2782 36212
rect 2820 36187 2872 36212
rect 2872 36187 2876 36212
rect 2914 36187 2924 36212
rect 2924 36187 2940 36212
rect 2940 36187 2970 36212
rect 3008 36236 3060 36239
rect 3060 36236 3064 36239
rect 3109 36238 3165 36294
rect 3193 36238 3249 36294
rect 3277 36238 3333 36294
rect 3360 36238 3416 36294
rect 3443 36238 3499 36294
rect 3526 36238 3582 36294
rect 3609 36238 3665 36294
rect 3692 36238 3748 36294
rect 3775 36290 3831 36294
rect 3858 36290 3914 36294
rect 3941 36290 3997 36294
rect 3775 36238 3792 36290
rect 3792 36238 3831 36290
rect 3858 36238 3860 36290
rect 3860 36238 3912 36290
rect 3912 36238 3914 36290
rect 3941 36238 3980 36290
rect 3980 36238 3997 36290
rect 4024 36238 4080 36294
rect 4107 36238 4163 36294
rect 4190 36238 4246 36294
rect 4273 36238 4329 36294
rect 4356 36238 4412 36294
rect 4439 36238 4495 36294
rect 4522 36238 4578 36294
rect 4605 36238 4661 36294
rect 4688 36290 4744 36294
rect 4771 36290 4827 36294
rect 4854 36290 4910 36294
rect 4688 36238 4712 36290
rect 4712 36238 4744 36290
rect 4771 36238 4780 36290
rect 4780 36238 4827 36290
rect 4854 36238 4900 36290
rect 4900 36238 4910 36290
rect 4937 36238 4993 36294
rect 5195 36238 5251 36294
rect 5277 36238 5333 36294
rect 5359 36238 5415 36294
rect 5441 36238 5497 36294
rect 5523 36238 5579 36294
rect 5605 36290 5661 36294
rect 5687 36290 5743 36294
rect 5769 36290 5825 36294
rect 5605 36238 5632 36290
rect 5632 36238 5661 36290
rect 5687 36238 5700 36290
rect 5700 36238 5743 36290
rect 5769 36238 5820 36290
rect 5820 36238 5825 36290
rect 5851 36238 5907 36294
rect 5933 36238 5989 36294
rect 6015 36238 6071 36294
rect 6097 36238 6153 36294
rect 6179 36238 6235 36294
rect 6261 36238 6317 36294
rect 6343 36238 6399 36294
rect 6425 36238 6481 36294
rect 6507 36290 6563 36294
rect 6589 36290 6645 36294
rect 6671 36290 6727 36294
rect 6507 36238 6552 36290
rect 6552 36238 6563 36290
rect 6589 36238 6604 36290
rect 6604 36238 6620 36290
rect 6620 36238 6645 36290
rect 6671 36238 6672 36290
rect 6672 36238 6688 36290
rect 6688 36238 6727 36290
rect 6753 36238 6809 36294
rect 3008 36187 3060 36212
rect 3060 36187 3064 36212
rect 2820 36174 2876 36187
rect 2914 36174 2970 36187
rect 3008 36174 3064 36187
rect 2820 36156 2872 36174
rect 2872 36156 2876 36174
rect 2914 36156 2924 36174
rect 2924 36156 2940 36174
rect 2940 36156 2970 36174
rect 2538 36076 2594 36132
rect 2632 36076 2688 36132
rect 2726 36076 2782 36132
rect 2820 36122 2872 36132
rect 2872 36122 2876 36132
rect 2914 36122 2924 36132
rect 2924 36122 2940 36132
rect 2940 36122 2970 36132
rect 3008 36156 3060 36174
rect 3060 36156 3064 36174
rect 3109 36158 3165 36214
rect 3193 36158 3249 36214
rect 3277 36158 3333 36214
rect 3360 36158 3416 36214
rect 3443 36158 3499 36214
rect 3526 36158 3582 36214
rect 3609 36158 3665 36214
rect 3692 36158 3748 36214
rect 3775 36174 3792 36214
rect 3792 36174 3831 36214
rect 3858 36174 3860 36214
rect 3860 36174 3912 36214
rect 3912 36174 3914 36214
rect 3941 36174 3980 36214
rect 3980 36174 3997 36214
rect 3775 36162 3831 36174
rect 3858 36162 3914 36174
rect 3941 36162 3997 36174
rect 3775 36158 3792 36162
rect 3792 36158 3831 36162
rect 3858 36158 3860 36162
rect 3860 36158 3912 36162
rect 3912 36158 3914 36162
rect 3941 36158 3980 36162
rect 3980 36158 3997 36162
rect 4024 36158 4080 36214
rect 4107 36158 4163 36214
rect 4190 36158 4246 36214
rect 4273 36158 4329 36214
rect 4356 36158 4412 36214
rect 4439 36158 4495 36214
rect 4522 36158 4578 36214
rect 4605 36158 4661 36214
rect 4688 36174 4712 36214
rect 4712 36174 4744 36214
rect 4771 36174 4780 36214
rect 4780 36174 4827 36214
rect 4854 36174 4900 36214
rect 4900 36174 4910 36214
rect 4688 36162 4744 36174
rect 4771 36162 4827 36174
rect 4854 36162 4910 36174
rect 4688 36158 4712 36162
rect 4712 36158 4744 36162
rect 4771 36158 4780 36162
rect 4780 36158 4827 36162
rect 3008 36122 3060 36132
rect 3060 36122 3064 36132
rect 2820 36109 2876 36122
rect 2914 36109 2970 36122
rect 3008 36109 3064 36122
rect 2820 36076 2872 36109
rect 2872 36076 2876 36109
rect 2914 36076 2924 36109
rect 2924 36076 2940 36109
rect 2940 36076 2970 36109
rect 3008 36076 3060 36109
rect 3060 36076 3064 36109
rect 3109 36078 3165 36134
rect 3193 36078 3249 36134
rect 3277 36078 3333 36134
rect 3360 36078 3416 36134
rect 3443 36078 3499 36134
rect 3526 36078 3582 36134
rect 3609 36078 3665 36134
rect 3692 36078 3748 36134
rect 3775 36110 3792 36134
rect 3792 36110 3831 36134
rect 3858 36110 3860 36134
rect 3860 36110 3912 36134
rect 3912 36110 3914 36134
rect 3941 36110 3980 36134
rect 3980 36110 3997 36134
rect 3775 36098 3831 36110
rect 3858 36098 3914 36110
rect 3941 36098 3997 36110
rect 3775 36078 3792 36098
rect 3792 36078 3831 36098
rect 3858 36078 3860 36098
rect 3860 36078 3912 36098
rect 3912 36078 3914 36098
rect 3941 36078 3980 36098
rect 3980 36078 3997 36098
rect 4024 36078 4080 36134
rect 4107 36078 4163 36134
rect 4190 36078 4246 36134
rect 4273 36078 4329 36134
rect 4356 36078 4412 36134
rect 4439 36078 4495 36134
rect 4522 36078 4578 36134
rect 4605 36078 4661 36134
rect 4688 36110 4712 36134
rect 4712 36110 4744 36134
rect 4771 36110 4780 36134
rect 4780 36110 4827 36134
rect 4854 36158 4900 36162
rect 4900 36158 4910 36162
rect 4937 36158 4993 36214
rect 5195 36158 5251 36214
rect 5277 36158 5333 36214
rect 5359 36158 5415 36214
rect 5441 36158 5497 36214
rect 5523 36158 5579 36214
rect 5605 36174 5632 36214
rect 5632 36174 5661 36214
rect 5687 36174 5700 36214
rect 5700 36174 5743 36214
rect 6853 36222 6909 36278
rect 6941 36222 6997 36278
rect 7029 36222 7085 36278
rect 7117 36222 7173 36278
rect 7205 36222 7261 36278
rect 7293 36222 7349 36278
rect 5769 36174 5820 36214
rect 5820 36174 5825 36214
rect 5605 36162 5661 36174
rect 5687 36162 5743 36174
rect 5769 36162 5825 36174
rect 5605 36158 5632 36162
rect 5632 36158 5661 36162
rect 5687 36158 5700 36162
rect 5700 36158 5743 36162
rect 4854 36110 4900 36134
rect 4900 36110 4910 36134
rect 4688 36098 4744 36110
rect 4771 36098 4827 36110
rect 4854 36098 4910 36110
rect 4688 36078 4712 36098
rect 4712 36078 4744 36098
rect 4771 36078 4780 36098
rect 4780 36078 4827 36098
rect 2538 35996 2594 36052
rect 2632 35996 2688 36052
rect 2726 35996 2782 36052
rect 2820 36044 2876 36052
rect 2914 36044 2970 36052
rect 3008 36044 3064 36052
rect 2820 35996 2872 36044
rect 2872 35996 2876 36044
rect 2914 35996 2924 36044
rect 2924 35996 2940 36044
rect 2940 35996 2970 36044
rect 3008 35996 3060 36044
rect 3060 35996 3064 36044
rect 3109 35998 3165 36054
rect 3193 35998 3249 36054
rect 3277 35998 3333 36054
rect 3360 35998 3416 36054
rect 3443 35998 3499 36054
rect 3526 35998 3582 36054
rect 3609 35998 3665 36054
rect 3692 35998 3748 36054
rect 3775 36046 3792 36054
rect 3792 36046 3831 36054
rect 3858 36046 3860 36054
rect 3860 36046 3912 36054
rect 3912 36046 3914 36054
rect 3941 36046 3980 36054
rect 3980 36046 3997 36054
rect 3775 36034 3831 36046
rect 3858 36034 3914 36046
rect 3941 36034 3997 36046
rect 3775 35998 3792 36034
rect 3792 35998 3831 36034
rect 3858 35998 3860 36034
rect 3860 35998 3912 36034
rect 3912 35998 3914 36034
rect 3941 35998 3980 36034
rect 3980 35998 3997 36034
rect 4024 35998 4080 36054
rect 4107 35998 4163 36054
rect 4190 35998 4246 36054
rect 4273 35998 4329 36054
rect 4356 35998 4412 36054
rect 4439 35998 4495 36054
rect 4522 35998 4578 36054
rect 4605 35998 4661 36054
rect 4688 36046 4712 36054
rect 4712 36046 4744 36054
rect 4771 36046 4780 36054
rect 4780 36046 4827 36054
rect 4854 36078 4900 36098
rect 4900 36078 4910 36098
rect 4937 36078 4993 36134
rect 5195 36078 5251 36134
rect 5277 36078 5333 36134
rect 5359 36078 5415 36134
rect 5441 36078 5497 36134
rect 5523 36078 5579 36134
rect 5605 36110 5632 36134
rect 5632 36110 5661 36134
rect 5687 36110 5700 36134
rect 5700 36110 5743 36134
rect 5769 36158 5820 36162
rect 5820 36158 5825 36162
rect 5851 36158 5907 36214
rect 5933 36158 5989 36214
rect 6015 36158 6071 36214
rect 6097 36158 6153 36214
rect 6179 36158 6235 36214
rect 6261 36158 6317 36214
rect 6343 36158 6399 36214
rect 6425 36158 6481 36214
rect 6507 36174 6552 36214
rect 6552 36174 6563 36214
rect 6589 36174 6604 36214
rect 6604 36174 6620 36214
rect 6620 36174 6645 36214
rect 6671 36174 6672 36214
rect 6672 36174 6688 36214
rect 6688 36174 6727 36214
rect 6507 36162 6563 36174
rect 6589 36162 6645 36174
rect 6671 36162 6727 36174
rect 6507 36158 6552 36162
rect 6552 36158 6563 36162
rect 6589 36158 6604 36162
rect 6604 36158 6620 36162
rect 6620 36158 6645 36162
rect 6671 36158 6672 36162
rect 6672 36158 6688 36162
rect 6688 36158 6727 36162
rect 6753 36158 6809 36214
rect 6853 36140 6909 36196
rect 6941 36140 6997 36196
rect 7029 36140 7085 36196
rect 7117 36140 7173 36196
rect 7205 36140 7261 36196
rect 7293 36140 7349 36196
rect 5769 36110 5820 36134
rect 5820 36110 5825 36134
rect 5605 36098 5661 36110
rect 5687 36098 5743 36110
rect 5769 36098 5825 36110
rect 5605 36078 5632 36098
rect 5632 36078 5661 36098
rect 5687 36078 5700 36098
rect 5700 36078 5743 36098
rect 4854 36046 4900 36054
rect 4900 36046 4910 36054
rect 4688 36034 4744 36046
rect 4771 36034 4827 36046
rect 4854 36034 4910 36046
rect 4688 35998 4712 36034
rect 4712 35998 4744 36034
rect 4771 35998 4780 36034
rect 4780 35998 4827 36034
rect 4854 35998 4900 36034
rect 4900 35998 4910 36034
rect 4937 35998 4993 36054
rect 5195 35998 5251 36054
rect 5277 35998 5333 36054
rect 5359 35998 5415 36054
rect 5441 35998 5497 36054
rect 5523 35998 5579 36054
rect 5605 36046 5632 36054
rect 5632 36046 5661 36054
rect 5687 36046 5700 36054
rect 5700 36046 5743 36054
rect 5769 36078 5820 36098
rect 5820 36078 5825 36098
rect 5851 36078 5907 36134
rect 5933 36078 5989 36134
rect 6015 36078 6071 36134
rect 6097 36078 6153 36134
rect 6179 36078 6235 36134
rect 6261 36078 6317 36134
rect 6343 36078 6399 36134
rect 6425 36078 6481 36134
rect 6507 36110 6552 36134
rect 6552 36110 6563 36134
rect 6589 36110 6604 36134
rect 6604 36110 6620 36134
rect 6620 36110 6645 36134
rect 6671 36110 6672 36134
rect 6672 36110 6688 36134
rect 6688 36110 6727 36134
rect 6507 36098 6563 36110
rect 6589 36098 6645 36110
rect 6671 36098 6727 36110
rect 6507 36078 6552 36098
rect 6552 36078 6563 36098
rect 6589 36078 6604 36098
rect 6604 36078 6620 36098
rect 6620 36078 6645 36098
rect 6671 36078 6672 36098
rect 6672 36078 6688 36098
rect 6688 36078 6727 36098
rect 6753 36078 6809 36134
rect 6853 36058 6909 36114
rect 6941 36058 6997 36114
rect 7029 36058 7085 36114
rect 7117 36058 7173 36114
rect 7205 36058 7261 36114
rect 7293 36058 7349 36114
rect 5769 36046 5820 36054
rect 5820 36046 5825 36054
rect 5605 36034 5661 36046
rect 5687 36034 5743 36046
rect 5769 36034 5825 36046
rect 5605 35998 5632 36034
rect 5632 35998 5661 36034
rect 5687 35998 5700 36034
rect 5700 35998 5743 36034
rect 5769 35998 5820 36034
rect 5820 35998 5825 36034
rect 5851 35998 5907 36054
rect 5933 35998 5989 36054
rect 6015 35998 6071 36054
rect 6097 35998 6153 36054
rect 6179 35998 6235 36054
rect 6261 35998 6317 36054
rect 6343 35998 6399 36054
rect 6425 35998 6481 36054
rect 6507 36046 6552 36054
rect 6552 36046 6563 36054
rect 6589 36046 6604 36054
rect 6604 36046 6620 36054
rect 6620 36046 6645 36054
rect 6671 36046 6672 36054
rect 6672 36046 6688 36054
rect 6688 36046 6727 36054
rect 6507 36034 6563 36046
rect 6589 36034 6645 36046
rect 6671 36034 6727 36046
rect 6507 35998 6552 36034
rect 6552 35998 6563 36034
rect 6589 35998 6604 36034
rect 6604 35998 6620 36034
rect 6620 35998 6645 36034
rect 6671 35998 6672 36034
rect 6672 35998 6688 36034
rect 6688 35998 6727 36034
rect 6753 35998 6809 36054
rect 2538 35916 2594 35972
rect 2632 35916 2688 35972
rect 2726 35916 2782 35972
rect 2820 35927 2872 35972
rect 2872 35927 2876 35972
rect 2914 35927 2924 35972
rect 2924 35927 2940 35972
rect 2940 35927 2970 35972
rect 6853 35976 6909 36032
rect 6941 35976 6997 36032
rect 7029 35976 7085 36032
rect 7117 35976 7173 36032
rect 7205 35976 7261 36032
rect 7293 35976 7349 36032
rect 3008 35927 3060 35972
rect 3060 35927 3064 35972
rect 2820 35916 2876 35927
rect 2914 35916 2970 35927
rect 3008 35916 3064 35927
rect 3109 35918 3165 35974
rect 3193 35918 3249 35974
rect 3277 35918 3333 35974
rect 3360 35918 3416 35974
rect 3443 35918 3499 35974
rect 3526 35918 3582 35974
rect 3609 35918 3665 35974
rect 3692 35918 3748 35974
rect 3775 35970 3831 35974
rect 3858 35970 3914 35974
rect 3941 35970 3997 35974
rect 3775 35918 3792 35970
rect 3792 35918 3831 35970
rect 3858 35918 3860 35970
rect 3860 35918 3912 35970
rect 3912 35918 3914 35970
rect 3941 35918 3980 35970
rect 3980 35918 3997 35970
rect 4024 35918 4080 35974
rect 4107 35918 4163 35974
rect 4190 35918 4246 35974
rect 4273 35918 4329 35974
rect 4356 35918 4412 35974
rect 4439 35918 4495 35974
rect 4522 35918 4578 35974
rect 4605 35918 4661 35974
rect 4688 35970 4744 35974
rect 4771 35970 4827 35974
rect 4854 35970 4910 35974
rect 4688 35918 4712 35970
rect 4712 35918 4744 35970
rect 4771 35918 4780 35970
rect 4780 35918 4827 35970
rect 4854 35918 4900 35970
rect 4900 35918 4910 35970
rect 4937 35918 4993 35974
rect 5195 35918 5251 35974
rect 5277 35918 5333 35974
rect 5359 35918 5415 35974
rect 5441 35918 5497 35974
rect 5523 35918 5579 35974
rect 5605 35970 5661 35974
rect 5687 35970 5743 35974
rect 5769 35970 5825 35974
rect 5605 35918 5632 35970
rect 5632 35918 5661 35970
rect 5687 35918 5700 35970
rect 5700 35918 5743 35970
rect 5769 35918 5820 35970
rect 5820 35918 5825 35970
rect 5851 35918 5907 35974
rect 5933 35918 5989 35974
rect 6015 35918 6071 35974
rect 6097 35918 6153 35974
rect 6179 35918 6235 35974
rect 6261 35918 6317 35974
rect 6343 35918 6399 35974
rect 6425 35918 6481 35974
rect 6507 35970 6563 35974
rect 6589 35970 6645 35974
rect 6671 35970 6727 35974
rect 6507 35918 6552 35970
rect 6552 35918 6563 35970
rect 6589 35918 6604 35970
rect 6604 35918 6620 35970
rect 6620 35918 6645 35970
rect 6671 35918 6672 35970
rect 6672 35918 6688 35970
rect 6688 35918 6727 35970
rect 6753 35918 6809 35974
rect 2538 35836 2594 35892
rect 2632 35836 2688 35892
rect 2726 35836 2782 35892
rect 2820 35862 2872 35892
rect 2872 35862 2876 35892
rect 2914 35862 2924 35892
rect 2924 35862 2940 35892
rect 2940 35862 2970 35892
rect 3008 35862 3060 35892
rect 3060 35862 3064 35892
rect 2820 35849 2876 35862
rect 2914 35849 2970 35862
rect 3008 35849 3064 35862
rect 2820 35836 2872 35849
rect 2872 35836 2876 35849
rect 2914 35836 2924 35849
rect 2924 35836 2940 35849
rect 2940 35836 2970 35849
rect 2538 35756 2594 35812
rect 2632 35756 2688 35812
rect 2726 35756 2782 35812
rect 2820 35797 2872 35812
rect 2872 35797 2876 35812
rect 2914 35797 2924 35812
rect 2924 35797 2940 35812
rect 2940 35797 2970 35812
rect 3008 35836 3060 35849
rect 3060 35836 3064 35849
rect 3109 35838 3165 35894
rect 3193 35838 3249 35894
rect 3277 35838 3333 35894
rect 3360 35838 3416 35894
rect 3443 35838 3499 35894
rect 3526 35838 3582 35894
rect 3609 35838 3665 35894
rect 3692 35838 3748 35894
rect 3775 35854 3792 35894
rect 3792 35854 3831 35894
rect 3858 35854 3860 35894
rect 3860 35854 3912 35894
rect 3912 35854 3914 35894
rect 3941 35854 3980 35894
rect 3980 35854 3997 35894
rect 3775 35842 3831 35854
rect 3858 35842 3914 35854
rect 3941 35842 3997 35854
rect 3775 35838 3792 35842
rect 3792 35838 3831 35842
rect 3858 35838 3860 35842
rect 3860 35838 3912 35842
rect 3912 35838 3914 35842
rect 3941 35838 3980 35842
rect 3980 35838 3997 35842
rect 4024 35838 4080 35894
rect 4107 35838 4163 35894
rect 4190 35838 4246 35894
rect 4273 35838 4329 35894
rect 4356 35838 4412 35894
rect 4439 35838 4495 35894
rect 4522 35838 4578 35894
rect 4605 35838 4661 35894
rect 4688 35854 4712 35894
rect 4712 35854 4744 35894
rect 4771 35854 4780 35894
rect 4780 35854 4827 35894
rect 4854 35854 4900 35894
rect 4900 35854 4910 35894
rect 4688 35842 4744 35854
rect 4771 35842 4827 35854
rect 4854 35842 4910 35854
rect 4688 35838 4712 35842
rect 4712 35838 4744 35842
rect 4771 35838 4780 35842
rect 4780 35838 4827 35842
rect 3008 35797 3060 35812
rect 3060 35797 3064 35812
rect 2820 35784 2876 35797
rect 2914 35784 2970 35797
rect 3008 35784 3064 35797
rect 2820 35756 2872 35784
rect 2872 35756 2876 35784
rect 2914 35756 2924 35784
rect 2924 35756 2940 35784
rect 2940 35756 2970 35784
rect 3008 35756 3060 35784
rect 3060 35756 3064 35784
rect 3109 35758 3165 35814
rect 3193 35758 3249 35814
rect 3277 35758 3333 35814
rect 3360 35758 3416 35814
rect 3443 35758 3499 35814
rect 3526 35758 3582 35814
rect 3609 35758 3665 35814
rect 3692 35758 3748 35814
rect 3775 35790 3792 35814
rect 3792 35790 3831 35814
rect 3858 35790 3860 35814
rect 3860 35790 3912 35814
rect 3912 35790 3914 35814
rect 3941 35790 3980 35814
rect 3980 35790 3997 35814
rect 3775 35778 3831 35790
rect 3858 35778 3914 35790
rect 3941 35778 3997 35790
rect 3775 35758 3792 35778
rect 3792 35758 3831 35778
rect 3858 35758 3860 35778
rect 3860 35758 3912 35778
rect 3912 35758 3914 35778
rect 3941 35758 3980 35778
rect 3980 35758 3997 35778
rect 4024 35758 4080 35814
rect 4107 35758 4163 35814
rect 4190 35758 4246 35814
rect 4273 35758 4329 35814
rect 4356 35758 4412 35814
rect 4439 35758 4495 35814
rect 4522 35758 4578 35814
rect 4605 35758 4661 35814
rect 4688 35790 4712 35814
rect 4712 35790 4744 35814
rect 4771 35790 4780 35814
rect 4780 35790 4827 35814
rect 4854 35838 4900 35842
rect 4900 35838 4910 35842
rect 4937 35838 4993 35894
rect 5195 35838 5251 35894
rect 5277 35838 5333 35894
rect 5359 35838 5415 35894
rect 5441 35838 5497 35894
rect 5523 35838 5579 35894
rect 5605 35854 5632 35894
rect 5632 35854 5661 35894
rect 5687 35854 5700 35894
rect 5700 35854 5743 35894
rect 6853 35894 6909 35950
rect 6941 35894 6997 35950
rect 7029 35894 7085 35950
rect 7117 35894 7173 35950
rect 7205 35894 7261 35950
rect 7293 35894 7349 35950
rect 5769 35854 5820 35894
rect 5820 35854 5825 35894
rect 5605 35842 5661 35854
rect 5687 35842 5743 35854
rect 5769 35842 5825 35854
rect 5605 35838 5632 35842
rect 5632 35838 5661 35842
rect 5687 35838 5700 35842
rect 5700 35838 5743 35842
rect 4854 35790 4900 35814
rect 4900 35790 4910 35814
rect 4688 35778 4744 35790
rect 4771 35778 4827 35790
rect 4854 35778 4910 35790
rect 4688 35758 4712 35778
rect 4712 35758 4744 35778
rect 4771 35758 4780 35778
rect 4780 35758 4827 35778
rect 2538 35676 2594 35732
rect 2632 35676 2688 35732
rect 2726 35676 2782 35732
rect 2820 35719 2876 35732
rect 2914 35719 2970 35732
rect 3008 35719 3064 35732
rect 2820 35676 2872 35719
rect 2872 35676 2876 35719
rect 2914 35676 2924 35719
rect 2924 35676 2940 35719
rect 2940 35676 2970 35719
rect 3008 35676 3060 35719
rect 3060 35676 3064 35719
rect 3109 35678 3165 35734
rect 3193 35678 3249 35734
rect 3277 35678 3333 35734
rect 3360 35678 3416 35734
rect 3443 35678 3499 35734
rect 3526 35678 3582 35734
rect 3609 35678 3665 35734
rect 3692 35678 3748 35734
rect 3775 35726 3792 35734
rect 3792 35726 3831 35734
rect 3858 35726 3860 35734
rect 3860 35726 3912 35734
rect 3912 35726 3914 35734
rect 3941 35726 3980 35734
rect 3980 35726 3997 35734
rect 3775 35714 3831 35726
rect 3858 35714 3914 35726
rect 3941 35714 3997 35726
rect 3775 35678 3792 35714
rect 3792 35678 3831 35714
rect 3858 35678 3860 35714
rect 3860 35678 3912 35714
rect 3912 35678 3914 35714
rect 3941 35678 3980 35714
rect 3980 35678 3997 35714
rect 4024 35678 4080 35734
rect 4107 35678 4163 35734
rect 4190 35678 4246 35734
rect 4273 35678 4329 35734
rect 4356 35678 4412 35734
rect 4439 35678 4495 35734
rect 4522 35678 4578 35734
rect 4605 35678 4661 35734
rect 4688 35726 4712 35734
rect 4712 35726 4744 35734
rect 4771 35726 4780 35734
rect 4780 35726 4827 35734
rect 4854 35758 4900 35778
rect 4900 35758 4910 35778
rect 4937 35758 4993 35814
rect 5195 35758 5251 35814
rect 5277 35758 5333 35814
rect 5359 35758 5415 35814
rect 5441 35758 5497 35814
rect 5523 35758 5579 35814
rect 5605 35790 5632 35814
rect 5632 35790 5661 35814
rect 5687 35790 5700 35814
rect 5700 35790 5743 35814
rect 5769 35838 5820 35842
rect 5820 35838 5825 35842
rect 5851 35838 5907 35894
rect 5933 35838 5989 35894
rect 6015 35838 6071 35894
rect 6097 35838 6153 35894
rect 6179 35838 6235 35894
rect 6261 35838 6317 35894
rect 6343 35838 6399 35894
rect 6425 35838 6481 35894
rect 6507 35854 6552 35894
rect 6552 35854 6563 35894
rect 6589 35854 6604 35894
rect 6604 35854 6620 35894
rect 6620 35854 6645 35894
rect 6671 35854 6672 35894
rect 6672 35854 6688 35894
rect 6688 35854 6727 35894
rect 6507 35842 6563 35854
rect 6589 35842 6645 35854
rect 6671 35842 6727 35854
rect 6507 35838 6552 35842
rect 6552 35838 6563 35842
rect 6589 35838 6604 35842
rect 6604 35838 6620 35842
rect 6620 35838 6645 35842
rect 6671 35838 6672 35842
rect 6672 35838 6688 35842
rect 6688 35838 6727 35842
rect 6753 35838 6809 35894
rect 5769 35790 5820 35814
rect 5820 35790 5825 35814
rect 5605 35778 5661 35790
rect 5687 35778 5743 35790
rect 5769 35778 5825 35790
rect 5605 35758 5632 35778
rect 5632 35758 5661 35778
rect 5687 35758 5700 35778
rect 5700 35758 5743 35778
rect 4854 35726 4900 35734
rect 4900 35726 4910 35734
rect 4688 35714 4744 35726
rect 4771 35714 4827 35726
rect 4854 35714 4910 35726
rect 4688 35678 4712 35714
rect 4712 35678 4744 35714
rect 4771 35678 4780 35714
rect 4780 35678 4827 35714
rect 4854 35678 4900 35714
rect 4900 35678 4910 35714
rect 4937 35678 4993 35734
rect 5195 35678 5251 35734
rect 5277 35678 5333 35734
rect 5359 35678 5415 35734
rect 5441 35678 5497 35734
rect 5523 35678 5579 35734
rect 5605 35726 5632 35734
rect 5632 35726 5661 35734
rect 5687 35726 5700 35734
rect 5700 35726 5743 35734
rect 5769 35758 5820 35778
rect 5820 35758 5825 35778
rect 5851 35758 5907 35814
rect 5933 35758 5989 35814
rect 6015 35758 6071 35814
rect 6097 35758 6153 35814
rect 6179 35758 6235 35814
rect 6261 35758 6317 35814
rect 6343 35758 6399 35814
rect 6425 35758 6481 35814
rect 6507 35790 6552 35814
rect 6552 35790 6563 35814
rect 6589 35790 6604 35814
rect 6604 35790 6620 35814
rect 6620 35790 6645 35814
rect 6671 35790 6672 35814
rect 6672 35790 6688 35814
rect 6688 35790 6727 35814
rect 6507 35778 6563 35790
rect 6589 35778 6645 35790
rect 6671 35778 6727 35790
rect 6507 35758 6552 35778
rect 6552 35758 6563 35778
rect 6589 35758 6604 35778
rect 6604 35758 6620 35778
rect 6620 35758 6645 35778
rect 6671 35758 6672 35778
rect 6672 35758 6688 35778
rect 6688 35758 6727 35778
rect 6753 35758 6809 35814
rect 6853 35812 6909 35868
rect 6941 35812 6997 35868
rect 7029 35812 7085 35868
rect 7117 35812 7173 35868
rect 7205 35812 7261 35868
rect 7293 35812 7349 35868
rect 5769 35726 5820 35734
rect 5820 35726 5825 35734
rect 5605 35714 5661 35726
rect 5687 35714 5743 35726
rect 5769 35714 5825 35726
rect 5605 35678 5632 35714
rect 5632 35678 5661 35714
rect 5687 35678 5700 35714
rect 5700 35678 5743 35714
rect 5769 35678 5820 35714
rect 5820 35678 5825 35714
rect 5851 35678 5907 35734
rect 5933 35678 5989 35734
rect 6015 35678 6071 35734
rect 6097 35678 6153 35734
rect 6179 35678 6235 35734
rect 6261 35678 6317 35734
rect 6343 35678 6399 35734
rect 6425 35678 6481 35734
rect 6507 35726 6552 35734
rect 6552 35726 6563 35734
rect 6589 35726 6604 35734
rect 6604 35726 6620 35734
rect 6620 35726 6645 35734
rect 6671 35726 6672 35734
rect 6672 35726 6688 35734
rect 6688 35726 6727 35734
rect 6507 35714 6563 35726
rect 6589 35714 6645 35726
rect 6671 35714 6727 35726
rect 6507 35678 6552 35714
rect 6552 35678 6563 35714
rect 6589 35678 6604 35714
rect 6604 35678 6620 35714
rect 6620 35678 6645 35714
rect 6671 35678 6672 35714
rect 6672 35678 6688 35714
rect 6688 35678 6727 35714
rect 6753 35678 6809 35734
rect 6853 35730 6909 35786
rect 6941 35730 6997 35786
rect 7029 35730 7085 35786
rect 7117 35730 7173 35786
rect 7205 35730 7261 35786
rect 7293 35730 7349 35786
rect 2538 35596 2594 35652
rect 2632 35596 2688 35652
rect 2726 35596 2782 35652
rect 2820 35602 2872 35652
rect 2872 35602 2876 35652
rect 2914 35602 2924 35652
rect 2924 35602 2940 35652
rect 2940 35602 2970 35652
rect 3008 35602 3060 35652
rect 3060 35602 3064 35652
rect 2820 35596 2876 35602
rect 2914 35596 2970 35602
rect 3008 35596 3064 35602
rect 3109 35598 3165 35654
rect 3193 35598 3249 35654
rect 3277 35598 3333 35654
rect 3360 35598 3416 35654
rect 3443 35598 3499 35654
rect 3526 35598 3582 35654
rect 3609 35598 3665 35654
rect 3692 35598 3748 35654
rect 3775 35650 3831 35654
rect 3858 35650 3914 35654
rect 3941 35650 3997 35654
rect 3775 35598 3792 35650
rect 3792 35598 3831 35650
rect 3858 35598 3860 35650
rect 3860 35598 3912 35650
rect 3912 35598 3914 35650
rect 3941 35598 3980 35650
rect 3980 35598 3997 35650
rect 4024 35598 4080 35654
rect 4107 35598 4163 35654
rect 4190 35598 4246 35654
rect 4273 35598 4329 35654
rect 4356 35598 4412 35654
rect 4439 35598 4495 35654
rect 4522 35598 4578 35654
rect 4605 35598 4661 35654
rect 4688 35650 4744 35654
rect 4771 35650 4827 35654
rect 4854 35650 4910 35654
rect 4688 35598 4712 35650
rect 4712 35598 4744 35650
rect 4771 35598 4780 35650
rect 4780 35598 4827 35650
rect 4854 35598 4900 35650
rect 4900 35598 4910 35650
rect 4937 35598 4993 35654
rect 5195 35598 5251 35654
rect 5277 35598 5333 35654
rect 5359 35598 5415 35654
rect 5441 35598 5497 35654
rect 5523 35598 5579 35654
rect 5605 35650 5661 35654
rect 5687 35650 5743 35654
rect 5769 35650 5825 35654
rect 5605 35598 5632 35650
rect 5632 35598 5661 35650
rect 5687 35598 5700 35650
rect 5700 35598 5743 35650
rect 5769 35598 5820 35650
rect 5820 35598 5825 35650
rect 5851 35598 5907 35654
rect 5933 35598 5989 35654
rect 6015 35598 6071 35654
rect 6097 35598 6153 35654
rect 6179 35598 6235 35654
rect 6261 35598 6317 35654
rect 6343 35598 6399 35654
rect 6425 35598 6481 35654
rect 6507 35650 6563 35654
rect 6589 35650 6645 35654
rect 6671 35650 6727 35654
rect 6507 35598 6552 35650
rect 6552 35598 6563 35650
rect 6589 35598 6604 35650
rect 6604 35598 6620 35650
rect 6620 35598 6645 35650
rect 6671 35598 6672 35650
rect 6672 35598 6688 35650
rect 6688 35598 6727 35650
rect 6753 35598 6809 35654
rect 6853 35648 6909 35704
rect 6941 35648 6997 35704
rect 7029 35648 7085 35704
rect 7117 35648 7173 35704
rect 7205 35648 7261 35704
rect 7293 35648 7349 35704
rect 2538 35516 2594 35572
rect 2632 35516 2688 35572
rect 2726 35516 2782 35572
rect 2820 35537 2872 35572
rect 2872 35537 2876 35572
rect 2914 35537 2924 35572
rect 2924 35537 2940 35572
rect 2940 35537 2970 35572
rect 3008 35537 3060 35572
rect 3060 35537 3064 35572
rect 2820 35524 2876 35537
rect 2914 35524 2970 35537
rect 3008 35524 3064 35537
rect 2820 35516 2872 35524
rect 2872 35516 2876 35524
rect 2914 35516 2924 35524
rect 2924 35516 2940 35524
rect 2940 35516 2970 35524
rect 2538 35435 2594 35491
rect 2632 35435 2688 35491
rect 2726 35435 2782 35491
rect 2820 35472 2872 35491
rect 2872 35472 2876 35491
rect 2914 35472 2924 35491
rect 2924 35472 2940 35491
rect 2940 35472 2970 35491
rect 3008 35516 3060 35524
rect 3060 35516 3064 35524
rect 3109 35518 3165 35574
rect 3193 35518 3249 35574
rect 3277 35518 3333 35574
rect 3360 35518 3416 35574
rect 3443 35518 3499 35574
rect 3526 35518 3582 35574
rect 3609 35518 3665 35574
rect 3692 35518 3748 35574
rect 3775 35534 3792 35574
rect 3792 35534 3831 35574
rect 3858 35534 3860 35574
rect 3860 35534 3912 35574
rect 3912 35534 3914 35574
rect 3941 35534 3980 35574
rect 3980 35534 3997 35574
rect 3775 35522 3831 35534
rect 3858 35522 3914 35534
rect 3941 35522 3997 35534
rect 3775 35518 3792 35522
rect 3792 35518 3831 35522
rect 3858 35518 3860 35522
rect 3860 35518 3912 35522
rect 3912 35518 3914 35522
rect 3941 35518 3980 35522
rect 3980 35518 3997 35522
rect 4024 35518 4080 35574
rect 4107 35518 4163 35574
rect 4190 35518 4246 35574
rect 4273 35518 4329 35574
rect 4356 35518 4412 35574
rect 4439 35518 4495 35574
rect 4522 35518 4578 35574
rect 4605 35518 4661 35574
rect 4688 35534 4712 35574
rect 4712 35534 4744 35574
rect 4771 35534 4780 35574
rect 4780 35534 4827 35574
rect 4854 35534 4900 35574
rect 4900 35534 4910 35574
rect 4688 35522 4744 35534
rect 4771 35522 4827 35534
rect 4854 35522 4910 35534
rect 4688 35518 4712 35522
rect 4712 35518 4744 35522
rect 4771 35518 4780 35522
rect 4780 35518 4827 35522
rect 3008 35472 3060 35491
rect 3060 35472 3064 35491
rect 2820 35459 2876 35472
rect 2914 35459 2970 35472
rect 3008 35459 3064 35472
rect 2820 35435 2872 35459
rect 2872 35435 2876 35459
rect 2914 35435 2924 35459
rect 2924 35435 2940 35459
rect 2940 35435 2970 35459
rect 2538 35354 2594 35410
rect 2632 35354 2688 35410
rect 2726 35354 2782 35410
rect 2820 35407 2872 35410
rect 2872 35407 2876 35410
rect 2914 35407 2924 35410
rect 2924 35407 2940 35410
rect 2940 35407 2970 35410
rect 3008 35435 3060 35459
rect 3060 35435 3064 35459
rect 3109 35438 3165 35494
rect 3193 35438 3249 35494
rect 3277 35438 3333 35494
rect 3360 35438 3416 35494
rect 3443 35438 3499 35494
rect 3526 35438 3582 35494
rect 3609 35438 3665 35494
rect 3692 35438 3748 35494
rect 3775 35470 3792 35494
rect 3792 35470 3831 35494
rect 3858 35470 3860 35494
rect 3860 35470 3912 35494
rect 3912 35470 3914 35494
rect 3941 35470 3980 35494
rect 3980 35470 3997 35494
rect 3775 35458 3831 35470
rect 3858 35458 3914 35470
rect 3941 35458 3997 35470
rect 3775 35438 3792 35458
rect 3792 35438 3831 35458
rect 3858 35438 3860 35458
rect 3860 35438 3912 35458
rect 3912 35438 3914 35458
rect 3941 35438 3980 35458
rect 3980 35438 3997 35458
rect 4024 35438 4080 35494
rect 4107 35438 4163 35494
rect 4190 35438 4246 35494
rect 4273 35438 4329 35494
rect 4356 35438 4412 35494
rect 4439 35438 4495 35494
rect 4522 35438 4578 35494
rect 4605 35438 4661 35494
rect 4688 35470 4712 35494
rect 4712 35470 4744 35494
rect 4771 35470 4780 35494
rect 4780 35470 4827 35494
rect 4854 35518 4900 35522
rect 4900 35518 4910 35522
rect 4937 35518 4993 35574
rect 5195 35518 5251 35574
rect 5277 35518 5333 35574
rect 5359 35518 5415 35574
rect 5441 35518 5497 35574
rect 5523 35518 5579 35574
rect 5605 35534 5632 35574
rect 5632 35534 5661 35574
rect 5687 35534 5700 35574
rect 5700 35534 5743 35574
rect 5769 35534 5820 35574
rect 5820 35534 5825 35574
rect 5605 35522 5661 35534
rect 5687 35522 5743 35534
rect 5769 35522 5825 35534
rect 5605 35518 5632 35522
rect 5632 35518 5661 35522
rect 5687 35518 5700 35522
rect 5700 35518 5743 35522
rect 4854 35470 4900 35494
rect 4900 35470 4910 35494
rect 4688 35458 4744 35470
rect 4771 35458 4827 35470
rect 4854 35458 4910 35470
rect 4688 35438 4712 35458
rect 4712 35438 4744 35458
rect 4771 35438 4780 35458
rect 4780 35438 4827 35458
rect 3008 35407 3060 35410
rect 3060 35407 3064 35410
rect 2820 35394 2876 35407
rect 2914 35394 2970 35407
rect 3008 35394 3064 35407
rect 2820 35354 2872 35394
rect 2872 35354 2876 35394
rect 2914 35354 2924 35394
rect 2924 35354 2940 35394
rect 2940 35354 2970 35394
rect 3008 35354 3060 35394
rect 3060 35354 3064 35394
rect 3109 35358 3165 35414
rect 3193 35358 3249 35414
rect 3277 35358 3333 35414
rect 3360 35358 3416 35414
rect 3443 35358 3499 35414
rect 3526 35358 3582 35414
rect 3609 35358 3665 35414
rect 3692 35358 3748 35414
rect 3775 35406 3792 35414
rect 3792 35406 3831 35414
rect 3858 35406 3860 35414
rect 3860 35406 3912 35414
rect 3912 35406 3914 35414
rect 3941 35406 3980 35414
rect 3980 35406 3997 35414
rect 3775 35394 3831 35406
rect 3858 35394 3914 35406
rect 3941 35394 3997 35406
rect 3775 35358 3792 35394
rect 3792 35358 3831 35394
rect 3858 35358 3860 35394
rect 3860 35358 3912 35394
rect 3912 35358 3914 35394
rect 3941 35358 3980 35394
rect 3980 35358 3997 35394
rect 4024 35358 4080 35414
rect 4107 35358 4163 35414
rect 4190 35358 4246 35414
rect 4273 35358 4329 35414
rect 4356 35358 4412 35414
rect 4439 35358 4495 35414
rect 4522 35358 4578 35414
rect 4605 35358 4661 35414
rect 4688 35406 4712 35414
rect 4712 35406 4744 35414
rect 4771 35406 4780 35414
rect 4780 35406 4827 35414
rect 4854 35438 4900 35458
rect 4900 35438 4910 35458
rect 4937 35438 4993 35494
rect 5195 35438 5251 35494
rect 5277 35438 5333 35494
rect 5359 35438 5415 35494
rect 5441 35438 5497 35494
rect 5523 35438 5579 35494
rect 5605 35470 5632 35494
rect 5632 35470 5661 35494
rect 5687 35470 5700 35494
rect 5700 35470 5743 35494
rect 5769 35518 5820 35522
rect 5820 35518 5825 35522
rect 5851 35518 5907 35574
rect 5933 35518 5989 35574
rect 6015 35518 6071 35574
rect 6097 35518 6153 35574
rect 6179 35518 6235 35574
rect 6261 35518 6317 35574
rect 6343 35518 6399 35574
rect 6425 35518 6481 35574
rect 6507 35534 6552 35574
rect 6552 35534 6563 35574
rect 6589 35534 6604 35574
rect 6604 35534 6620 35574
rect 6620 35534 6645 35574
rect 6671 35534 6672 35574
rect 6672 35534 6688 35574
rect 6688 35534 6727 35574
rect 6507 35522 6563 35534
rect 6589 35522 6645 35534
rect 6671 35522 6727 35534
rect 6507 35518 6552 35522
rect 6552 35518 6563 35522
rect 6589 35518 6604 35522
rect 6604 35518 6620 35522
rect 6620 35518 6645 35522
rect 6671 35518 6672 35522
rect 6672 35518 6688 35522
rect 6688 35518 6727 35522
rect 6753 35518 6809 35574
rect 6853 35566 6909 35622
rect 6941 35566 6997 35622
rect 7029 35566 7085 35622
rect 7117 35566 7173 35622
rect 7205 35566 7261 35622
rect 7293 35566 7349 35622
rect 5769 35470 5820 35494
rect 5820 35470 5825 35494
rect 5605 35458 5661 35470
rect 5687 35458 5743 35470
rect 5769 35458 5825 35470
rect 5605 35438 5632 35458
rect 5632 35438 5661 35458
rect 5687 35438 5700 35458
rect 5700 35438 5743 35458
rect 4854 35406 4900 35414
rect 4900 35406 4910 35414
rect 4688 35394 4744 35406
rect 4771 35394 4827 35406
rect 4854 35394 4910 35406
rect 4688 35358 4712 35394
rect 4712 35358 4744 35394
rect 4771 35358 4780 35394
rect 4780 35358 4827 35394
rect 4854 35358 4900 35394
rect 4900 35358 4910 35394
rect 4937 35358 4993 35414
rect 5195 35358 5251 35414
rect 5277 35358 5333 35414
rect 5359 35358 5415 35414
rect 5441 35358 5497 35414
rect 5523 35358 5579 35414
rect 5605 35406 5632 35414
rect 5632 35406 5661 35414
rect 5687 35406 5700 35414
rect 5700 35406 5743 35414
rect 5769 35438 5820 35458
rect 5820 35438 5825 35458
rect 5851 35438 5907 35494
rect 5933 35438 5989 35494
rect 6015 35438 6071 35494
rect 6097 35438 6153 35494
rect 6179 35438 6235 35494
rect 6261 35438 6317 35494
rect 6343 35438 6399 35494
rect 6425 35438 6481 35494
rect 6507 35470 6552 35494
rect 6552 35470 6563 35494
rect 6589 35470 6604 35494
rect 6604 35470 6620 35494
rect 6620 35470 6645 35494
rect 6671 35470 6672 35494
rect 6672 35470 6688 35494
rect 6688 35470 6727 35494
rect 6507 35458 6563 35470
rect 6589 35458 6645 35470
rect 6671 35458 6727 35470
rect 6507 35438 6552 35458
rect 6552 35438 6563 35458
rect 6589 35438 6604 35458
rect 6604 35438 6620 35458
rect 6620 35438 6645 35458
rect 6671 35438 6672 35458
rect 6672 35438 6688 35458
rect 6688 35438 6727 35458
rect 6753 35438 6809 35494
rect 6853 35483 6909 35539
rect 6941 35483 6997 35539
rect 7029 35483 7085 35539
rect 7117 35483 7173 35539
rect 7205 35483 7261 35539
rect 7293 35483 7349 35539
rect 5769 35406 5820 35414
rect 5820 35406 5825 35414
rect 5605 35394 5661 35406
rect 5687 35394 5743 35406
rect 5769 35394 5825 35406
rect 5605 35358 5632 35394
rect 5632 35358 5661 35394
rect 5687 35358 5700 35394
rect 5700 35358 5743 35394
rect 5769 35358 5820 35394
rect 5820 35358 5825 35394
rect 5851 35358 5907 35414
rect 5933 35358 5989 35414
rect 6015 35358 6071 35414
rect 6097 35358 6153 35414
rect 6179 35358 6235 35414
rect 6261 35358 6317 35414
rect 6343 35358 6399 35414
rect 6425 35358 6481 35414
rect 6507 35406 6552 35414
rect 6552 35406 6563 35414
rect 6589 35406 6604 35414
rect 6604 35406 6620 35414
rect 6620 35406 6645 35414
rect 6671 35406 6672 35414
rect 6672 35406 6688 35414
rect 6688 35406 6727 35414
rect 6507 35394 6563 35406
rect 6589 35394 6645 35406
rect 6671 35394 6727 35406
rect 6507 35358 6552 35394
rect 6552 35358 6563 35394
rect 6589 35358 6604 35394
rect 6604 35358 6620 35394
rect 6620 35358 6645 35394
rect 6671 35358 6672 35394
rect 6672 35358 6688 35394
rect 6688 35358 6727 35394
rect 6753 35358 6809 35414
rect 6853 35400 6909 35456
rect 6941 35400 6997 35456
rect 7029 35400 7085 35456
rect 7117 35400 7173 35456
rect 7205 35400 7261 35456
rect 7293 35400 7349 35456
rect 2538 35273 2594 35329
rect 2632 35273 2688 35329
rect 2726 35273 2782 35329
rect 2820 35277 2872 35329
rect 2872 35277 2876 35329
rect 2914 35277 2924 35329
rect 2924 35277 2940 35329
rect 2940 35277 2970 35329
rect 3008 35277 3060 35329
rect 3060 35277 3064 35329
rect 3109 35278 3165 35334
rect 3193 35278 3249 35334
rect 3277 35278 3333 35334
rect 3360 35278 3416 35334
rect 3443 35278 3499 35334
rect 3526 35278 3582 35334
rect 3609 35278 3665 35334
rect 3692 35278 3748 35334
rect 3775 35329 3831 35334
rect 3858 35329 3914 35334
rect 3941 35329 3997 35334
rect 3775 35278 3792 35329
rect 3792 35278 3831 35329
rect 3858 35278 3860 35329
rect 3860 35278 3912 35329
rect 3912 35278 3914 35329
rect 3941 35278 3980 35329
rect 3980 35278 3997 35329
rect 4024 35278 4080 35334
rect 4107 35278 4163 35334
rect 4190 35278 4246 35334
rect 4273 35278 4329 35334
rect 4356 35278 4412 35334
rect 4439 35278 4495 35334
rect 4522 35278 4578 35334
rect 4605 35278 4661 35334
rect 4688 35329 4744 35334
rect 4771 35329 4827 35334
rect 4854 35329 4910 35334
rect 4688 35278 4712 35329
rect 4712 35278 4744 35329
rect 4771 35278 4780 35329
rect 4780 35278 4827 35329
rect 4854 35278 4900 35329
rect 4900 35278 4910 35329
rect 4937 35278 4993 35334
rect 5195 35278 5251 35334
rect 5277 35278 5333 35334
rect 5359 35278 5415 35334
rect 5441 35278 5497 35334
rect 5523 35278 5579 35334
rect 5605 35329 5661 35334
rect 5687 35329 5743 35334
rect 5769 35329 5825 35334
rect 5605 35278 5632 35329
rect 5632 35278 5661 35329
rect 5687 35278 5700 35329
rect 5700 35278 5743 35329
rect 5769 35278 5820 35329
rect 5820 35278 5825 35329
rect 5851 35278 5907 35334
rect 5933 35278 5989 35334
rect 6015 35278 6071 35334
rect 6097 35278 6153 35334
rect 6179 35278 6235 35334
rect 6261 35278 6317 35334
rect 6343 35278 6399 35334
rect 6425 35278 6481 35334
rect 6507 35329 6563 35334
rect 6589 35329 6645 35334
rect 6671 35329 6727 35334
rect 6507 35278 6552 35329
rect 6552 35278 6563 35329
rect 6589 35278 6604 35329
rect 6604 35278 6620 35329
rect 6620 35278 6645 35329
rect 6671 35278 6672 35329
rect 6672 35278 6688 35329
rect 6688 35278 6727 35329
rect 6753 35278 6809 35334
rect 6853 35317 6909 35373
rect 6941 35317 6997 35373
rect 7029 35317 7085 35373
rect 7117 35317 7173 35373
rect 7205 35317 7261 35373
rect 7293 35317 7349 35373
rect 2820 35273 2876 35277
rect 2914 35273 2970 35277
rect 3008 35273 3064 35277
rect 2538 35192 2594 35248
rect 2632 35192 2688 35248
rect 2726 35192 2782 35248
rect 2820 35212 2872 35248
rect 2872 35212 2876 35248
rect 2914 35212 2924 35248
rect 2924 35212 2940 35248
rect 2940 35212 2970 35248
rect 3008 35212 3060 35248
rect 3060 35212 3064 35248
rect 2820 35199 2876 35212
rect 2914 35199 2970 35212
rect 3008 35199 3064 35212
rect 2820 35192 2872 35199
rect 2872 35192 2876 35199
rect 2914 35192 2924 35199
rect 2924 35192 2940 35199
rect 2940 35192 2970 35199
rect 3008 35192 3060 35199
rect 3060 35192 3064 35199
rect 3109 35198 3165 35254
rect 3193 35198 3249 35254
rect 3277 35198 3333 35254
rect 3360 35198 3416 35254
rect 3443 35198 3499 35254
rect 3526 35198 3582 35254
rect 3609 35198 3665 35254
rect 3692 35198 3748 35254
rect 3775 35212 3792 35254
rect 3792 35212 3831 35254
rect 3858 35212 3860 35254
rect 3860 35212 3912 35254
rect 3912 35212 3914 35254
rect 3941 35212 3980 35254
rect 3980 35212 3997 35254
rect 3775 35199 3831 35212
rect 3858 35199 3914 35212
rect 3941 35199 3997 35212
rect 3775 35198 3792 35199
rect 3792 35198 3831 35199
rect 3858 35198 3860 35199
rect 3860 35198 3912 35199
rect 3912 35198 3914 35199
rect 3941 35198 3980 35199
rect 3980 35198 3997 35199
rect 4024 35198 4080 35254
rect 4107 35198 4163 35254
rect 4190 35198 4246 35254
rect 4273 35198 4329 35254
rect 4356 35198 4412 35254
rect 4439 35198 4495 35254
rect 4522 35198 4578 35254
rect 4605 35198 4661 35254
rect 4688 35212 4712 35254
rect 4712 35212 4744 35254
rect 4771 35212 4780 35254
rect 4780 35212 4827 35254
rect 4854 35212 4900 35254
rect 4900 35212 4910 35254
rect 4688 35199 4744 35212
rect 4771 35199 4827 35212
rect 4854 35199 4910 35212
rect 4688 35198 4712 35199
rect 4712 35198 4744 35199
rect 4771 35198 4780 35199
rect 4780 35198 4827 35199
rect 2821 35147 2872 35150
rect 2872 35147 2877 35150
rect 2914 35147 2924 35150
rect 2924 35147 2940 35150
rect 2940 35147 2970 35150
rect 3006 35147 3008 35150
rect 3008 35147 3060 35150
rect 3060 35147 3062 35150
rect 2675 35083 2731 35139
rect 2821 35134 2877 35147
rect 2914 35134 2970 35147
rect 3006 35134 3062 35147
rect 2821 35094 2872 35134
rect 2872 35094 2877 35134
rect 2914 35094 2924 35134
rect 2924 35094 2940 35134
rect 2940 35094 2970 35134
rect 3006 35094 3008 35134
rect 3008 35094 3060 35134
rect 3060 35094 3062 35134
rect 3109 35118 3165 35174
rect 3193 35118 3249 35174
rect 3277 35118 3333 35174
rect 3360 35118 3416 35174
rect 3443 35118 3499 35174
rect 3526 35118 3582 35174
rect 3609 35118 3665 35174
rect 3692 35118 3748 35174
rect 3775 35147 3792 35174
rect 3792 35147 3831 35174
rect 3858 35147 3860 35174
rect 3860 35147 3912 35174
rect 3912 35147 3914 35174
rect 3941 35147 3980 35174
rect 3980 35147 3997 35174
rect 3775 35134 3831 35147
rect 3858 35134 3914 35147
rect 3941 35134 3997 35147
rect 3775 35118 3792 35134
rect 3792 35118 3831 35134
rect 3858 35118 3860 35134
rect 3860 35118 3912 35134
rect 3912 35118 3914 35134
rect 3941 35118 3980 35134
rect 3980 35118 3997 35134
rect 4024 35118 4080 35174
rect 4107 35118 4163 35174
rect 4190 35118 4246 35174
rect 4273 35118 4329 35174
rect 4356 35118 4412 35174
rect 4439 35118 4495 35174
rect 4522 35118 4578 35174
rect 4605 35118 4661 35174
rect 4688 35147 4712 35174
rect 4712 35147 4744 35174
rect 4771 35147 4780 35174
rect 4780 35147 4827 35174
rect 4854 35198 4900 35199
rect 4900 35198 4910 35199
rect 4937 35198 4993 35254
rect 5195 35198 5251 35254
rect 5277 35198 5333 35254
rect 5359 35198 5415 35254
rect 5441 35198 5497 35254
rect 5523 35198 5579 35254
rect 5605 35212 5632 35254
rect 5632 35212 5661 35254
rect 5687 35212 5700 35254
rect 5700 35212 5743 35254
rect 5769 35212 5820 35254
rect 5820 35212 5825 35254
rect 5605 35199 5661 35212
rect 5687 35199 5743 35212
rect 5769 35199 5825 35212
rect 5605 35198 5632 35199
rect 5632 35198 5661 35199
rect 5687 35198 5700 35199
rect 5700 35198 5743 35199
rect 4854 35147 4900 35174
rect 4900 35147 4910 35174
rect 4688 35134 4744 35147
rect 4771 35134 4827 35147
rect 4854 35134 4910 35147
rect 4688 35118 4712 35134
rect 4712 35118 4744 35134
rect 4771 35118 4780 35134
rect 4780 35118 4827 35134
rect 2821 35017 2872 35058
rect 2872 35017 2877 35058
rect 2914 35017 2924 35058
rect 2924 35017 2940 35058
rect 2940 35017 2970 35058
rect 3006 35017 3008 35058
rect 3008 35017 3060 35058
rect 3060 35017 3062 35058
rect 3109 35038 3165 35094
rect 3193 35038 3249 35094
rect 3277 35038 3333 35094
rect 3360 35038 3416 35094
rect 3443 35038 3499 35094
rect 3526 35038 3582 35094
rect 3609 35038 3665 35094
rect 3692 35038 3748 35094
rect 3775 35082 3792 35094
rect 3792 35082 3831 35094
rect 3858 35082 3860 35094
rect 3860 35082 3912 35094
rect 3912 35082 3914 35094
rect 3941 35082 3980 35094
rect 3980 35082 3997 35094
rect 3775 35069 3831 35082
rect 3858 35069 3914 35082
rect 3941 35069 3997 35082
rect 3775 35038 3792 35069
rect 3792 35038 3831 35069
rect 3858 35038 3860 35069
rect 3860 35038 3912 35069
rect 3912 35038 3914 35069
rect 3941 35038 3980 35069
rect 3980 35038 3997 35069
rect 4024 35038 4080 35094
rect 4107 35038 4163 35094
rect 4190 35038 4246 35094
rect 4273 35038 4329 35094
rect 4356 35038 4412 35094
rect 4439 35038 4495 35094
rect 4522 35038 4578 35094
rect 4605 35038 4661 35094
rect 4688 35082 4712 35094
rect 4712 35082 4744 35094
rect 4771 35082 4780 35094
rect 4780 35082 4827 35094
rect 4854 35118 4900 35134
rect 4900 35118 4910 35134
rect 4937 35118 4993 35174
rect 5195 35118 5251 35174
rect 5277 35118 5333 35174
rect 5359 35118 5415 35174
rect 5441 35118 5497 35174
rect 5523 35118 5579 35174
rect 5605 35147 5632 35174
rect 5632 35147 5661 35174
rect 5687 35147 5700 35174
rect 5700 35147 5743 35174
rect 5769 35198 5820 35199
rect 5820 35198 5825 35199
rect 5851 35198 5907 35254
rect 5933 35198 5989 35254
rect 6015 35198 6071 35254
rect 6097 35198 6153 35254
rect 6179 35198 6235 35254
rect 6261 35198 6317 35254
rect 6343 35198 6399 35254
rect 6425 35198 6481 35254
rect 6507 35212 6552 35254
rect 6552 35212 6563 35254
rect 6589 35212 6604 35254
rect 6604 35212 6620 35254
rect 6620 35212 6645 35254
rect 6671 35212 6672 35254
rect 6672 35212 6688 35254
rect 6688 35212 6727 35254
rect 6507 35199 6563 35212
rect 6589 35199 6645 35212
rect 6671 35199 6727 35212
rect 6507 35198 6552 35199
rect 6552 35198 6563 35199
rect 6589 35198 6604 35199
rect 6604 35198 6620 35199
rect 6620 35198 6645 35199
rect 6671 35198 6672 35199
rect 6672 35198 6688 35199
rect 6688 35198 6727 35199
rect 6753 35198 6809 35254
rect 6853 35234 6909 35290
rect 6941 35234 6997 35290
rect 7029 35234 7085 35290
rect 7117 35234 7173 35290
rect 7205 35234 7261 35290
rect 7293 35234 7349 35290
rect 5769 35147 5820 35174
rect 5820 35147 5825 35174
rect 5605 35134 5661 35147
rect 5687 35134 5743 35147
rect 5769 35134 5825 35147
rect 5605 35118 5632 35134
rect 5632 35118 5661 35134
rect 5687 35118 5700 35134
rect 5700 35118 5743 35134
rect 4854 35082 4900 35094
rect 4900 35082 4910 35094
rect 4688 35069 4744 35082
rect 4771 35069 4827 35082
rect 4854 35069 4910 35082
rect 4688 35038 4712 35069
rect 4712 35038 4744 35069
rect 4771 35038 4780 35069
rect 4780 35038 4827 35069
rect 4854 35038 4900 35069
rect 4900 35038 4910 35069
rect 4937 35038 4993 35094
rect 5195 35038 5251 35094
rect 5277 35038 5333 35094
rect 5359 35038 5415 35094
rect 5441 35038 5497 35094
rect 5523 35038 5579 35094
rect 5605 35082 5632 35094
rect 5632 35082 5661 35094
rect 5687 35082 5700 35094
rect 5700 35082 5743 35094
rect 5769 35118 5820 35134
rect 5820 35118 5825 35134
rect 5851 35118 5907 35174
rect 5933 35118 5989 35174
rect 6015 35118 6071 35174
rect 6097 35118 6153 35174
rect 6179 35118 6235 35174
rect 6261 35118 6317 35174
rect 6343 35118 6399 35174
rect 6425 35118 6481 35174
rect 6507 35147 6552 35174
rect 6552 35147 6563 35174
rect 6589 35147 6604 35174
rect 6604 35147 6620 35174
rect 6620 35147 6645 35174
rect 6671 35147 6672 35174
rect 6672 35147 6688 35174
rect 6688 35147 6727 35174
rect 6507 35134 6563 35147
rect 6589 35134 6645 35147
rect 6671 35134 6727 35147
rect 6507 35118 6552 35134
rect 6552 35118 6563 35134
rect 6589 35118 6604 35134
rect 6604 35118 6620 35134
rect 6620 35118 6645 35134
rect 6671 35118 6672 35134
rect 6672 35118 6688 35134
rect 6688 35118 6727 35134
rect 6753 35118 6809 35174
rect 6853 35151 6909 35207
rect 6941 35151 6997 35207
rect 7029 35151 7085 35207
rect 7117 35151 7173 35207
rect 7205 35151 7261 35207
rect 7293 35151 7349 35207
rect 5769 35082 5820 35094
rect 5820 35082 5825 35094
rect 5605 35069 5661 35082
rect 5687 35069 5743 35082
rect 5769 35069 5825 35082
rect 5605 35038 5632 35069
rect 5632 35038 5661 35069
rect 5687 35038 5700 35069
rect 5700 35038 5743 35069
rect 5769 35038 5820 35069
rect 5820 35038 5825 35069
rect 5851 35038 5907 35094
rect 5933 35038 5989 35094
rect 6015 35038 6071 35094
rect 6097 35038 6153 35094
rect 6179 35038 6235 35094
rect 6261 35038 6317 35094
rect 6343 35038 6399 35094
rect 6425 35038 6481 35094
rect 6507 35082 6552 35094
rect 6552 35082 6563 35094
rect 6589 35082 6604 35094
rect 6604 35082 6620 35094
rect 6620 35082 6645 35094
rect 6671 35082 6672 35094
rect 6672 35082 6688 35094
rect 6688 35082 6727 35094
rect 6507 35069 6563 35082
rect 6589 35069 6645 35082
rect 6671 35069 6727 35082
rect 6507 35038 6552 35069
rect 6552 35038 6563 35069
rect 6589 35038 6604 35069
rect 6604 35038 6620 35069
rect 6620 35038 6645 35069
rect 6671 35038 6672 35069
rect 6672 35038 6688 35069
rect 6688 35038 6727 35069
rect 6753 35038 6809 35094
rect 6853 35068 6909 35124
rect 6941 35068 6997 35124
rect 7029 35068 7085 35124
rect 7117 35068 7173 35124
rect 7205 35068 7261 35124
rect 7293 35068 7349 35124
rect 2821 35004 2877 35017
rect 2914 35004 2970 35017
rect 3006 35004 3062 35017
rect 2821 35002 2872 35004
rect 2872 35002 2877 35004
rect 2914 35002 2924 35004
rect 2924 35002 2940 35004
rect 2940 35002 2970 35004
rect 3006 35002 3008 35004
rect 3008 35002 3060 35004
rect 3060 35002 3062 35004
rect 2821 34952 2872 34966
rect 2872 34952 2877 34966
rect 2914 34952 2924 34966
rect 2924 34952 2940 34966
rect 2940 34952 2970 34966
rect 3006 34952 3008 34966
rect 3008 34952 3060 34966
rect 3060 34952 3062 34966
rect 3109 34958 3165 35014
rect 3193 34958 3249 35014
rect 3277 34958 3333 35014
rect 3360 34958 3416 35014
rect 3443 34958 3499 35014
rect 3526 34958 3582 35014
rect 3609 34958 3665 35014
rect 3692 34958 3748 35014
rect 3775 35004 3831 35014
rect 3858 35004 3914 35014
rect 3941 35004 3997 35014
rect 3775 34958 3792 35004
rect 3792 34958 3831 35004
rect 3858 34958 3860 35004
rect 3860 34958 3912 35004
rect 3912 34958 3914 35004
rect 3941 34958 3980 35004
rect 3980 34958 3997 35004
rect 4024 34958 4080 35014
rect 4107 34958 4163 35014
rect 4190 34958 4246 35014
rect 4273 34958 4329 35014
rect 4356 34958 4412 35014
rect 4439 34958 4495 35014
rect 4522 34958 4578 35014
rect 4605 34958 4661 35014
rect 4688 35004 4744 35014
rect 4771 35004 4827 35014
rect 4854 35004 4910 35014
rect 4688 34958 4712 35004
rect 4712 34958 4744 35004
rect 4771 34958 4780 35004
rect 4780 34958 4827 35004
rect 4854 34958 4900 35004
rect 4900 34958 4910 35004
rect 4937 34958 4993 35014
rect 5195 34958 5251 35014
rect 5277 34958 5333 35014
rect 5359 34958 5415 35014
rect 5441 34958 5497 35014
rect 5523 34958 5579 35014
rect 5605 35004 5661 35014
rect 5687 35004 5743 35014
rect 5769 35004 5825 35014
rect 5605 34958 5632 35004
rect 5632 34958 5661 35004
rect 5687 34958 5700 35004
rect 5700 34958 5743 35004
rect 5769 34958 5820 35004
rect 5820 34958 5825 35004
rect 5851 34958 5907 35014
rect 5933 34958 5989 35014
rect 6015 34958 6071 35014
rect 6097 34958 6153 35014
rect 6179 34958 6235 35014
rect 6261 34958 6317 35014
rect 6343 34958 6399 35014
rect 6425 34958 6481 35014
rect 6507 35004 6563 35014
rect 6589 35004 6645 35014
rect 6671 35004 6727 35014
rect 6507 34958 6552 35004
rect 6552 34958 6563 35004
rect 6589 34958 6604 35004
rect 6604 34958 6620 35004
rect 6620 34958 6645 35004
rect 6671 34958 6672 35004
rect 6672 34958 6688 35004
rect 6688 34958 6727 35004
rect 6753 34958 6809 35014
rect 6847 34954 6903 35010
rect 6989 34954 7045 35010
rect 2821 34939 2877 34952
rect 2914 34939 2970 34952
rect 3006 34939 3062 34952
rect 2821 34910 2872 34939
rect 2872 34910 2877 34939
rect 2914 34910 2924 34939
rect 2924 34910 2940 34939
rect 2940 34910 2970 34939
rect 3006 34910 3008 34939
rect 3008 34910 3060 34939
rect 3060 34910 3062 34939
rect 3109 34878 3165 34934
rect 3193 34878 3249 34934
rect 3277 34878 3333 34934
rect 3360 34878 3416 34934
rect 3443 34878 3499 34934
rect 3526 34878 3582 34934
rect 3609 34878 3665 34934
rect 3692 34878 3748 34934
rect 3775 34887 3792 34934
rect 3792 34887 3831 34934
rect 3858 34887 3860 34934
rect 3860 34887 3912 34934
rect 3912 34887 3914 34934
rect 3941 34887 3980 34934
rect 3980 34887 3997 34934
rect 3775 34878 3831 34887
rect 3858 34878 3914 34887
rect 3941 34878 3997 34887
rect 4024 34878 4080 34934
rect 4107 34878 4163 34934
rect 4190 34878 4246 34934
rect 4273 34878 4329 34934
rect 4356 34878 4412 34934
rect 4439 34878 4495 34934
rect 4522 34878 4578 34934
rect 4605 34878 4661 34934
rect 4688 34887 4712 34934
rect 4712 34887 4744 34934
rect 4771 34887 4780 34934
rect 4780 34887 4827 34934
rect 4854 34887 4900 34934
rect 4900 34887 4910 34934
rect 4688 34878 4744 34887
rect 4771 34878 4827 34887
rect 4854 34878 4910 34887
rect 4937 34878 4993 34934
rect 5195 34878 5251 34934
rect 5277 34878 5333 34934
rect 5359 34878 5415 34934
rect 5441 34878 5497 34934
rect 5523 34878 5579 34934
rect 5605 34887 5632 34934
rect 5632 34887 5661 34934
rect 5687 34887 5700 34934
rect 5700 34887 5743 34934
rect 5769 34887 5820 34934
rect 5820 34887 5825 34934
rect 5605 34878 5661 34887
rect 5687 34878 5743 34887
rect 5769 34878 5825 34887
rect 5851 34878 5907 34934
rect 5933 34878 5989 34934
rect 6015 34878 6071 34934
rect 6097 34878 6153 34934
rect 6179 34878 6235 34934
rect 6261 34878 6317 34934
rect 6343 34878 6399 34934
rect 6425 34878 6481 34934
rect 6507 34887 6552 34934
rect 6552 34887 6563 34934
rect 6589 34887 6604 34934
rect 6604 34887 6620 34934
rect 6620 34887 6645 34934
rect 6671 34887 6672 34934
rect 6672 34887 6688 34934
rect 6688 34887 6727 34934
rect 6507 34878 6563 34887
rect 6589 34878 6645 34887
rect 6671 34878 6727 34887
rect 6753 34878 6809 34934
rect 7102 34924 7158 34980
rect 2963 34822 2992 34851
rect 2992 34822 3008 34851
rect 3008 34822 3019 34851
rect 2963 34809 3019 34822
rect 2963 34795 2992 34809
rect 2992 34795 3008 34809
rect 3008 34795 3019 34809
rect 3109 34798 3165 34854
rect 3193 34798 3249 34854
rect 3277 34798 3333 34854
rect 3360 34798 3416 34854
rect 3443 34798 3499 34854
rect 3526 34798 3582 34854
rect 3609 34798 3665 34854
rect 3692 34798 3748 34854
rect 3775 34822 3792 34854
rect 3792 34822 3831 34854
rect 3858 34822 3860 34854
rect 3860 34822 3912 34854
rect 3912 34822 3914 34854
rect 3941 34822 3980 34854
rect 3980 34822 3997 34854
rect 3775 34809 3831 34822
rect 3858 34809 3914 34822
rect 3941 34809 3997 34822
rect 3775 34798 3792 34809
rect 3792 34798 3831 34809
rect 3858 34798 3860 34809
rect 3860 34798 3912 34809
rect 3912 34798 3914 34809
rect 3941 34798 3980 34809
rect 3980 34798 3997 34809
rect 4024 34798 4080 34854
rect 4107 34798 4163 34854
rect 4190 34798 4246 34854
rect 4273 34798 4329 34854
rect 4356 34798 4412 34854
rect 4439 34798 4495 34854
rect 4522 34798 4578 34854
rect 4605 34798 4661 34854
rect 4688 34822 4712 34854
rect 4712 34822 4744 34854
rect 4771 34822 4780 34854
rect 4780 34822 4827 34854
rect 4854 34822 4900 34854
rect 4900 34822 4910 34854
rect 4688 34809 4744 34822
rect 4771 34809 4827 34822
rect 4854 34809 4910 34822
rect 4688 34798 4712 34809
rect 4712 34798 4744 34809
rect 4771 34798 4780 34809
rect 4780 34798 4827 34809
rect 3109 34718 3165 34774
rect 3193 34718 3249 34774
rect 3277 34718 3333 34774
rect 3360 34718 3416 34774
rect 3443 34718 3499 34774
rect 3526 34718 3582 34774
rect 3609 34718 3665 34774
rect 3692 34718 3748 34774
rect 3775 34757 3792 34774
rect 3792 34757 3831 34774
rect 3858 34757 3860 34774
rect 3860 34757 3912 34774
rect 3912 34757 3914 34774
rect 3941 34757 3980 34774
rect 3980 34757 3997 34774
rect 3775 34744 3831 34757
rect 3858 34744 3914 34757
rect 3941 34744 3997 34757
rect 3775 34718 3792 34744
rect 3792 34718 3831 34744
rect 3858 34718 3860 34744
rect 3860 34718 3912 34744
rect 3912 34718 3914 34744
rect 3941 34718 3980 34744
rect 3980 34718 3997 34744
rect 4024 34718 4080 34774
rect 4107 34718 4163 34774
rect 4190 34718 4246 34774
rect 4273 34718 4329 34774
rect 4356 34718 4412 34774
rect 4439 34718 4495 34774
rect 4522 34718 4578 34774
rect 4605 34718 4661 34774
rect 4688 34757 4712 34774
rect 4712 34757 4744 34774
rect 4771 34757 4780 34774
rect 4780 34757 4827 34774
rect 4854 34798 4900 34809
rect 4900 34798 4910 34809
rect 4937 34798 4993 34854
rect 5195 34798 5251 34854
rect 5277 34798 5333 34854
rect 5359 34798 5415 34854
rect 5441 34798 5497 34854
rect 5523 34798 5579 34854
rect 5605 34822 5632 34854
rect 5632 34822 5661 34854
rect 5687 34822 5700 34854
rect 5700 34822 5743 34854
rect 6847 34867 6903 34923
rect 6989 34867 7045 34923
rect 5769 34822 5820 34854
rect 5820 34822 5825 34854
rect 5605 34809 5661 34822
rect 5687 34809 5743 34822
rect 5769 34809 5825 34822
rect 5605 34798 5632 34809
rect 5632 34798 5661 34809
rect 5687 34798 5700 34809
rect 5700 34798 5743 34809
rect 4854 34757 4900 34774
rect 4900 34757 4910 34774
rect 4688 34744 4744 34757
rect 4771 34744 4827 34757
rect 4854 34744 4910 34757
rect 4688 34718 4712 34744
rect 4712 34718 4744 34744
rect 4771 34718 4780 34744
rect 4780 34718 4827 34744
rect 3109 34638 3165 34694
rect 3193 34638 3249 34694
rect 3277 34638 3333 34694
rect 3360 34638 3416 34694
rect 3443 34638 3499 34694
rect 3526 34638 3582 34694
rect 3609 34638 3665 34694
rect 3692 34638 3748 34694
rect 3775 34692 3792 34694
rect 3792 34692 3831 34694
rect 3858 34692 3860 34694
rect 3860 34692 3912 34694
rect 3912 34692 3914 34694
rect 3941 34692 3980 34694
rect 3980 34692 3997 34694
rect 3775 34679 3831 34692
rect 3858 34679 3914 34692
rect 3941 34679 3997 34692
rect 3775 34638 3792 34679
rect 3792 34638 3831 34679
rect 3858 34638 3860 34679
rect 3860 34638 3912 34679
rect 3912 34638 3914 34679
rect 3941 34638 3980 34679
rect 3980 34638 3997 34679
rect 4024 34638 4080 34694
rect 4107 34638 4163 34694
rect 4190 34638 4246 34694
rect 4273 34638 4329 34694
rect 4356 34638 4412 34694
rect 4439 34638 4495 34694
rect 4522 34638 4578 34694
rect 4605 34638 4661 34694
rect 4688 34692 4712 34694
rect 4712 34692 4744 34694
rect 4771 34692 4780 34694
rect 4780 34692 4827 34694
rect 4854 34718 4900 34744
rect 4900 34718 4910 34744
rect 4937 34718 4993 34774
rect 5195 34718 5251 34774
rect 5277 34718 5333 34774
rect 5359 34718 5415 34774
rect 5441 34718 5497 34774
rect 5523 34718 5579 34774
rect 5605 34757 5632 34774
rect 5632 34757 5661 34774
rect 5687 34757 5700 34774
rect 5700 34757 5743 34774
rect 5769 34798 5820 34809
rect 5820 34798 5825 34809
rect 5851 34798 5907 34854
rect 5933 34798 5989 34854
rect 6015 34798 6071 34854
rect 6097 34798 6153 34854
rect 6179 34798 6235 34854
rect 6261 34798 6317 34854
rect 6343 34798 6399 34854
rect 6425 34798 6481 34854
rect 6507 34822 6552 34854
rect 6552 34822 6563 34854
rect 6589 34822 6604 34854
rect 6604 34822 6620 34854
rect 6620 34822 6645 34854
rect 6671 34822 6672 34854
rect 6672 34822 6688 34854
rect 6688 34822 6727 34854
rect 6507 34809 6563 34822
rect 6589 34809 6645 34822
rect 6671 34809 6727 34822
rect 6507 34798 6552 34809
rect 6552 34798 6563 34809
rect 6589 34798 6604 34809
rect 6604 34798 6620 34809
rect 6620 34798 6645 34809
rect 6671 34798 6672 34809
rect 6672 34798 6688 34809
rect 6688 34798 6727 34809
rect 6753 34798 6809 34854
rect 6847 34779 6903 34835
rect 6989 34779 7045 34835
rect 5769 34757 5820 34774
rect 5820 34757 5825 34774
rect 5605 34744 5661 34757
rect 5687 34744 5743 34757
rect 5769 34744 5825 34757
rect 5605 34718 5632 34744
rect 5632 34718 5661 34744
rect 5687 34718 5700 34744
rect 5700 34718 5743 34744
rect 4854 34692 4900 34694
rect 4900 34692 4910 34694
rect 4688 34679 4744 34692
rect 4771 34679 4827 34692
rect 4854 34679 4910 34692
rect 4688 34638 4712 34679
rect 4712 34638 4744 34679
rect 4771 34638 4780 34679
rect 4780 34638 4827 34679
rect 4854 34638 4900 34679
rect 4900 34638 4910 34679
rect 4937 34638 4993 34694
rect 5195 34638 5251 34694
rect 5277 34638 5333 34694
rect 5359 34638 5415 34694
rect 5441 34638 5497 34694
rect 5523 34638 5579 34694
rect 5605 34692 5632 34694
rect 5632 34692 5661 34694
rect 5687 34692 5700 34694
rect 5700 34692 5743 34694
rect 5769 34718 5820 34744
rect 5820 34718 5825 34744
rect 5851 34718 5907 34774
rect 5933 34718 5989 34774
rect 6015 34718 6071 34774
rect 6097 34718 6153 34774
rect 6179 34718 6235 34774
rect 6261 34718 6317 34774
rect 6343 34718 6399 34774
rect 6425 34718 6481 34774
rect 6507 34757 6552 34774
rect 6552 34757 6563 34774
rect 6589 34757 6604 34774
rect 6604 34757 6620 34774
rect 6620 34757 6645 34774
rect 6671 34757 6672 34774
rect 6672 34757 6688 34774
rect 6688 34757 6727 34774
rect 6507 34744 6563 34757
rect 6589 34744 6645 34757
rect 6671 34744 6727 34757
rect 6507 34718 6552 34744
rect 6552 34718 6563 34744
rect 6589 34718 6604 34744
rect 6604 34718 6620 34744
rect 6620 34718 6645 34744
rect 6671 34718 6672 34744
rect 6672 34718 6688 34744
rect 6688 34718 6727 34744
rect 6753 34718 6809 34774
rect 5769 34692 5820 34694
rect 5820 34692 5825 34694
rect 5605 34679 5661 34692
rect 5687 34679 5743 34692
rect 5769 34679 5825 34692
rect 5605 34638 5632 34679
rect 5632 34638 5661 34679
rect 5687 34638 5700 34679
rect 5700 34638 5743 34679
rect 5769 34638 5820 34679
rect 5820 34638 5825 34679
rect 5851 34638 5907 34694
rect 5933 34638 5989 34694
rect 6015 34638 6071 34694
rect 6097 34638 6153 34694
rect 6179 34638 6235 34694
rect 6261 34638 6317 34694
rect 6343 34638 6399 34694
rect 6425 34638 6481 34694
rect 6507 34692 6552 34694
rect 6552 34692 6563 34694
rect 6589 34692 6604 34694
rect 6604 34692 6620 34694
rect 6620 34692 6645 34694
rect 6671 34692 6672 34694
rect 6672 34692 6688 34694
rect 6688 34692 6727 34694
rect 6507 34679 6563 34692
rect 6589 34679 6645 34692
rect 6671 34679 6727 34692
rect 6507 34638 6552 34679
rect 6552 34638 6563 34679
rect 6589 34638 6604 34679
rect 6604 34638 6620 34679
rect 6620 34638 6645 34679
rect 6671 34638 6672 34679
rect 6672 34638 6688 34679
rect 6688 34638 6727 34679
rect 6753 34638 6809 34694
rect 6847 34639 6903 34695
rect 3109 34558 3165 34614
rect 3193 34558 3249 34614
rect 3277 34558 3333 34614
rect 3360 34558 3416 34614
rect 3443 34558 3499 34614
rect 3526 34558 3582 34614
rect 3609 34558 3665 34614
rect 3692 34558 3748 34614
rect 3775 34562 3792 34614
rect 3792 34562 3831 34614
rect 3858 34562 3860 34614
rect 3860 34562 3912 34614
rect 3912 34562 3914 34614
rect 3941 34562 3980 34614
rect 3980 34562 3997 34614
rect 3775 34558 3831 34562
rect 3858 34558 3914 34562
rect 3941 34558 3997 34562
rect 4024 34558 4080 34614
rect 4107 34558 4163 34614
rect 4190 34558 4246 34614
rect 4273 34558 4329 34614
rect 4356 34558 4412 34614
rect 4439 34558 4495 34614
rect 4522 34558 4578 34614
rect 4605 34558 4661 34614
rect 4688 34562 4712 34614
rect 4712 34562 4744 34614
rect 4771 34562 4780 34614
rect 4780 34562 4827 34614
rect 4854 34562 4900 34614
rect 4900 34562 4910 34614
rect 4688 34558 4744 34562
rect 4771 34558 4827 34562
rect 4854 34558 4910 34562
rect 4937 34558 4993 34614
rect 5195 34558 5251 34614
rect 5277 34558 5333 34614
rect 5359 34558 5415 34614
rect 5441 34558 5497 34614
rect 5523 34558 5579 34614
rect 5605 34562 5632 34614
rect 5632 34562 5661 34614
rect 5687 34562 5700 34614
rect 5700 34562 5743 34614
rect 5769 34562 5820 34614
rect 5820 34562 5825 34614
rect 5605 34558 5661 34562
rect 5687 34558 5743 34562
rect 5769 34558 5825 34562
rect 5851 34558 5907 34614
rect 5933 34558 5989 34614
rect 6015 34558 6071 34614
rect 6097 34558 6153 34614
rect 6179 34558 6235 34614
rect 6261 34558 6317 34614
rect 6343 34558 6399 34614
rect 6425 34558 6481 34614
rect 6507 34562 6552 34614
rect 6552 34562 6563 34614
rect 6589 34562 6604 34614
rect 6604 34562 6620 34614
rect 6620 34562 6645 34614
rect 6671 34562 6672 34614
rect 6672 34562 6688 34614
rect 6688 34562 6727 34614
rect 6507 34558 6563 34562
rect 6589 34558 6645 34562
rect 6671 34558 6727 34562
rect 6753 34558 6809 34614
rect 8580 34173 8636 34229
rect 8661 34173 8717 34229
rect 8742 34173 8798 34229
rect 8823 34173 8879 34229
rect 8904 34225 8960 34229
rect 8985 34225 9041 34229
rect 8904 34173 8933 34225
rect 8933 34173 8959 34225
rect 8959 34173 8960 34225
rect 8985 34173 9011 34225
rect 9011 34173 9041 34225
rect 8580 34093 8636 34149
rect 8661 34093 8717 34149
rect 8742 34093 8798 34149
rect 8823 34093 8879 34149
rect 8904 34109 8933 34149
rect 8933 34109 8959 34149
rect 8959 34109 8960 34149
rect 8985 34109 9011 34149
rect 9011 34109 9041 34149
rect 8904 34097 8960 34109
rect 8985 34097 9041 34109
rect 8904 34093 8933 34097
rect 8933 34093 8959 34097
rect 8959 34093 8960 34097
rect 8985 34093 9011 34097
rect 9011 34093 9041 34097
rect 8580 34013 8636 34069
rect 8661 34013 8717 34069
rect 8742 34013 8798 34069
rect 8823 34013 8879 34069
rect 8904 34045 8933 34069
rect 8933 34045 8959 34069
rect 8959 34045 8960 34069
rect 8985 34045 9011 34069
rect 9011 34045 9041 34069
rect 8904 34033 8960 34045
rect 8985 34033 9041 34045
rect 8904 34013 8933 34033
rect 8933 34013 8959 34033
rect 8959 34013 8960 34033
rect 8985 34013 9011 34033
rect 9011 34013 9041 34033
rect 8580 33933 8636 33989
rect 8661 33933 8717 33989
rect 8742 33933 8798 33989
rect 8823 33933 8879 33989
rect 8904 33981 8933 33989
rect 8933 33981 8959 33989
rect 8959 33981 8960 33989
rect 8985 33981 9011 33989
rect 9011 33981 9041 33989
rect 8904 33969 8960 33981
rect 8985 33969 9041 33981
rect 8904 33933 8933 33969
rect 8933 33933 8959 33969
rect 8959 33933 8960 33969
rect 8985 33933 9011 33969
rect 9011 33933 9041 33969
rect 8580 33853 8636 33909
rect 8661 33853 8717 33909
rect 8742 33853 8798 33909
rect 8823 33853 8879 33909
rect 8904 33905 8960 33909
rect 8985 33905 9041 33909
rect 8904 33853 8933 33905
rect 8933 33853 8959 33905
rect 8959 33853 8960 33905
rect 8985 33853 9011 33905
rect 9011 33853 9041 33905
rect 8580 33773 8636 33829
rect 8661 33773 8717 33829
rect 8742 33773 8798 33829
rect 8823 33773 8879 33829
rect 8904 33789 8933 33829
rect 8933 33789 8959 33829
rect 8959 33789 8960 33829
rect 8985 33789 9011 33829
rect 9011 33789 9041 33829
rect 8904 33777 8960 33789
rect 8985 33777 9041 33789
rect 8904 33773 8933 33777
rect 8933 33773 8959 33777
rect 8959 33773 8960 33777
rect 8985 33773 9011 33777
rect 9011 33773 9041 33777
rect 8580 33693 8636 33749
rect 8661 33693 8717 33749
rect 8742 33693 8798 33749
rect 8823 33693 8879 33749
rect 8904 33725 8933 33749
rect 8933 33725 8959 33749
rect 8959 33725 8960 33749
rect 8985 33725 9011 33749
rect 9011 33725 9041 33749
rect 8904 33713 8960 33725
rect 8985 33713 9041 33725
rect 8904 33693 8933 33713
rect 8933 33693 8959 33713
rect 8959 33693 8960 33713
rect 8985 33693 9011 33713
rect 9011 33693 9041 33713
rect 8580 33613 8636 33669
rect 8661 33613 8717 33669
rect 8742 33613 8798 33669
rect 8823 33613 8879 33669
rect 8904 33661 8933 33669
rect 8933 33661 8959 33669
rect 8959 33661 8960 33669
rect 8985 33661 9011 33669
rect 9011 33661 9041 33669
rect 8904 33649 8960 33661
rect 8985 33649 9041 33661
rect 8904 33613 8933 33649
rect 8933 33613 8959 33649
rect 8959 33613 8960 33649
rect 8985 33613 9011 33649
rect 9011 33613 9041 33649
rect 8580 33533 8636 33589
rect 8661 33533 8717 33589
rect 8742 33533 8798 33589
rect 8823 33533 8879 33589
rect 8904 33585 8960 33589
rect 8985 33585 9041 33589
rect 8904 33533 8933 33585
rect 8933 33533 8959 33585
rect 8959 33533 8960 33585
rect 8985 33533 9011 33585
rect 9011 33533 9041 33585
rect 8580 33453 8636 33509
rect 8661 33453 8717 33509
rect 8742 33453 8798 33509
rect 8823 33453 8879 33509
rect 8904 33469 8933 33509
rect 8933 33469 8959 33509
rect 8959 33469 8960 33509
rect 8985 33469 9011 33509
rect 9011 33469 9041 33509
rect 8904 33457 8960 33469
rect 8985 33457 9041 33469
rect 8904 33453 8933 33457
rect 8933 33453 8959 33457
rect 8959 33453 8960 33457
rect 8985 33453 9011 33457
rect 9011 33453 9041 33457
rect 8580 33373 8636 33429
rect 8661 33373 8717 33429
rect 8742 33373 8798 33429
rect 8823 33373 8879 33429
rect 8904 33405 8933 33429
rect 8933 33405 8959 33429
rect 8959 33405 8960 33429
rect 8985 33405 9011 33429
rect 9011 33405 9041 33429
rect 8904 33393 8960 33405
rect 8985 33393 9041 33405
rect 8904 33373 8933 33393
rect 8933 33373 8959 33393
rect 8959 33373 8960 33393
rect 8985 33373 9011 33393
rect 9011 33373 9041 33393
rect 8580 33293 8636 33349
rect 8661 33293 8717 33349
rect 8742 33293 8798 33349
rect 8823 33293 8879 33349
rect 8904 33341 8933 33349
rect 8933 33341 8959 33349
rect 8959 33341 8960 33349
rect 8985 33341 9011 33349
rect 9011 33341 9041 33349
rect 8904 33329 8960 33341
rect 8985 33329 9041 33341
rect 8904 33293 8933 33329
rect 8933 33293 8959 33329
rect 8959 33293 8960 33329
rect 8985 33293 9011 33329
rect 9011 33293 9041 33329
rect 8580 33213 8636 33269
rect 8661 33213 8717 33269
rect 8742 33213 8798 33269
rect 8823 33213 8879 33269
rect 8904 33264 8960 33269
rect 8985 33264 9041 33269
rect 8904 33213 8933 33264
rect 8933 33213 8959 33264
rect 8959 33213 8960 33264
rect 8985 33213 9011 33264
rect 9011 33213 9041 33264
rect 8580 33133 8636 33189
rect 8661 33133 8717 33189
rect 8742 33133 8798 33189
rect 8823 33133 8879 33189
rect 8904 33147 8933 33189
rect 8933 33147 8959 33189
rect 8959 33147 8960 33189
rect 8985 33147 9011 33189
rect 9011 33147 9041 33189
rect 8904 33134 8960 33147
rect 8985 33134 9041 33147
rect 8904 33133 8933 33134
rect 8933 33133 8959 33134
rect 8959 33133 8960 33134
rect 8985 33133 9011 33134
rect 9011 33133 9041 33134
rect 8580 33053 8636 33109
rect 8661 33053 8717 33109
rect 8742 33053 8798 33109
rect 8823 33053 8879 33109
rect 8904 33082 8933 33109
rect 8933 33082 8959 33109
rect 8959 33082 8960 33109
rect 8985 33082 9011 33109
rect 9011 33082 9041 33109
rect 8904 33069 8960 33082
rect 8985 33069 9041 33082
rect 8904 33053 8933 33069
rect 8933 33053 8959 33069
rect 8959 33053 8960 33069
rect 8985 33053 9011 33069
rect 9011 33053 9041 33069
rect 8580 32973 8636 33029
rect 8661 32973 8717 33029
rect 8742 32973 8798 33029
rect 8823 32973 8879 33029
rect 8904 33017 8933 33029
rect 8933 33017 8959 33029
rect 8959 33017 8960 33029
rect 8985 33017 9011 33029
rect 9011 33017 9041 33029
rect 8904 33004 8960 33017
rect 8985 33004 9041 33017
rect 8904 32973 8933 33004
rect 8933 32973 8959 33004
rect 8959 32973 8960 33004
rect 8985 32973 9011 33004
rect 9011 32973 9041 33004
rect 8580 32893 8636 32949
rect 8661 32893 8717 32949
rect 8742 32893 8798 32949
rect 8823 32893 8879 32949
rect 8904 32939 8960 32949
rect 8985 32939 9041 32949
rect 8904 32893 8933 32939
rect 8933 32893 8959 32939
rect 8959 32893 8960 32939
rect 8985 32893 9011 32939
rect 9011 32893 9041 32939
rect 8580 32813 8636 32869
rect 8661 32813 8717 32869
rect 8742 32813 8798 32869
rect 8823 32813 8879 32869
rect 8904 32822 8933 32869
rect 8933 32822 8959 32869
rect 8959 32822 8960 32869
rect 8985 32822 9011 32869
rect 9011 32822 9041 32869
rect 8904 32813 8960 32822
rect 8985 32813 9041 32822
rect 8580 32733 8636 32789
rect 8661 32733 8717 32789
rect 8742 32733 8798 32789
rect 8823 32733 8879 32789
rect 8904 32757 8933 32789
rect 8933 32757 8959 32789
rect 8959 32757 8960 32789
rect 8985 32757 9011 32789
rect 9011 32757 9041 32789
rect 8904 32744 8960 32757
rect 8985 32744 9041 32757
rect 8904 32733 8933 32744
rect 8933 32733 8959 32744
rect 8959 32733 8960 32744
rect 8985 32733 9011 32744
rect 9011 32733 9041 32744
rect 8580 32653 8636 32709
rect 8661 32653 8717 32709
rect 8742 32653 8798 32709
rect 8823 32653 8879 32709
rect 8904 32692 8933 32709
rect 8933 32692 8959 32709
rect 8959 32692 8960 32709
rect 8985 32692 9011 32709
rect 9011 32692 9041 32709
rect 8904 32679 8960 32692
rect 8985 32679 9041 32692
rect 8904 32653 8933 32679
rect 8933 32653 8959 32679
rect 8959 32653 8960 32679
rect 8985 32653 9011 32679
rect 9011 32653 9041 32679
rect 8580 32573 8636 32629
rect 8661 32573 8717 32629
rect 8742 32573 8798 32629
rect 8823 32573 8879 32629
rect 8904 32627 8933 32629
rect 8933 32627 8959 32629
rect 8959 32627 8960 32629
rect 8985 32627 9011 32629
rect 9011 32627 9041 32629
rect 8904 32614 8960 32627
rect 8985 32614 9041 32627
rect 8904 32573 8933 32614
rect 8933 32573 8959 32614
rect 8959 32573 8960 32614
rect 8985 32573 9011 32614
rect 9011 32573 9041 32614
rect 8580 32493 8636 32549
rect 8661 32493 8717 32549
rect 8742 32493 8798 32549
rect 8823 32493 8879 32549
rect 8904 32497 8933 32549
rect 8933 32497 8959 32549
rect 8959 32497 8960 32549
rect 8985 32497 9011 32549
rect 9011 32497 9041 32549
rect 8904 32493 8960 32497
rect 8985 32493 9041 32497
rect 9066 32493 9762 34229
rect 10666 34225 10722 34229
rect 10747 34225 10803 34229
rect 10828 34225 10884 34229
rect 10666 34173 10721 34225
rect 10721 34173 10722 34225
rect 10747 34173 10773 34225
rect 10773 34173 10799 34225
rect 10799 34173 10803 34225
rect 10828 34173 10851 34225
rect 10851 34173 10884 34225
rect 10909 34173 10965 34229
rect 10990 34173 11046 34229
rect 11071 34173 11127 34229
rect 11152 34225 11848 34229
rect 11152 34173 11641 34225
rect 11641 34173 11693 34225
rect 11693 34173 11719 34225
rect 11719 34173 11771 34225
rect 11771 34173 11848 34225
rect 11152 34161 11848 34173
rect 10666 34109 10721 34149
rect 10721 34109 10722 34149
rect 10747 34109 10773 34149
rect 10773 34109 10799 34149
rect 10799 34109 10803 34149
rect 10828 34109 10851 34149
rect 10851 34109 10884 34149
rect 10666 34097 10722 34109
rect 10747 34097 10803 34109
rect 10828 34097 10884 34109
rect 10666 34093 10721 34097
rect 10721 34093 10722 34097
rect 10747 34093 10773 34097
rect 10773 34093 10799 34097
rect 10799 34093 10803 34097
rect 10828 34093 10851 34097
rect 10851 34093 10884 34097
rect 10909 34093 10965 34149
rect 10990 34093 11046 34149
rect 11071 34093 11127 34149
rect 11152 34109 11641 34161
rect 11641 34109 11693 34161
rect 11693 34109 11719 34161
rect 11719 34109 11771 34161
rect 11771 34109 11848 34161
rect 11152 34097 11848 34109
rect 10666 34045 10721 34069
rect 10721 34045 10722 34069
rect 10747 34045 10773 34069
rect 10773 34045 10799 34069
rect 10799 34045 10803 34069
rect 10828 34045 10851 34069
rect 10851 34045 10884 34069
rect 10666 34033 10722 34045
rect 10747 34033 10803 34045
rect 10828 34033 10884 34045
rect 10666 34013 10721 34033
rect 10721 34013 10722 34033
rect 10747 34013 10773 34033
rect 10773 34013 10799 34033
rect 10799 34013 10803 34033
rect 10828 34013 10851 34033
rect 10851 34013 10884 34033
rect 10909 34013 10965 34069
rect 10990 34013 11046 34069
rect 11071 34013 11127 34069
rect 11152 34045 11641 34097
rect 11641 34045 11693 34097
rect 11693 34045 11719 34097
rect 11719 34045 11771 34097
rect 11771 34045 11848 34097
rect 11152 34033 11848 34045
rect 10666 33981 10721 33989
rect 10721 33981 10722 33989
rect 10747 33981 10773 33989
rect 10773 33981 10799 33989
rect 10799 33981 10803 33989
rect 10828 33981 10851 33989
rect 10851 33981 10884 33989
rect 10666 33969 10722 33981
rect 10747 33969 10803 33981
rect 10828 33969 10884 33981
rect 10666 33933 10721 33969
rect 10721 33933 10722 33969
rect 10747 33933 10773 33969
rect 10773 33933 10799 33969
rect 10799 33933 10803 33969
rect 10828 33933 10851 33969
rect 10851 33933 10884 33969
rect 10909 33933 10965 33989
rect 10990 33933 11046 33989
rect 11071 33933 11127 33989
rect 11152 33981 11641 34033
rect 11641 33981 11693 34033
rect 11693 33981 11719 34033
rect 11719 33981 11771 34033
rect 11771 33981 11848 34033
rect 11152 33969 11848 33981
rect 11152 33917 11641 33969
rect 11641 33917 11693 33969
rect 11693 33917 11719 33969
rect 11719 33917 11771 33969
rect 11771 33917 11848 33969
rect 10666 33905 10722 33909
rect 10747 33905 10803 33909
rect 10828 33905 10884 33909
rect 10666 33853 10721 33905
rect 10721 33853 10722 33905
rect 10747 33853 10773 33905
rect 10773 33853 10799 33905
rect 10799 33853 10803 33905
rect 10828 33853 10851 33905
rect 10851 33853 10884 33905
rect 10909 33853 10965 33909
rect 10990 33853 11046 33909
rect 11071 33853 11127 33909
rect 11152 33905 11848 33917
rect 11152 33853 11641 33905
rect 11641 33853 11693 33905
rect 11693 33853 11719 33905
rect 11719 33853 11771 33905
rect 11771 33853 11848 33905
rect 11152 33841 11848 33853
rect 10666 33789 10721 33829
rect 10721 33789 10722 33829
rect 10747 33789 10773 33829
rect 10773 33789 10799 33829
rect 10799 33789 10803 33829
rect 10828 33789 10851 33829
rect 10851 33789 10884 33829
rect 10666 33777 10722 33789
rect 10747 33777 10803 33789
rect 10828 33777 10884 33789
rect 10666 33773 10721 33777
rect 10721 33773 10722 33777
rect 10747 33773 10773 33777
rect 10773 33773 10799 33777
rect 10799 33773 10803 33777
rect 10828 33773 10851 33777
rect 10851 33773 10884 33777
rect 10909 33773 10965 33829
rect 10990 33773 11046 33829
rect 11071 33773 11127 33829
rect 11152 33789 11641 33841
rect 11641 33789 11693 33841
rect 11693 33789 11719 33841
rect 11719 33789 11771 33841
rect 11771 33789 11848 33841
rect 11152 33777 11848 33789
rect 10666 33725 10721 33749
rect 10721 33725 10722 33749
rect 10747 33725 10773 33749
rect 10773 33725 10799 33749
rect 10799 33725 10803 33749
rect 10828 33725 10851 33749
rect 10851 33725 10884 33749
rect 10666 33713 10722 33725
rect 10747 33713 10803 33725
rect 10828 33713 10884 33725
rect 10666 33693 10721 33713
rect 10721 33693 10722 33713
rect 10747 33693 10773 33713
rect 10773 33693 10799 33713
rect 10799 33693 10803 33713
rect 10828 33693 10851 33713
rect 10851 33693 10884 33713
rect 10909 33693 10965 33749
rect 10990 33693 11046 33749
rect 11071 33693 11127 33749
rect 11152 33725 11641 33777
rect 11641 33725 11693 33777
rect 11693 33725 11719 33777
rect 11719 33725 11771 33777
rect 11771 33725 11848 33777
rect 11152 33713 11848 33725
rect 10666 33661 10721 33669
rect 10721 33661 10722 33669
rect 10747 33661 10773 33669
rect 10773 33661 10799 33669
rect 10799 33661 10803 33669
rect 10828 33661 10851 33669
rect 10851 33661 10884 33669
rect 10666 33649 10722 33661
rect 10747 33649 10803 33661
rect 10828 33649 10884 33661
rect 10666 33613 10721 33649
rect 10721 33613 10722 33649
rect 10747 33613 10773 33649
rect 10773 33613 10799 33649
rect 10799 33613 10803 33649
rect 10828 33613 10851 33649
rect 10851 33613 10884 33649
rect 10909 33613 10965 33669
rect 10990 33613 11046 33669
rect 11071 33613 11127 33669
rect 11152 33661 11641 33713
rect 11641 33661 11693 33713
rect 11693 33661 11719 33713
rect 11719 33661 11771 33713
rect 11771 33661 11848 33713
rect 11152 33649 11848 33661
rect 11152 33597 11641 33649
rect 11641 33597 11693 33649
rect 11693 33597 11719 33649
rect 11719 33597 11771 33649
rect 11771 33597 11848 33649
rect 10666 33585 10722 33589
rect 10747 33585 10803 33589
rect 10828 33585 10884 33589
rect 10666 33533 10721 33585
rect 10721 33533 10722 33585
rect 10747 33533 10773 33585
rect 10773 33533 10799 33585
rect 10799 33533 10803 33585
rect 10828 33533 10851 33585
rect 10851 33533 10884 33585
rect 10909 33533 10965 33589
rect 10990 33533 11046 33589
rect 11071 33533 11127 33589
rect 11152 33585 11848 33597
rect 11152 33533 11641 33585
rect 11641 33533 11693 33585
rect 11693 33533 11719 33585
rect 11719 33533 11771 33585
rect 11771 33533 11848 33585
rect 11152 33521 11848 33533
rect 10666 33469 10721 33509
rect 10721 33469 10722 33509
rect 10747 33469 10773 33509
rect 10773 33469 10799 33509
rect 10799 33469 10803 33509
rect 10828 33469 10851 33509
rect 10851 33469 10884 33509
rect 10666 33457 10722 33469
rect 10747 33457 10803 33469
rect 10828 33457 10884 33469
rect 10666 33453 10721 33457
rect 10721 33453 10722 33457
rect 10747 33453 10773 33457
rect 10773 33453 10799 33457
rect 10799 33453 10803 33457
rect 10828 33453 10851 33457
rect 10851 33453 10884 33457
rect 10909 33453 10965 33509
rect 10990 33453 11046 33509
rect 11071 33453 11127 33509
rect 11152 33469 11641 33521
rect 11641 33469 11693 33521
rect 11693 33469 11719 33521
rect 11719 33469 11771 33521
rect 11771 33469 11848 33521
rect 11152 33457 11848 33469
rect 10666 33405 10721 33429
rect 10721 33405 10722 33429
rect 10747 33405 10773 33429
rect 10773 33405 10799 33429
rect 10799 33405 10803 33429
rect 10828 33405 10851 33429
rect 10851 33405 10884 33429
rect 10666 33393 10722 33405
rect 10747 33393 10803 33405
rect 10828 33393 10884 33405
rect 10666 33373 10721 33393
rect 10721 33373 10722 33393
rect 10747 33373 10773 33393
rect 10773 33373 10799 33393
rect 10799 33373 10803 33393
rect 10828 33373 10851 33393
rect 10851 33373 10884 33393
rect 10909 33373 10965 33429
rect 10990 33373 11046 33429
rect 11071 33373 11127 33429
rect 11152 33405 11641 33457
rect 11641 33405 11693 33457
rect 11693 33405 11719 33457
rect 11719 33405 11771 33457
rect 11771 33405 11848 33457
rect 11152 33393 11848 33405
rect 10666 33341 10721 33349
rect 10721 33341 10722 33349
rect 10747 33341 10773 33349
rect 10773 33341 10799 33349
rect 10799 33341 10803 33349
rect 10828 33341 10851 33349
rect 10851 33341 10884 33349
rect 10666 33329 10722 33341
rect 10747 33329 10803 33341
rect 10828 33329 10884 33341
rect 10666 33293 10721 33329
rect 10721 33293 10722 33329
rect 10747 33293 10773 33329
rect 10773 33293 10799 33329
rect 10799 33293 10803 33329
rect 10828 33293 10851 33329
rect 10851 33293 10884 33329
rect 10909 33293 10965 33349
rect 10990 33293 11046 33349
rect 11071 33293 11127 33349
rect 11152 33341 11641 33393
rect 11641 33341 11693 33393
rect 11693 33341 11719 33393
rect 11719 33341 11771 33393
rect 11771 33341 11848 33393
rect 11152 33329 11848 33341
rect 11152 33277 11641 33329
rect 11641 33277 11693 33329
rect 11693 33277 11719 33329
rect 11719 33277 11771 33329
rect 11771 33277 11848 33329
rect 10666 33264 10722 33269
rect 10747 33264 10803 33269
rect 10828 33264 10884 33269
rect 10666 33213 10721 33264
rect 10721 33213 10722 33264
rect 10747 33213 10773 33264
rect 10773 33213 10799 33264
rect 10799 33213 10803 33264
rect 10828 33213 10851 33264
rect 10851 33213 10884 33264
rect 10909 33213 10965 33269
rect 10990 33213 11046 33269
rect 11071 33213 11127 33269
rect 11152 33264 11848 33277
rect 11152 33212 11641 33264
rect 11641 33212 11693 33264
rect 11693 33212 11719 33264
rect 11719 33212 11771 33264
rect 11771 33212 11848 33264
rect 11152 33199 11848 33212
rect 10666 33147 10721 33189
rect 10721 33147 10722 33189
rect 10747 33147 10773 33189
rect 10773 33147 10799 33189
rect 10799 33147 10803 33189
rect 10828 33147 10851 33189
rect 10851 33147 10884 33189
rect 10666 33134 10722 33147
rect 10747 33134 10803 33147
rect 10828 33134 10884 33147
rect 10666 33133 10721 33134
rect 10721 33133 10722 33134
rect 10747 33133 10773 33134
rect 10773 33133 10799 33134
rect 10799 33133 10803 33134
rect 10828 33133 10851 33134
rect 10851 33133 10884 33134
rect 10909 33133 10965 33189
rect 10990 33133 11046 33189
rect 11071 33133 11127 33189
rect 11152 33147 11641 33199
rect 11641 33147 11693 33199
rect 11693 33147 11719 33199
rect 11719 33147 11771 33199
rect 11771 33147 11848 33199
rect 11152 33134 11848 33147
rect 10666 33082 10721 33109
rect 10721 33082 10722 33109
rect 10747 33082 10773 33109
rect 10773 33082 10799 33109
rect 10799 33082 10803 33109
rect 10828 33082 10851 33109
rect 10851 33082 10884 33109
rect 10666 33069 10722 33082
rect 10747 33069 10803 33082
rect 10828 33069 10884 33082
rect 10666 33053 10721 33069
rect 10721 33053 10722 33069
rect 10747 33053 10773 33069
rect 10773 33053 10799 33069
rect 10799 33053 10803 33069
rect 10828 33053 10851 33069
rect 10851 33053 10884 33069
rect 10909 33053 10965 33109
rect 10990 33053 11046 33109
rect 11071 33053 11127 33109
rect 11152 33082 11641 33134
rect 11641 33082 11693 33134
rect 11693 33082 11719 33134
rect 11719 33082 11771 33134
rect 11771 33082 11848 33134
rect 11152 33069 11848 33082
rect 10666 33017 10721 33029
rect 10721 33017 10722 33029
rect 10747 33017 10773 33029
rect 10773 33017 10799 33029
rect 10799 33017 10803 33029
rect 10828 33017 10851 33029
rect 10851 33017 10884 33029
rect 10666 33004 10722 33017
rect 10747 33004 10803 33017
rect 10828 33004 10884 33017
rect 10666 32973 10721 33004
rect 10721 32973 10722 33004
rect 10747 32973 10773 33004
rect 10773 32973 10799 33004
rect 10799 32973 10803 33004
rect 10828 32973 10851 33004
rect 10851 32973 10884 33004
rect 10909 32973 10965 33029
rect 10990 32973 11046 33029
rect 11071 32973 11127 33029
rect 11152 33017 11641 33069
rect 11641 33017 11693 33069
rect 11693 33017 11719 33069
rect 11719 33017 11771 33069
rect 11771 33017 11848 33069
rect 11152 33004 11848 33017
rect 11152 32952 11641 33004
rect 11641 32952 11693 33004
rect 11693 32952 11719 33004
rect 11719 32952 11771 33004
rect 11771 32952 11848 33004
rect 10666 32939 10722 32949
rect 10747 32939 10803 32949
rect 10828 32939 10884 32949
rect 10666 32893 10721 32939
rect 10721 32893 10722 32939
rect 10747 32893 10773 32939
rect 10773 32893 10799 32939
rect 10799 32893 10803 32939
rect 10828 32893 10851 32939
rect 10851 32893 10884 32939
rect 10909 32893 10965 32949
rect 10990 32893 11046 32949
rect 11071 32893 11127 32949
rect 11152 32939 11848 32952
rect 11152 32887 11641 32939
rect 11641 32887 11693 32939
rect 11693 32887 11719 32939
rect 11719 32887 11771 32939
rect 11771 32887 11848 32939
rect 11152 32874 11848 32887
rect 10666 32822 10721 32869
rect 10721 32822 10722 32869
rect 10747 32822 10773 32869
rect 10773 32822 10799 32869
rect 10799 32822 10803 32869
rect 10828 32822 10851 32869
rect 10851 32822 10884 32869
rect 10666 32813 10722 32822
rect 10747 32813 10803 32822
rect 10828 32813 10884 32822
rect 10909 32813 10965 32869
rect 10990 32813 11046 32869
rect 11071 32813 11127 32869
rect 11152 32822 11641 32874
rect 11641 32822 11693 32874
rect 11693 32822 11719 32874
rect 11719 32822 11771 32874
rect 11771 32822 11848 32874
rect 11152 32809 11848 32822
rect 10666 32757 10721 32789
rect 10721 32757 10722 32789
rect 10747 32757 10773 32789
rect 10773 32757 10799 32789
rect 10799 32757 10803 32789
rect 10828 32757 10851 32789
rect 10851 32757 10884 32789
rect 10666 32744 10722 32757
rect 10747 32744 10803 32757
rect 10828 32744 10884 32757
rect 10666 32733 10721 32744
rect 10721 32733 10722 32744
rect 10747 32733 10773 32744
rect 10773 32733 10799 32744
rect 10799 32733 10803 32744
rect 10828 32733 10851 32744
rect 10851 32733 10884 32744
rect 10909 32733 10965 32789
rect 10990 32733 11046 32789
rect 11071 32733 11127 32789
rect 11152 32757 11641 32809
rect 11641 32757 11693 32809
rect 11693 32757 11719 32809
rect 11719 32757 11771 32809
rect 11771 32757 11848 32809
rect 11152 32744 11848 32757
rect 10666 32692 10721 32709
rect 10721 32692 10722 32709
rect 10747 32692 10773 32709
rect 10773 32692 10799 32709
rect 10799 32692 10803 32709
rect 10828 32692 10851 32709
rect 10851 32692 10884 32709
rect 10666 32679 10722 32692
rect 10747 32679 10803 32692
rect 10828 32679 10884 32692
rect 10666 32653 10721 32679
rect 10721 32653 10722 32679
rect 10747 32653 10773 32679
rect 10773 32653 10799 32679
rect 10799 32653 10803 32679
rect 10828 32653 10851 32679
rect 10851 32653 10884 32679
rect 10909 32653 10965 32709
rect 10990 32653 11046 32709
rect 11071 32653 11127 32709
rect 11152 32692 11641 32744
rect 11641 32692 11693 32744
rect 11693 32692 11719 32744
rect 11719 32692 11771 32744
rect 11771 32692 11848 32744
rect 11152 32679 11848 32692
rect 10666 32627 10721 32629
rect 10721 32627 10722 32629
rect 10747 32627 10773 32629
rect 10773 32627 10799 32629
rect 10799 32627 10803 32629
rect 10828 32627 10851 32629
rect 10851 32627 10884 32629
rect 10666 32614 10722 32627
rect 10747 32614 10803 32627
rect 10828 32614 10884 32627
rect 10666 32573 10721 32614
rect 10721 32573 10722 32614
rect 10747 32573 10773 32614
rect 10773 32573 10799 32614
rect 10799 32573 10803 32614
rect 10828 32573 10851 32614
rect 10851 32573 10884 32614
rect 10909 32573 10965 32629
rect 10990 32573 11046 32629
rect 11071 32573 11127 32629
rect 11152 32627 11641 32679
rect 11641 32627 11693 32679
rect 11693 32627 11719 32679
rect 11719 32627 11771 32679
rect 11771 32627 11848 32679
rect 11152 32614 11848 32627
rect 11152 32562 11641 32614
rect 11641 32562 11693 32614
rect 11693 32562 11719 32614
rect 11719 32562 11771 32614
rect 11771 32562 11848 32614
rect 11152 32549 11848 32562
rect 10666 32497 10721 32549
rect 10721 32497 10722 32549
rect 10747 32497 10773 32549
rect 10773 32497 10799 32549
rect 10799 32497 10803 32549
rect 10828 32497 10851 32549
rect 10851 32497 10884 32549
rect 10666 32493 10722 32497
rect 10747 32493 10803 32497
rect 10828 32493 10884 32497
rect 10909 32493 10965 32549
rect 10990 32493 11046 32549
rect 11071 32493 11127 32549
rect 11152 32497 11641 32549
rect 11641 32497 11693 32549
rect 11693 32497 11719 32549
rect 11719 32497 11771 32549
rect 11771 32497 11848 32549
rect 11152 32493 11848 32497
rect 3109 31638 3165 31694
rect 3190 31638 3246 31694
rect 3271 31638 3327 31694
rect 3352 31638 3408 31694
rect 3433 31638 3489 31694
rect 3514 31690 4290 31694
rect 3514 31638 3792 31690
rect 3792 31638 3844 31690
rect 3844 31638 3860 31690
rect 3860 31638 3912 31690
rect 3912 31638 3928 31690
rect 3928 31638 3980 31690
rect 3980 31638 4290 31690
rect 5195 31638 5251 31694
rect 5276 31638 5332 31694
rect 5357 31638 5413 31694
rect 5438 31638 5494 31694
rect 5519 31638 5575 31694
rect 5600 31690 6376 31694
rect 5600 31638 5632 31690
rect 5632 31638 5684 31690
rect 5684 31638 5700 31690
rect 5700 31638 5752 31690
rect 5752 31638 5768 31690
rect 5768 31638 5820 31690
rect 5820 31638 6376 31690
rect 3514 31626 4290 31638
rect 5600 31626 6376 31638
rect 3109 31558 3165 31614
rect 3190 31558 3246 31614
rect 3271 31558 3327 31614
rect 3352 31558 3408 31614
rect 3433 31558 3489 31614
rect 3514 31574 3792 31626
rect 3792 31574 3844 31626
rect 3844 31574 3860 31626
rect 3860 31574 3912 31626
rect 3912 31574 3928 31626
rect 3928 31574 3980 31626
rect 3980 31574 4290 31626
rect 3514 31562 4290 31574
rect 3109 31478 3165 31534
rect 3190 31478 3246 31534
rect 3271 31478 3327 31534
rect 3352 31478 3408 31534
rect 3433 31478 3489 31534
rect 3514 31510 3792 31562
rect 3792 31510 3844 31562
rect 3844 31510 3860 31562
rect 3860 31510 3912 31562
rect 3912 31510 3928 31562
rect 3928 31510 3980 31562
rect 3980 31510 4290 31562
rect 5195 31558 5251 31614
rect 5276 31558 5332 31614
rect 5357 31558 5413 31614
rect 5438 31558 5494 31614
rect 5519 31558 5575 31614
rect 5600 31574 5632 31626
rect 5632 31574 5684 31626
rect 5684 31574 5700 31626
rect 5700 31574 5752 31626
rect 5752 31574 5768 31626
rect 5768 31574 5820 31626
rect 5820 31574 6376 31626
rect 5600 31562 6376 31574
rect 3514 31498 4290 31510
rect 3109 31398 3165 31454
rect 3190 31398 3246 31454
rect 3271 31398 3327 31454
rect 3352 31398 3408 31454
rect 3433 31398 3489 31454
rect 3514 31446 3792 31498
rect 3792 31446 3844 31498
rect 3844 31446 3860 31498
rect 3860 31446 3912 31498
rect 3912 31446 3928 31498
rect 3928 31446 3980 31498
rect 3980 31446 4290 31498
rect 5195 31478 5251 31534
rect 5276 31478 5332 31534
rect 5357 31478 5413 31534
rect 5438 31478 5494 31534
rect 5519 31478 5575 31534
rect 5600 31510 5632 31562
rect 5632 31510 5684 31562
rect 5684 31510 5700 31562
rect 5700 31510 5752 31562
rect 5752 31510 5768 31562
rect 5768 31510 5820 31562
rect 5820 31510 6376 31562
rect 5600 31498 6376 31510
rect 3514 31434 4290 31446
rect 3514 31382 3792 31434
rect 3792 31382 3844 31434
rect 3844 31382 3860 31434
rect 3860 31382 3912 31434
rect 3912 31382 3928 31434
rect 3928 31382 3980 31434
rect 3980 31382 4290 31434
rect 5195 31398 5251 31454
rect 5276 31398 5332 31454
rect 5357 31398 5413 31454
rect 5438 31398 5494 31454
rect 5519 31398 5575 31454
rect 5600 31446 5632 31498
rect 5632 31446 5684 31498
rect 5684 31446 5700 31498
rect 5700 31446 5752 31498
rect 5752 31446 5768 31498
rect 5768 31446 5820 31498
rect 5820 31446 6376 31498
rect 5600 31434 6376 31446
rect 5600 31382 5632 31434
rect 5632 31382 5684 31434
rect 5684 31382 5700 31434
rect 5700 31382 5752 31434
rect 5752 31382 5768 31434
rect 5768 31382 5820 31434
rect 5820 31382 6376 31434
rect 3109 31318 3165 31374
rect 3190 31318 3246 31374
rect 3271 31318 3327 31374
rect 3352 31318 3408 31374
rect 3433 31318 3489 31374
rect 3514 31370 4290 31382
rect 3514 31318 3792 31370
rect 3792 31318 3844 31370
rect 3844 31318 3860 31370
rect 3860 31318 3912 31370
rect 3912 31318 3928 31370
rect 3928 31318 3980 31370
rect 3980 31318 4290 31370
rect 5195 31318 5251 31374
rect 5276 31318 5332 31374
rect 5357 31318 5413 31374
rect 5438 31318 5494 31374
rect 5519 31318 5575 31374
rect 5600 31370 6376 31382
rect 5600 31318 5632 31370
rect 5632 31318 5684 31370
rect 5684 31318 5700 31370
rect 5700 31318 5752 31370
rect 5752 31318 5768 31370
rect 5768 31318 5820 31370
rect 5820 31318 6376 31370
rect 3514 31306 4290 31318
rect 5600 31306 6376 31318
rect 3109 31238 3165 31294
rect 3190 31238 3246 31294
rect 3271 31238 3327 31294
rect 3352 31238 3408 31294
rect 3433 31238 3489 31294
rect 3514 31254 3792 31306
rect 3792 31254 3844 31306
rect 3844 31254 3860 31306
rect 3860 31254 3912 31306
rect 3912 31254 3928 31306
rect 3928 31254 3980 31306
rect 3980 31254 4290 31306
rect 3514 31242 4290 31254
rect 3109 31158 3165 31214
rect 3190 31158 3246 31214
rect 3271 31158 3327 31214
rect 3352 31158 3408 31214
rect 3433 31158 3489 31214
rect 3514 31190 3792 31242
rect 3792 31190 3844 31242
rect 3844 31190 3860 31242
rect 3860 31190 3912 31242
rect 3912 31190 3928 31242
rect 3928 31190 3980 31242
rect 3980 31190 4290 31242
rect 5195 31238 5251 31294
rect 5276 31238 5332 31294
rect 5357 31238 5413 31294
rect 5438 31238 5494 31294
rect 5519 31238 5575 31294
rect 5600 31254 5632 31306
rect 5632 31254 5684 31306
rect 5684 31254 5700 31306
rect 5700 31254 5752 31306
rect 5752 31254 5768 31306
rect 5768 31254 5820 31306
rect 5820 31254 6376 31306
rect 5600 31242 6376 31254
rect 3514 31178 4290 31190
rect 3109 31078 3165 31134
rect 3190 31078 3246 31134
rect 3271 31078 3327 31134
rect 3352 31078 3408 31134
rect 3433 31078 3489 31134
rect 3514 31126 3792 31178
rect 3792 31126 3844 31178
rect 3844 31126 3860 31178
rect 3860 31126 3912 31178
rect 3912 31126 3928 31178
rect 3928 31126 3980 31178
rect 3980 31126 4290 31178
rect 5195 31158 5251 31214
rect 5276 31158 5332 31214
rect 5357 31158 5413 31214
rect 5438 31158 5494 31214
rect 5519 31158 5575 31214
rect 5600 31190 5632 31242
rect 5632 31190 5684 31242
rect 5684 31190 5700 31242
rect 5700 31190 5752 31242
rect 5752 31190 5768 31242
rect 5768 31190 5820 31242
rect 5820 31190 6376 31242
rect 5600 31178 6376 31190
rect 3514 31114 4290 31126
rect 3514 31062 3792 31114
rect 3792 31062 3844 31114
rect 3844 31062 3860 31114
rect 3860 31062 3912 31114
rect 3912 31062 3928 31114
rect 3928 31062 3980 31114
rect 3980 31062 4290 31114
rect 5195 31078 5251 31134
rect 5276 31078 5332 31134
rect 5357 31078 5413 31134
rect 5438 31078 5494 31134
rect 5519 31078 5575 31134
rect 5600 31126 5632 31178
rect 5632 31126 5684 31178
rect 5684 31126 5700 31178
rect 5700 31126 5752 31178
rect 5752 31126 5768 31178
rect 5768 31126 5820 31178
rect 5820 31126 6376 31178
rect 5600 31114 6376 31126
rect 5600 31062 5632 31114
rect 5632 31062 5684 31114
rect 5684 31062 5700 31114
rect 5700 31062 5752 31114
rect 5752 31062 5768 31114
rect 5768 31062 5820 31114
rect 5820 31062 6376 31114
rect 3109 30998 3165 31054
rect 3190 30998 3246 31054
rect 3271 30998 3327 31054
rect 3352 30998 3408 31054
rect 3433 30998 3489 31054
rect 3514 31050 4290 31062
rect 3514 30998 3792 31050
rect 3792 30998 3844 31050
rect 3844 30998 3860 31050
rect 3860 30998 3912 31050
rect 3912 30998 3928 31050
rect 3928 30998 3980 31050
rect 3980 30998 4290 31050
rect 5195 30998 5251 31054
rect 5276 30998 5332 31054
rect 5357 30998 5413 31054
rect 5438 30998 5494 31054
rect 5519 30998 5575 31054
rect 5600 31050 6376 31062
rect 5600 30998 5632 31050
rect 5632 30998 5684 31050
rect 5684 30998 5700 31050
rect 5700 30998 5752 31050
rect 5752 30998 5768 31050
rect 5768 30998 5820 31050
rect 5820 30998 6376 31050
rect 3514 30986 4290 30998
rect 5600 30986 6376 30998
rect 3109 30918 3165 30974
rect 3190 30918 3246 30974
rect 3271 30918 3327 30974
rect 3352 30918 3408 30974
rect 3433 30918 3489 30974
rect 3514 30934 3792 30986
rect 3792 30934 3844 30986
rect 3844 30934 3860 30986
rect 3860 30934 3912 30986
rect 3912 30934 3928 30986
rect 3928 30934 3980 30986
rect 3980 30934 4290 30986
rect 3514 30922 4290 30934
rect 3109 30838 3165 30894
rect 3190 30838 3246 30894
rect 3271 30838 3327 30894
rect 3352 30838 3408 30894
rect 3433 30838 3489 30894
rect 3514 30870 3792 30922
rect 3792 30870 3844 30922
rect 3844 30870 3860 30922
rect 3860 30870 3912 30922
rect 3912 30870 3928 30922
rect 3928 30870 3980 30922
rect 3980 30870 4290 30922
rect 5195 30918 5251 30974
rect 5276 30918 5332 30974
rect 5357 30918 5413 30974
rect 5438 30918 5494 30974
rect 5519 30918 5575 30974
rect 5600 30934 5632 30986
rect 5632 30934 5684 30986
rect 5684 30934 5700 30986
rect 5700 30934 5752 30986
rect 5752 30934 5768 30986
rect 5768 30934 5820 30986
rect 5820 30934 6376 30986
rect 5600 30922 6376 30934
rect 3514 30858 4290 30870
rect 3109 30758 3165 30814
rect 3190 30758 3246 30814
rect 3271 30758 3327 30814
rect 3352 30758 3408 30814
rect 3433 30758 3489 30814
rect 3514 30806 3792 30858
rect 3792 30806 3844 30858
rect 3844 30806 3860 30858
rect 3860 30806 3912 30858
rect 3912 30806 3928 30858
rect 3928 30806 3980 30858
rect 3980 30806 4290 30858
rect 5195 30838 5251 30894
rect 5276 30838 5332 30894
rect 5357 30838 5413 30894
rect 5438 30838 5494 30894
rect 5519 30838 5575 30894
rect 5600 30870 5632 30922
rect 5632 30870 5684 30922
rect 5684 30870 5700 30922
rect 5700 30870 5752 30922
rect 5752 30870 5768 30922
rect 5768 30870 5820 30922
rect 5820 30870 6376 30922
rect 5600 30858 6376 30870
rect 3514 30794 4290 30806
rect 3514 30742 3792 30794
rect 3792 30742 3844 30794
rect 3844 30742 3860 30794
rect 3860 30742 3912 30794
rect 3912 30742 3928 30794
rect 3928 30742 3980 30794
rect 3980 30742 4290 30794
rect 5195 30758 5251 30814
rect 5276 30758 5332 30814
rect 5357 30758 5413 30814
rect 5438 30758 5494 30814
rect 5519 30758 5575 30814
rect 5600 30806 5632 30858
rect 5632 30806 5684 30858
rect 5684 30806 5700 30858
rect 5700 30806 5752 30858
rect 5752 30806 5768 30858
rect 5768 30806 5820 30858
rect 5820 30806 6376 30858
rect 5600 30794 6376 30806
rect 5600 30742 5632 30794
rect 5632 30742 5684 30794
rect 5684 30742 5700 30794
rect 5700 30742 5752 30794
rect 5752 30742 5768 30794
rect 5768 30742 5820 30794
rect 5820 30742 6376 30794
rect 3109 30678 3165 30734
rect 3190 30678 3246 30734
rect 3271 30678 3327 30734
rect 3352 30678 3408 30734
rect 3433 30678 3489 30734
rect 3514 30729 4290 30742
rect 3514 30677 3792 30729
rect 3792 30677 3844 30729
rect 3844 30677 3860 30729
rect 3860 30677 3912 30729
rect 3912 30677 3928 30729
rect 3928 30677 3980 30729
rect 3980 30677 4290 30729
rect 5195 30678 5251 30734
rect 5276 30678 5332 30734
rect 5357 30678 5413 30734
rect 5438 30678 5494 30734
rect 5519 30678 5575 30734
rect 5600 30729 6376 30742
rect 5600 30677 5632 30729
rect 5632 30677 5684 30729
rect 5684 30677 5700 30729
rect 5700 30677 5752 30729
rect 5752 30677 5768 30729
rect 5768 30677 5820 30729
rect 5820 30677 6376 30729
rect 3514 30664 4290 30677
rect 5600 30664 6376 30677
rect 3109 30598 3165 30654
rect 3190 30598 3246 30654
rect 3271 30598 3327 30654
rect 3352 30598 3408 30654
rect 3433 30598 3489 30654
rect 3514 30612 3792 30664
rect 3792 30612 3844 30664
rect 3844 30612 3860 30664
rect 3860 30612 3912 30664
rect 3912 30612 3928 30664
rect 3928 30612 3980 30664
rect 3980 30612 4290 30664
rect 3514 30599 4290 30612
rect 3109 30518 3165 30574
rect 3190 30518 3246 30574
rect 3271 30518 3327 30574
rect 3352 30518 3408 30574
rect 3433 30518 3489 30574
rect 3514 30547 3792 30599
rect 3792 30547 3844 30599
rect 3844 30547 3860 30599
rect 3860 30547 3912 30599
rect 3912 30547 3928 30599
rect 3928 30547 3980 30599
rect 3980 30547 4290 30599
rect 5195 30598 5251 30654
rect 5276 30598 5332 30654
rect 5357 30598 5413 30654
rect 5438 30598 5494 30654
rect 5519 30598 5575 30654
rect 5600 30612 5632 30664
rect 5632 30612 5684 30664
rect 5684 30612 5700 30664
rect 5700 30612 5752 30664
rect 5752 30612 5768 30664
rect 5768 30612 5820 30664
rect 5820 30612 6376 30664
rect 5600 30599 6376 30612
rect 3514 30534 4290 30547
rect 3109 30438 3165 30494
rect 3190 30438 3246 30494
rect 3271 30438 3327 30494
rect 3352 30438 3408 30494
rect 3433 30438 3489 30494
rect 3514 30482 3792 30534
rect 3792 30482 3844 30534
rect 3844 30482 3860 30534
rect 3860 30482 3912 30534
rect 3912 30482 3928 30534
rect 3928 30482 3980 30534
rect 3980 30482 4290 30534
rect 5195 30518 5251 30574
rect 5276 30518 5332 30574
rect 5357 30518 5413 30574
rect 5438 30518 5494 30574
rect 5519 30518 5575 30574
rect 5600 30547 5632 30599
rect 5632 30547 5684 30599
rect 5684 30547 5700 30599
rect 5700 30547 5752 30599
rect 5752 30547 5768 30599
rect 5768 30547 5820 30599
rect 5820 30547 6376 30599
rect 5600 30534 6376 30547
rect 3514 30469 4290 30482
rect 3514 30417 3792 30469
rect 3792 30417 3844 30469
rect 3844 30417 3860 30469
rect 3860 30417 3912 30469
rect 3912 30417 3928 30469
rect 3928 30417 3980 30469
rect 3980 30417 4290 30469
rect 5195 30438 5251 30494
rect 5276 30438 5332 30494
rect 5357 30438 5413 30494
rect 5438 30438 5494 30494
rect 5519 30438 5575 30494
rect 5600 30482 5632 30534
rect 5632 30482 5684 30534
rect 5684 30482 5700 30534
rect 5700 30482 5752 30534
rect 5752 30482 5768 30534
rect 5768 30482 5820 30534
rect 5820 30482 6376 30534
rect 5600 30469 6376 30482
rect 5600 30417 5632 30469
rect 5632 30417 5684 30469
rect 5684 30417 5700 30469
rect 5700 30417 5752 30469
rect 5752 30417 5768 30469
rect 5768 30417 5820 30469
rect 5820 30417 6376 30469
rect 3109 30358 3165 30414
rect 3190 30358 3246 30414
rect 3271 30358 3327 30414
rect 3352 30358 3408 30414
rect 3433 30358 3489 30414
rect 3514 30404 4290 30417
rect 3514 30352 3792 30404
rect 3792 30352 3844 30404
rect 3844 30352 3860 30404
rect 3860 30352 3912 30404
rect 3912 30352 3928 30404
rect 3928 30352 3980 30404
rect 3980 30352 4290 30404
rect 5195 30358 5251 30414
rect 5276 30358 5332 30414
rect 5357 30358 5413 30414
rect 5438 30358 5494 30414
rect 5519 30358 5575 30414
rect 5600 30404 6376 30417
rect 5600 30352 5632 30404
rect 5632 30352 5684 30404
rect 5684 30352 5700 30404
rect 5700 30352 5752 30404
rect 5752 30352 5768 30404
rect 5768 30352 5820 30404
rect 5820 30352 6376 30404
rect 3514 30339 4290 30352
rect 5600 30339 6376 30352
rect 3109 30278 3165 30334
rect 3190 30278 3246 30334
rect 3271 30278 3327 30334
rect 3352 30278 3408 30334
rect 3433 30278 3489 30334
rect 3514 30287 3792 30339
rect 3792 30287 3844 30339
rect 3844 30287 3860 30339
rect 3860 30287 3912 30339
rect 3912 30287 3928 30339
rect 3928 30287 3980 30339
rect 3980 30287 4290 30339
rect 3514 30274 4290 30287
rect 5195 30278 5251 30334
rect 5276 30278 5332 30334
rect 5357 30278 5413 30334
rect 5438 30278 5494 30334
rect 5519 30278 5575 30334
rect 5600 30287 5632 30339
rect 5632 30287 5684 30339
rect 5684 30287 5700 30339
rect 5700 30287 5752 30339
rect 5752 30287 5768 30339
rect 5768 30287 5820 30339
rect 5820 30287 6376 30339
rect 5600 30274 6376 30287
rect 3109 30198 3165 30254
rect 3190 30198 3246 30254
rect 3271 30198 3327 30254
rect 3352 30198 3408 30254
rect 3433 30198 3489 30254
rect 3514 30222 3792 30274
rect 3792 30222 3844 30274
rect 3844 30222 3860 30274
rect 3860 30222 3912 30274
rect 3912 30222 3928 30274
rect 3928 30222 3980 30274
rect 3980 30222 4290 30274
rect 3514 30209 4290 30222
rect 3109 30118 3165 30174
rect 3190 30118 3246 30174
rect 3271 30118 3327 30174
rect 3352 30118 3408 30174
rect 3433 30118 3489 30174
rect 3514 30157 3792 30209
rect 3792 30157 3844 30209
rect 3844 30157 3860 30209
rect 3860 30157 3912 30209
rect 3912 30157 3928 30209
rect 3928 30157 3980 30209
rect 3980 30157 4290 30209
rect 5195 30198 5251 30254
rect 5276 30198 5332 30254
rect 5357 30198 5413 30254
rect 5438 30198 5494 30254
rect 5519 30198 5575 30254
rect 5600 30222 5632 30274
rect 5632 30222 5684 30274
rect 5684 30222 5700 30274
rect 5700 30222 5752 30274
rect 5752 30222 5768 30274
rect 5768 30222 5820 30274
rect 5820 30222 6376 30274
rect 5600 30209 6376 30222
rect 3514 30144 4290 30157
rect 3109 30038 3165 30094
rect 3190 30038 3246 30094
rect 3271 30038 3327 30094
rect 3352 30038 3408 30094
rect 3433 30038 3489 30094
rect 3514 30092 3792 30144
rect 3792 30092 3844 30144
rect 3844 30092 3860 30144
rect 3860 30092 3912 30144
rect 3912 30092 3928 30144
rect 3928 30092 3980 30144
rect 3980 30092 4290 30144
rect 5195 30118 5251 30174
rect 5276 30118 5332 30174
rect 5357 30118 5413 30174
rect 5438 30118 5494 30174
rect 5519 30118 5575 30174
rect 5600 30157 5632 30209
rect 5632 30157 5684 30209
rect 5684 30157 5700 30209
rect 5700 30157 5752 30209
rect 5752 30157 5768 30209
rect 5768 30157 5820 30209
rect 5820 30157 6376 30209
rect 5600 30144 6376 30157
rect 3514 30079 4290 30092
rect 3514 30027 3792 30079
rect 3792 30027 3844 30079
rect 3844 30027 3860 30079
rect 3860 30027 3912 30079
rect 3912 30027 3928 30079
rect 3928 30027 3980 30079
rect 3980 30027 4290 30079
rect 5195 30038 5251 30094
rect 5276 30038 5332 30094
rect 5357 30038 5413 30094
rect 5438 30038 5494 30094
rect 5519 30038 5575 30094
rect 5600 30092 5632 30144
rect 5632 30092 5684 30144
rect 5684 30092 5700 30144
rect 5700 30092 5752 30144
rect 5752 30092 5768 30144
rect 5768 30092 5820 30144
rect 5820 30092 6376 30144
rect 5600 30079 6376 30092
rect 5600 30027 5632 30079
rect 5632 30027 5684 30079
rect 5684 30027 5700 30079
rect 5700 30027 5752 30079
rect 5752 30027 5768 30079
rect 5768 30027 5820 30079
rect 5820 30027 6376 30079
rect 3514 30014 4290 30027
rect 5600 30014 6376 30027
rect 3109 29958 3165 30014
rect 3190 29958 3246 30014
rect 3271 29958 3327 30014
rect 3352 29958 3408 30014
rect 3433 29958 3489 30014
rect 3514 29962 3792 30014
rect 3792 29962 3844 30014
rect 3844 29962 3860 30014
rect 3860 29962 3912 30014
rect 3912 29962 3928 30014
rect 3928 29962 3980 30014
rect 3980 29962 4290 30014
rect 3514 29958 4290 29962
rect 5195 29958 5251 30014
rect 5276 29958 5332 30014
rect 5357 29958 5413 30014
rect 5438 29958 5494 30014
rect 5519 29958 5575 30014
rect 5600 29962 5632 30014
rect 5632 29962 5684 30014
rect 5684 29962 5700 30014
rect 5700 29962 5752 30014
rect 5752 29962 5768 30014
rect 5768 29962 5820 30014
rect 5820 29962 6376 30014
rect 5600 29958 6376 29962
rect 8580 29573 8636 29629
rect 8661 29573 8717 29629
rect 8742 29573 8798 29629
rect 8823 29573 8879 29629
rect 8904 29625 8960 29629
rect 8985 29625 9041 29629
rect 8904 29573 8933 29625
rect 8933 29573 8959 29625
rect 8959 29573 8960 29625
rect 8985 29573 9011 29625
rect 9011 29573 9041 29625
rect 8580 29493 8636 29549
rect 8661 29493 8717 29549
rect 8742 29493 8798 29549
rect 8823 29493 8879 29549
rect 8904 29509 8933 29549
rect 8933 29509 8959 29549
rect 8959 29509 8960 29549
rect 8985 29509 9011 29549
rect 9011 29509 9041 29549
rect 8904 29497 8960 29509
rect 8985 29497 9041 29509
rect 8904 29493 8933 29497
rect 8933 29493 8959 29497
rect 8959 29493 8960 29497
rect 8985 29493 9011 29497
rect 9011 29493 9041 29497
rect 8580 29413 8636 29469
rect 8661 29413 8717 29469
rect 8742 29413 8798 29469
rect 8823 29413 8879 29469
rect 8904 29445 8933 29469
rect 8933 29445 8959 29469
rect 8959 29445 8960 29469
rect 8985 29445 9011 29469
rect 9011 29445 9041 29469
rect 8904 29433 8960 29445
rect 8985 29433 9041 29445
rect 8904 29413 8933 29433
rect 8933 29413 8959 29433
rect 8959 29413 8960 29433
rect 8985 29413 9011 29433
rect 9011 29413 9041 29433
rect 8580 29333 8636 29389
rect 8661 29333 8717 29389
rect 8742 29333 8798 29389
rect 8823 29333 8879 29389
rect 8904 29381 8933 29389
rect 8933 29381 8959 29389
rect 8959 29381 8960 29389
rect 8985 29381 9011 29389
rect 9011 29381 9041 29389
rect 8904 29369 8960 29381
rect 8985 29369 9041 29381
rect 8904 29333 8933 29369
rect 8933 29333 8959 29369
rect 8959 29333 8960 29369
rect 8985 29333 9011 29369
rect 9011 29333 9041 29369
rect 8580 29253 8636 29309
rect 8661 29253 8717 29309
rect 8742 29253 8798 29309
rect 8823 29253 8879 29309
rect 8904 29305 8960 29309
rect 8985 29305 9041 29309
rect 8904 29253 8933 29305
rect 8933 29253 8959 29305
rect 8959 29253 8960 29305
rect 8985 29253 9011 29305
rect 9011 29253 9041 29305
rect 8580 29173 8636 29229
rect 8661 29173 8717 29229
rect 8742 29173 8798 29229
rect 8823 29173 8879 29229
rect 8904 29189 8933 29229
rect 8933 29189 8959 29229
rect 8959 29189 8960 29229
rect 8985 29189 9011 29229
rect 9011 29189 9041 29229
rect 8904 29177 8960 29189
rect 8985 29177 9041 29189
rect 8904 29173 8933 29177
rect 8933 29173 8959 29177
rect 8959 29173 8960 29177
rect 8985 29173 9011 29177
rect 9011 29173 9041 29177
rect 8580 29093 8636 29149
rect 8661 29093 8717 29149
rect 8742 29093 8798 29149
rect 8823 29093 8879 29149
rect 8904 29125 8933 29149
rect 8933 29125 8959 29149
rect 8959 29125 8960 29149
rect 8985 29125 9011 29149
rect 9011 29125 9041 29149
rect 8904 29113 8960 29125
rect 8985 29113 9041 29125
rect 8904 29093 8933 29113
rect 8933 29093 8959 29113
rect 8959 29093 8960 29113
rect 8985 29093 9011 29113
rect 9011 29093 9041 29113
rect 8580 29013 8636 29069
rect 8661 29013 8717 29069
rect 8742 29013 8798 29069
rect 8823 29013 8879 29069
rect 8904 29061 8933 29069
rect 8933 29061 8959 29069
rect 8959 29061 8960 29069
rect 8985 29061 9011 29069
rect 9011 29061 9041 29069
rect 8904 29049 8960 29061
rect 8985 29049 9041 29061
rect 8904 29013 8933 29049
rect 8933 29013 8959 29049
rect 8959 29013 8960 29049
rect 8985 29013 9011 29049
rect 9011 29013 9041 29049
rect 8580 28933 8636 28989
rect 8661 28933 8717 28989
rect 8742 28933 8798 28989
rect 8823 28933 8879 28989
rect 8904 28985 8960 28989
rect 8985 28985 9041 28989
rect 8904 28933 8933 28985
rect 8933 28933 8959 28985
rect 8959 28933 8960 28985
rect 8985 28933 9011 28985
rect 9011 28933 9041 28985
rect 8580 28853 8636 28909
rect 8661 28853 8717 28909
rect 8742 28853 8798 28909
rect 8823 28853 8879 28909
rect 8904 28869 8933 28909
rect 8933 28869 8959 28909
rect 8959 28869 8960 28909
rect 8985 28869 9011 28909
rect 9011 28869 9041 28909
rect 8904 28857 8960 28869
rect 8985 28857 9041 28869
rect 8904 28853 8933 28857
rect 8933 28853 8959 28857
rect 8959 28853 8960 28857
rect 8985 28853 9011 28857
rect 9011 28853 9041 28857
rect 8580 28773 8636 28829
rect 8661 28773 8717 28829
rect 8742 28773 8798 28829
rect 8823 28773 8879 28829
rect 8904 28805 8933 28829
rect 8933 28805 8959 28829
rect 8959 28805 8960 28829
rect 8985 28805 9011 28829
rect 9011 28805 9041 28829
rect 8904 28793 8960 28805
rect 8985 28793 9041 28805
rect 8904 28773 8933 28793
rect 8933 28773 8959 28793
rect 8959 28773 8960 28793
rect 8985 28773 9011 28793
rect 9011 28773 9041 28793
rect 8580 28693 8636 28749
rect 8661 28693 8717 28749
rect 8742 28693 8798 28749
rect 8823 28693 8879 28749
rect 8904 28741 8933 28749
rect 8933 28741 8959 28749
rect 8959 28741 8960 28749
rect 8985 28741 9011 28749
rect 9011 28741 9041 28749
rect 8904 28729 8960 28741
rect 8985 28729 9041 28741
rect 8904 28693 8933 28729
rect 8933 28693 8959 28729
rect 8959 28693 8960 28729
rect 8985 28693 9011 28729
rect 9011 28693 9041 28729
rect 8580 28613 8636 28669
rect 8661 28613 8717 28669
rect 8742 28613 8798 28669
rect 8823 28613 8879 28669
rect 8904 28664 8960 28669
rect 8985 28664 9041 28669
rect 8904 28613 8933 28664
rect 8933 28613 8959 28664
rect 8959 28613 8960 28664
rect 8985 28613 9011 28664
rect 9011 28613 9041 28664
rect 8580 28533 8636 28589
rect 8661 28533 8717 28589
rect 8742 28533 8798 28589
rect 8823 28533 8879 28589
rect 8904 28547 8933 28589
rect 8933 28547 8959 28589
rect 8959 28547 8960 28589
rect 8985 28547 9011 28589
rect 9011 28547 9041 28589
rect 8904 28534 8960 28547
rect 8985 28534 9041 28547
rect 8904 28533 8933 28534
rect 8933 28533 8959 28534
rect 8959 28533 8960 28534
rect 8985 28533 9011 28534
rect 9011 28533 9041 28534
rect 8580 28453 8636 28509
rect 8661 28453 8717 28509
rect 8742 28453 8798 28509
rect 8823 28453 8879 28509
rect 8904 28482 8933 28509
rect 8933 28482 8959 28509
rect 8959 28482 8960 28509
rect 8985 28482 9011 28509
rect 9011 28482 9041 28509
rect 8904 28469 8960 28482
rect 8985 28469 9041 28482
rect 8904 28453 8933 28469
rect 8933 28453 8959 28469
rect 8959 28453 8960 28469
rect 8985 28453 9011 28469
rect 9011 28453 9041 28469
rect 8580 28373 8636 28429
rect 8661 28373 8717 28429
rect 8742 28373 8798 28429
rect 8823 28373 8879 28429
rect 8904 28417 8933 28429
rect 8933 28417 8959 28429
rect 8959 28417 8960 28429
rect 8985 28417 9011 28429
rect 9011 28417 9041 28429
rect 8904 28404 8960 28417
rect 8985 28404 9041 28417
rect 8904 28373 8933 28404
rect 8933 28373 8959 28404
rect 8959 28373 8960 28404
rect 8985 28373 9011 28404
rect 9011 28373 9041 28404
rect 8580 28293 8636 28349
rect 8661 28293 8717 28349
rect 8742 28293 8798 28349
rect 8823 28293 8879 28349
rect 8904 28339 8960 28349
rect 8985 28339 9041 28349
rect 8904 28293 8933 28339
rect 8933 28293 8959 28339
rect 8959 28293 8960 28339
rect 8985 28293 9011 28339
rect 9011 28293 9041 28339
rect 8580 28213 8636 28269
rect 8661 28213 8717 28269
rect 8742 28213 8798 28269
rect 8823 28213 8879 28269
rect 8904 28222 8933 28269
rect 8933 28222 8959 28269
rect 8959 28222 8960 28269
rect 8985 28222 9011 28269
rect 9011 28222 9041 28269
rect 8904 28213 8960 28222
rect 8985 28213 9041 28222
rect 8580 28133 8636 28189
rect 8661 28133 8717 28189
rect 8742 28133 8798 28189
rect 8823 28133 8879 28189
rect 8904 28157 8933 28189
rect 8933 28157 8959 28189
rect 8959 28157 8960 28189
rect 8985 28157 9011 28189
rect 9011 28157 9041 28189
rect 8904 28144 8960 28157
rect 8985 28144 9041 28157
rect 8904 28133 8933 28144
rect 8933 28133 8959 28144
rect 8959 28133 8960 28144
rect 8985 28133 9011 28144
rect 9011 28133 9041 28144
rect 8580 28053 8636 28109
rect 8661 28053 8717 28109
rect 8742 28053 8798 28109
rect 8823 28053 8879 28109
rect 8904 28092 8933 28109
rect 8933 28092 8959 28109
rect 8959 28092 8960 28109
rect 8985 28092 9011 28109
rect 9011 28092 9041 28109
rect 8904 28079 8960 28092
rect 8985 28079 9041 28092
rect 8904 28053 8933 28079
rect 8933 28053 8959 28079
rect 8959 28053 8960 28079
rect 8985 28053 9011 28079
rect 9011 28053 9041 28079
rect 8580 27973 8636 28029
rect 8661 27973 8717 28029
rect 8742 27973 8798 28029
rect 8823 27973 8879 28029
rect 8904 28027 8933 28029
rect 8933 28027 8959 28029
rect 8959 28027 8960 28029
rect 8985 28027 9011 28029
rect 9011 28027 9041 28029
rect 8904 28014 8960 28027
rect 8985 28014 9041 28027
rect 8904 27973 8933 28014
rect 8933 27973 8959 28014
rect 8959 27973 8960 28014
rect 8985 27973 9011 28014
rect 9011 27973 9041 28014
rect 8580 27893 8636 27949
rect 8661 27893 8717 27949
rect 8742 27893 8798 27949
rect 8823 27893 8879 27949
rect 8904 27897 8933 27949
rect 8933 27897 8959 27949
rect 8959 27897 8960 27949
rect 8985 27897 9011 27949
rect 9011 27897 9041 27949
rect 8904 27893 8960 27897
rect 8985 27893 9041 27897
rect 9066 27893 9762 29629
rect 10666 29625 10722 29629
rect 10747 29625 10803 29629
rect 10828 29625 10884 29629
rect 10666 29573 10721 29625
rect 10721 29573 10722 29625
rect 10747 29573 10773 29625
rect 10773 29573 10799 29625
rect 10799 29573 10803 29625
rect 10828 29573 10851 29625
rect 10851 29573 10884 29625
rect 10909 29573 10965 29629
rect 10990 29573 11046 29629
rect 11071 29573 11127 29629
rect 11152 29625 11848 29629
rect 11152 29573 11641 29625
rect 11641 29573 11693 29625
rect 11693 29573 11719 29625
rect 11719 29573 11771 29625
rect 11771 29573 11848 29625
rect 11152 29561 11848 29573
rect 10666 29509 10721 29549
rect 10721 29509 10722 29549
rect 10747 29509 10773 29549
rect 10773 29509 10799 29549
rect 10799 29509 10803 29549
rect 10828 29509 10851 29549
rect 10851 29509 10884 29549
rect 10666 29497 10722 29509
rect 10747 29497 10803 29509
rect 10828 29497 10884 29509
rect 10666 29493 10721 29497
rect 10721 29493 10722 29497
rect 10747 29493 10773 29497
rect 10773 29493 10799 29497
rect 10799 29493 10803 29497
rect 10828 29493 10851 29497
rect 10851 29493 10884 29497
rect 10909 29493 10965 29549
rect 10990 29493 11046 29549
rect 11071 29493 11127 29549
rect 11152 29509 11641 29561
rect 11641 29509 11693 29561
rect 11693 29509 11719 29561
rect 11719 29509 11771 29561
rect 11771 29509 11848 29561
rect 11152 29497 11848 29509
rect 10666 29445 10721 29469
rect 10721 29445 10722 29469
rect 10747 29445 10773 29469
rect 10773 29445 10799 29469
rect 10799 29445 10803 29469
rect 10828 29445 10851 29469
rect 10851 29445 10884 29469
rect 10666 29433 10722 29445
rect 10747 29433 10803 29445
rect 10828 29433 10884 29445
rect 10666 29413 10721 29433
rect 10721 29413 10722 29433
rect 10747 29413 10773 29433
rect 10773 29413 10799 29433
rect 10799 29413 10803 29433
rect 10828 29413 10851 29433
rect 10851 29413 10884 29433
rect 10909 29413 10965 29469
rect 10990 29413 11046 29469
rect 11071 29413 11127 29469
rect 11152 29445 11641 29497
rect 11641 29445 11693 29497
rect 11693 29445 11719 29497
rect 11719 29445 11771 29497
rect 11771 29445 11848 29497
rect 11152 29433 11848 29445
rect 10666 29381 10721 29389
rect 10721 29381 10722 29389
rect 10747 29381 10773 29389
rect 10773 29381 10799 29389
rect 10799 29381 10803 29389
rect 10828 29381 10851 29389
rect 10851 29381 10884 29389
rect 10666 29369 10722 29381
rect 10747 29369 10803 29381
rect 10828 29369 10884 29381
rect 10666 29333 10721 29369
rect 10721 29333 10722 29369
rect 10747 29333 10773 29369
rect 10773 29333 10799 29369
rect 10799 29333 10803 29369
rect 10828 29333 10851 29369
rect 10851 29333 10884 29369
rect 10909 29333 10965 29389
rect 10990 29333 11046 29389
rect 11071 29333 11127 29389
rect 11152 29381 11641 29433
rect 11641 29381 11693 29433
rect 11693 29381 11719 29433
rect 11719 29381 11771 29433
rect 11771 29381 11848 29433
rect 11152 29369 11848 29381
rect 11152 29317 11641 29369
rect 11641 29317 11693 29369
rect 11693 29317 11719 29369
rect 11719 29317 11771 29369
rect 11771 29317 11848 29369
rect 10666 29305 10722 29309
rect 10747 29305 10803 29309
rect 10828 29305 10884 29309
rect 10666 29253 10721 29305
rect 10721 29253 10722 29305
rect 10747 29253 10773 29305
rect 10773 29253 10799 29305
rect 10799 29253 10803 29305
rect 10828 29253 10851 29305
rect 10851 29253 10884 29305
rect 10909 29253 10965 29309
rect 10990 29253 11046 29309
rect 11071 29253 11127 29309
rect 11152 29305 11848 29317
rect 11152 29253 11641 29305
rect 11641 29253 11693 29305
rect 11693 29253 11719 29305
rect 11719 29253 11771 29305
rect 11771 29253 11848 29305
rect 11152 29241 11848 29253
rect 10666 29189 10721 29229
rect 10721 29189 10722 29229
rect 10747 29189 10773 29229
rect 10773 29189 10799 29229
rect 10799 29189 10803 29229
rect 10828 29189 10851 29229
rect 10851 29189 10884 29229
rect 10666 29177 10722 29189
rect 10747 29177 10803 29189
rect 10828 29177 10884 29189
rect 10666 29173 10721 29177
rect 10721 29173 10722 29177
rect 10747 29173 10773 29177
rect 10773 29173 10799 29177
rect 10799 29173 10803 29177
rect 10828 29173 10851 29177
rect 10851 29173 10884 29177
rect 10909 29173 10965 29229
rect 10990 29173 11046 29229
rect 11071 29173 11127 29229
rect 11152 29189 11641 29241
rect 11641 29189 11693 29241
rect 11693 29189 11719 29241
rect 11719 29189 11771 29241
rect 11771 29189 11848 29241
rect 11152 29177 11848 29189
rect 10666 29125 10721 29149
rect 10721 29125 10722 29149
rect 10747 29125 10773 29149
rect 10773 29125 10799 29149
rect 10799 29125 10803 29149
rect 10828 29125 10851 29149
rect 10851 29125 10884 29149
rect 10666 29113 10722 29125
rect 10747 29113 10803 29125
rect 10828 29113 10884 29125
rect 10666 29093 10721 29113
rect 10721 29093 10722 29113
rect 10747 29093 10773 29113
rect 10773 29093 10799 29113
rect 10799 29093 10803 29113
rect 10828 29093 10851 29113
rect 10851 29093 10884 29113
rect 10909 29093 10965 29149
rect 10990 29093 11046 29149
rect 11071 29093 11127 29149
rect 11152 29125 11641 29177
rect 11641 29125 11693 29177
rect 11693 29125 11719 29177
rect 11719 29125 11771 29177
rect 11771 29125 11848 29177
rect 11152 29113 11848 29125
rect 10666 29061 10721 29069
rect 10721 29061 10722 29069
rect 10747 29061 10773 29069
rect 10773 29061 10799 29069
rect 10799 29061 10803 29069
rect 10828 29061 10851 29069
rect 10851 29061 10884 29069
rect 10666 29049 10722 29061
rect 10747 29049 10803 29061
rect 10828 29049 10884 29061
rect 10666 29013 10721 29049
rect 10721 29013 10722 29049
rect 10747 29013 10773 29049
rect 10773 29013 10799 29049
rect 10799 29013 10803 29049
rect 10828 29013 10851 29049
rect 10851 29013 10884 29049
rect 10909 29013 10965 29069
rect 10990 29013 11046 29069
rect 11071 29013 11127 29069
rect 11152 29061 11641 29113
rect 11641 29061 11693 29113
rect 11693 29061 11719 29113
rect 11719 29061 11771 29113
rect 11771 29061 11848 29113
rect 11152 29049 11848 29061
rect 11152 28997 11641 29049
rect 11641 28997 11693 29049
rect 11693 28997 11719 29049
rect 11719 28997 11771 29049
rect 11771 28997 11848 29049
rect 10666 28985 10722 28989
rect 10747 28985 10803 28989
rect 10828 28985 10884 28989
rect 10666 28933 10721 28985
rect 10721 28933 10722 28985
rect 10747 28933 10773 28985
rect 10773 28933 10799 28985
rect 10799 28933 10803 28985
rect 10828 28933 10851 28985
rect 10851 28933 10884 28985
rect 10909 28933 10965 28989
rect 10990 28933 11046 28989
rect 11071 28933 11127 28989
rect 11152 28985 11848 28997
rect 11152 28933 11641 28985
rect 11641 28933 11693 28985
rect 11693 28933 11719 28985
rect 11719 28933 11771 28985
rect 11771 28933 11848 28985
rect 11152 28921 11848 28933
rect 10666 28869 10721 28909
rect 10721 28869 10722 28909
rect 10747 28869 10773 28909
rect 10773 28869 10799 28909
rect 10799 28869 10803 28909
rect 10828 28869 10851 28909
rect 10851 28869 10884 28909
rect 10666 28857 10722 28869
rect 10747 28857 10803 28869
rect 10828 28857 10884 28869
rect 10666 28853 10721 28857
rect 10721 28853 10722 28857
rect 10747 28853 10773 28857
rect 10773 28853 10799 28857
rect 10799 28853 10803 28857
rect 10828 28853 10851 28857
rect 10851 28853 10884 28857
rect 10909 28853 10965 28909
rect 10990 28853 11046 28909
rect 11071 28853 11127 28909
rect 11152 28869 11641 28921
rect 11641 28869 11693 28921
rect 11693 28869 11719 28921
rect 11719 28869 11771 28921
rect 11771 28869 11848 28921
rect 11152 28857 11848 28869
rect 10666 28805 10721 28829
rect 10721 28805 10722 28829
rect 10747 28805 10773 28829
rect 10773 28805 10799 28829
rect 10799 28805 10803 28829
rect 10828 28805 10851 28829
rect 10851 28805 10884 28829
rect 10666 28793 10722 28805
rect 10747 28793 10803 28805
rect 10828 28793 10884 28805
rect 10666 28773 10721 28793
rect 10721 28773 10722 28793
rect 10747 28773 10773 28793
rect 10773 28773 10799 28793
rect 10799 28773 10803 28793
rect 10828 28773 10851 28793
rect 10851 28773 10884 28793
rect 10909 28773 10965 28829
rect 10990 28773 11046 28829
rect 11071 28773 11127 28829
rect 11152 28805 11641 28857
rect 11641 28805 11693 28857
rect 11693 28805 11719 28857
rect 11719 28805 11771 28857
rect 11771 28805 11848 28857
rect 11152 28793 11848 28805
rect 10666 28741 10721 28749
rect 10721 28741 10722 28749
rect 10747 28741 10773 28749
rect 10773 28741 10799 28749
rect 10799 28741 10803 28749
rect 10828 28741 10851 28749
rect 10851 28741 10884 28749
rect 10666 28729 10722 28741
rect 10747 28729 10803 28741
rect 10828 28729 10884 28741
rect 10666 28693 10721 28729
rect 10721 28693 10722 28729
rect 10747 28693 10773 28729
rect 10773 28693 10799 28729
rect 10799 28693 10803 28729
rect 10828 28693 10851 28729
rect 10851 28693 10884 28729
rect 10909 28693 10965 28749
rect 10990 28693 11046 28749
rect 11071 28693 11127 28749
rect 11152 28741 11641 28793
rect 11641 28741 11693 28793
rect 11693 28741 11719 28793
rect 11719 28741 11771 28793
rect 11771 28741 11848 28793
rect 11152 28729 11848 28741
rect 11152 28677 11641 28729
rect 11641 28677 11693 28729
rect 11693 28677 11719 28729
rect 11719 28677 11771 28729
rect 11771 28677 11848 28729
rect 10666 28664 10722 28669
rect 10747 28664 10803 28669
rect 10828 28664 10884 28669
rect 10666 28613 10721 28664
rect 10721 28613 10722 28664
rect 10747 28613 10773 28664
rect 10773 28613 10799 28664
rect 10799 28613 10803 28664
rect 10828 28613 10851 28664
rect 10851 28613 10884 28664
rect 10909 28613 10965 28669
rect 10990 28613 11046 28669
rect 11071 28613 11127 28669
rect 11152 28664 11848 28677
rect 11152 28612 11641 28664
rect 11641 28612 11693 28664
rect 11693 28612 11719 28664
rect 11719 28612 11771 28664
rect 11771 28612 11848 28664
rect 11152 28599 11848 28612
rect 10666 28547 10721 28589
rect 10721 28547 10722 28589
rect 10747 28547 10773 28589
rect 10773 28547 10799 28589
rect 10799 28547 10803 28589
rect 10828 28547 10851 28589
rect 10851 28547 10884 28589
rect 10666 28534 10722 28547
rect 10747 28534 10803 28547
rect 10828 28534 10884 28547
rect 10666 28533 10721 28534
rect 10721 28533 10722 28534
rect 10747 28533 10773 28534
rect 10773 28533 10799 28534
rect 10799 28533 10803 28534
rect 10828 28533 10851 28534
rect 10851 28533 10884 28534
rect 10909 28533 10965 28589
rect 10990 28533 11046 28589
rect 11071 28533 11127 28589
rect 11152 28547 11641 28599
rect 11641 28547 11693 28599
rect 11693 28547 11719 28599
rect 11719 28547 11771 28599
rect 11771 28547 11848 28599
rect 11152 28534 11848 28547
rect 10666 28482 10721 28509
rect 10721 28482 10722 28509
rect 10747 28482 10773 28509
rect 10773 28482 10799 28509
rect 10799 28482 10803 28509
rect 10828 28482 10851 28509
rect 10851 28482 10884 28509
rect 10666 28469 10722 28482
rect 10747 28469 10803 28482
rect 10828 28469 10884 28482
rect 10666 28453 10721 28469
rect 10721 28453 10722 28469
rect 10747 28453 10773 28469
rect 10773 28453 10799 28469
rect 10799 28453 10803 28469
rect 10828 28453 10851 28469
rect 10851 28453 10884 28469
rect 10909 28453 10965 28509
rect 10990 28453 11046 28509
rect 11071 28453 11127 28509
rect 11152 28482 11641 28534
rect 11641 28482 11693 28534
rect 11693 28482 11719 28534
rect 11719 28482 11771 28534
rect 11771 28482 11848 28534
rect 11152 28469 11848 28482
rect 10666 28417 10721 28429
rect 10721 28417 10722 28429
rect 10747 28417 10773 28429
rect 10773 28417 10799 28429
rect 10799 28417 10803 28429
rect 10828 28417 10851 28429
rect 10851 28417 10884 28429
rect 10666 28404 10722 28417
rect 10747 28404 10803 28417
rect 10828 28404 10884 28417
rect 10666 28373 10721 28404
rect 10721 28373 10722 28404
rect 10747 28373 10773 28404
rect 10773 28373 10799 28404
rect 10799 28373 10803 28404
rect 10828 28373 10851 28404
rect 10851 28373 10884 28404
rect 10909 28373 10965 28429
rect 10990 28373 11046 28429
rect 11071 28373 11127 28429
rect 11152 28417 11641 28469
rect 11641 28417 11693 28469
rect 11693 28417 11719 28469
rect 11719 28417 11771 28469
rect 11771 28417 11848 28469
rect 11152 28404 11848 28417
rect 11152 28352 11641 28404
rect 11641 28352 11693 28404
rect 11693 28352 11719 28404
rect 11719 28352 11771 28404
rect 11771 28352 11848 28404
rect 10666 28339 10722 28349
rect 10747 28339 10803 28349
rect 10828 28339 10884 28349
rect 10666 28293 10721 28339
rect 10721 28293 10722 28339
rect 10747 28293 10773 28339
rect 10773 28293 10799 28339
rect 10799 28293 10803 28339
rect 10828 28293 10851 28339
rect 10851 28293 10884 28339
rect 10909 28293 10965 28349
rect 10990 28293 11046 28349
rect 11071 28293 11127 28349
rect 11152 28339 11848 28352
rect 11152 28287 11641 28339
rect 11641 28287 11693 28339
rect 11693 28287 11719 28339
rect 11719 28287 11771 28339
rect 11771 28287 11848 28339
rect 11152 28274 11848 28287
rect 10666 28222 10721 28269
rect 10721 28222 10722 28269
rect 10747 28222 10773 28269
rect 10773 28222 10799 28269
rect 10799 28222 10803 28269
rect 10828 28222 10851 28269
rect 10851 28222 10884 28269
rect 10666 28213 10722 28222
rect 10747 28213 10803 28222
rect 10828 28213 10884 28222
rect 10909 28213 10965 28269
rect 10990 28213 11046 28269
rect 11071 28213 11127 28269
rect 11152 28222 11641 28274
rect 11641 28222 11693 28274
rect 11693 28222 11719 28274
rect 11719 28222 11771 28274
rect 11771 28222 11848 28274
rect 11152 28209 11848 28222
rect 10666 28157 10721 28189
rect 10721 28157 10722 28189
rect 10747 28157 10773 28189
rect 10773 28157 10799 28189
rect 10799 28157 10803 28189
rect 10828 28157 10851 28189
rect 10851 28157 10884 28189
rect 10666 28144 10722 28157
rect 10747 28144 10803 28157
rect 10828 28144 10884 28157
rect 10666 28133 10721 28144
rect 10721 28133 10722 28144
rect 10747 28133 10773 28144
rect 10773 28133 10799 28144
rect 10799 28133 10803 28144
rect 10828 28133 10851 28144
rect 10851 28133 10884 28144
rect 10909 28133 10965 28189
rect 10990 28133 11046 28189
rect 11071 28133 11127 28189
rect 11152 28157 11641 28209
rect 11641 28157 11693 28209
rect 11693 28157 11719 28209
rect 11719 28157 11771 28209
rect 11771 28157 11848 28209
rect 11152 28144 11848 28157
rect 10666 28092 10721 28109
rect 10721 28092 10722 28109
rect 10747 28092 10773 28109
rect 10773 28092 10799 28109
rect 10799 28092 10803 28109
rect 10828 28092 10851 28109
rect 10851 28092 10884 28109
rect 10666 28079 10722 28092
rect 10747 28079 10803 28092
rect 10828 28079 10884 28092
rect 10666 28053 10721 28079
rect 10721 28053 10722 28079
rect 10747 28053 10773 28079
rect 10773 28053 10799 28079
rect 10799 28053 10803 28079
rect 10828 28053 10851 28079
rect 10851 28053 10884 28079
rect 10909 28053 10965 28109
rect 10990 28053 11046 28109
rect 11071 28053 11127 28109
rect 11152 28092 11641 28144
rect 11641 28092 11693 28144
rect 11693 28092 11719 28144
rect 11719 28092 11771 28144
rect 11771 28092 11848 28144
rect 11152 28079 11848 28092
rect 10666 28027 10721 28029
rect 10721 28027 10722 28029
rect 10747 28027 10773 28029
rect 10773 28027 10799 28029
rect 10799 28027 10803 28029
rect 10828 28027 10851 28029
rect 10851 28027 10884 28029
rect 10666 28014 10722 28027
rect 10747 28014 10803 28027
rect 10828 28014 10884 28027
rect 10666 27973 10721 28014
rect 10721 27973 10722 28014
rect 10747 27973 10773 28014
rect 10773 27973 10799 28014
rect 10799 27973 10803 28014
rect 10828 27973 10851 28014
rect 10851 27973 10884 28014
rect 10909 27973 10965 28029
rect 10990 27973 11046 28029
rect 11071 27973 11127 28029
rect 11152 28027 11641 28079
rect 11641 28027 11693 28079
rect 11693 28027 11719 28079
rect 11719 28027 11771 28079
rect 11771 28027 11848 28079
rect 11152 28014 11848 28027
rect 11152 27962 11641 28014
rect 11641 27962 11693 28014
rect 11693 27962 11719 28014
rect 11719 27962 11771 28014
rect 11771 27962 11848 28014
rect 11152 27949 11848 27962
rect 10666 27897 10721 27949
rect 10721 27897 10722 27949
rect 10747 27897 10773 27949
rect 10773 27897 10799 27949
rect 10799 27897 10803 27949
rect 10828 27897 10851 27949
rect 10851 27897 10884 27949
rect 10666 27893 10722 27897
rect 10747 27893 10803 27897
rect 10828 27893 10884 27897
rect 10909 27893 10965 27949
rect 10990 27893 11046 27949
rect 11071 27893 11127 27949
rect 11152 27897 11641 27949
rect 11641 27897 11693 27949
rect 11693 27897 11719 27949
rect 11719 27897 11771 27949
rect 11771 27897 11848 27949
rect 11152 27893 11848 27897
rect 3109 27038 3165 27094
rect 3190 27038 3246 27094
rect 3271 27038 3327 27094
rect 3352 27038 3408 27094
rect 3433 27038 3489 27094
rect 3109 26958 3165 27014
rect 3190 26958 3246 27014
rect 3271 26958 3327 27014
rect 3352 26958 3408 27014
rect 3433 26958 3489 27014
rect 3109 26878 3165 26934
rect 3190 26878 3246 26934
rect 3271 26878 3327 26934
rect 3352 26878 3408 26934
rect 3433 26878 3489 26934
rect 3109 26798 3165 26854
rect 3190 26798 3246 26854
rect 3271 26798 3327 26854
rect 3352 26798 3408 26854
rect 3433 26798 3489 26854
rect 3109 26718 3165 26774
rect 3190 26718 3246 26774
rect 3271 26718 3327 26774
rect 3352 26718 3408 26774
rect 3433 26718 3489 26774
rect 3109 26638 3165 26694
rect 3190 26638 3246 26694
rect 3271 26638 3327 26694
rect 3352 26638 3408 26694
rect 3433 26638 3489 26694
rect 3109 26558 3165 26614
rect 3190 26558 3246 26614
rect 3271 26558 3327 26614
rect 3352 26558 3408 26614
rect 3433 26558 3489 26614
rect 3109 26478 3165 26534
rect 3190 26478 3246 26534
rect 3271 26478 3327 26534
rect 3352 26478 3408 26534
rect 3433 26478 3489 26534
rect 3109 26398 3165 26454
rect 3190 26398 3246 26454
rect 3271 26398 3327 26454
rect 3352 26398 3408 26454
rect 3433 26398 3489 26454
rect 3109 26318 3165 26374
rect 3190 26318 3246 26374
rect 3271 26318 3327 26374
rect 3352 26318 3408 26374
rect 3433 26318 3489 26374
rect 3109 26238 3165 26294
rect 3190 26238 3246 26294
rect 3271 26238 3327 26294
rect 3352 26238 3408 26294
rect 3433 26238 3489 26294
rect 3109 26158 3165 26214
rect 3190 26158 3246 26214
rect 3271 26158 3327 26214
rect 3352 26158 3408 26214
rect 3433 26158 3489 26214
rect 3109 26078 3165 26134
rect 3190 26078 3246 26134
rect 3271 26078 3327 26134
rect 3352 26078 3408 26134
rect 3433 26078 3489 26134
rect 3109 25998 3165 26054
rect 3190 25998 3246 26054
rect 3271 25998 3327 26054
rect 3352 25998 3408 26054
rect 3433 25998 3489 26054
rect 3109 25918 3165 25974
rect 3190 25918 3246 25974
rect 3271 25918 3327 25974
rect 3352 25918 3408 25974
rect 3433 25918 3489 25974
rect 3109 25838 3165 25894
rect 3190 25838 3246 25894
rect 3271 25838 3327 25894
rect 3352 25838 3408 25894
rect 3433 25838 3489 25894
rect 3109 25758 3165 25814
rect 3190 25758 3246 25814
rect 3271 25758 3327 25814
rect 3352 25758 3408 25814
rect 3433 25758 3489 25814
rect 3109 25678 3165 25734
rect 3190 25678 3246 25734
rect 3271 25678 3327 25734
rect 3352 25678 3408 25734
rect 3433 25678 3489 25734
rect 3109 25598 3165 25654
rect 3190 25598 3246 25654
rect 3271 25598 3327 25654
rect 3352 25598 3408 25654
rect 3433 25598 3489 25654
rect 3109 25518 3165 25574
rect 3190 25518 3246 25574
rect 3271 25518 3327 25574
rect 3352 25518 3408 25574
rect 3433 25518 3489 25574
rect 3109 25438 3165 25494
rect 3190 25438 3246 25494
rect 3271 25438 3327 25494
rect 3352 25438 3408 25494
rect 3433 25438 3489 25494
rect 3109 25358 3165 25414
rect 3190 25358 3246 25414
rect 3271 25358 3327 25414
rect 3352 25358 3408 25414
rect 3433 25358 3489 25414
rect 3514 25358 4290 27094
rect 5195 27038 5251 27094
rect 5276 27038 5332 27094
rect 5357 27038 5413 27094
rect 5438 27038 5494 27094
rect 5519 27038 5575 27094
rect 5600 27090 6376 27094
rect 5600 27038 5632 27090
rect 5632 27038 5684 27090
rect 5684 27038 5700 27090
rect 5700 27038 5752 27090
rect 5752 27038 5768 27090
rect 5768 27038 5820 27090
rect 5820 27038 6376 27090
rect 5600 27026 6376 27038
rect 5195 26958 5251 27014
rect 5276 26958 5332 27014
rect 5357 26958 5413 27014
rect 5438 26958 5494 27014
rect 5519 26958 5575 27014
rect 5600 26974 5632 27026
rect 5632 26974 5684 27026
rect 5684 26974 5700 27026
rect 5700 26974 5752 27026
rect 5752 26974 5768 27026
rect 5768 26974 5820 27026
rect 5820 26974 6376 27026
rect 5600 26962 6376 26974
rect 5195 26878 5251 26934
rect 5276 26878 5332 26934
rect 5357 26878 5413 26934
rect 5438 26878 5494 26934
rect 5519 26878 5575 26934
rect 5600 26910 5632 26962
rect 5632 26910 5684 26962
rect 5684 26910 5700 26962
rect 5700 26910 5752 26962
rect 5752 26910 5768 26962
rect 5768 26910 5820 26962
rect 5820 26910 6376 26962
rect 5600 26898 6376 26910
rect 5195 26798 5251 26854
rect 5276 26798 5332 26854
rect 5357 26798 5413 26854
rect 5438 26798 5494 26854
rect 5519 26798 5575 26854
rect 5600 26846 5632 26898
rect 5632 26846 5684 26898
rect 5684 26846 5700 26898
rect 5700 26846 5752 26898
rect 5752 26846 5768 26898
rect 5768 26846 5820 26898
rect 5820 26846 6376 26898
rect 5600 26834 6376 26846
rect 5600 26782 5632 26834
rect 5632 26782 5684 26834
rect 5684 26782 5700 26834
rect 5700 26782 5752 26834
rect 5752 26782 5768 26834
rect 5768 26782 5820 26834
rect 5820 26782 6376 26834
rect 5195 26718 5251 26774
rect 5276 26718 5332 26774
rect 5357 26718 5413 26774
rect 5438 26718 5494 26774
rect 5519 26718 5575 26774
rect 5600 26770 6376 26782
rect 5600 26718 5632 26770
rect 5632 26718 5684 26770
rect 5684 26718 5700 26770
rect 5700 26718 5752 26770
rect 5752 26718 5768 26770
rect 5768 26718 5820 26770
rect 5820 26718 6376 26770
rect 5600 26706 6376 26718
rect 5195 26638 5251 26694
rect 5276 26638 5332 26694
rect 5357 26638 5413 26694
rect 5438 26638 5494 26694
rect 5519 26638 5575 26694
rect 5600 26654 5632 26706
rect 5632 26654 5684 26706
rect 5684 26654 5700 26706
rect 5700 26654 5752 26706
rect 5752 26654 5768 26706
rect 5768 26654 5820 26706
rect 5820 26654 6376 26706
rect 5600 26642 6376 26654
rect 5195 26558 5251 26614
rect 5276 26558 5332 26614
rect 5357 26558 5413 26614
rect 5438 26558 5494 26614
rect 5519 26558 5575 26614
rect 5600 26590 5632 26642
rect 5632 26590 5684 26642
rect 5684 26590 5700 26642
rect 5700 26590 5752 26642
rect 5752 26590 5768 26642
rect 5768 26590 5820 26642
rect 5820 26590 6376 26642
rect 5600 26578 6376 26590
rect 5195 26478 5251 26534
rect 5276 26478 5332 26534
rect 5357 26478 5413 26534
rect 5438 26478 5494 26534
rect 5519 26478 5575 26534
rect 5600 26526 5632 26578
rect 5632 26526 5684 26578
rect 5684 26526 5700 26578
rect 5700 26526 5752 26578
rect 5752 26526 5768 26578
rect 5768 26526 5820 26578
rect 5820 26526 6376 26578
rect 5600 26514 6376 26526
rect 5600 26462 5632 26514
rect 5632 26462 5684 26514
rect 5684 26462 5700 26514
rect 5700 26462 5752 26514
rect 5752 26462 5768 26514
rect 5768 26462 5820 26514
rect 5820 26462 6376 26514
rect 5195 26398 5251 26454
rect 5276 26398 5332 26454
rect 5357 26398 5413 26454
rect 5438 26398 5494 26454
rect 5519 26398 5575 26454
rect 5600 26450 6376 26462
rect 5600 26398 5632 26450
rect 5632 26398 5684 26450
rect 5684 26398 5700 26450
rect 5700 26398 5752 26450
rect 5752 26398 5768 26450
rect 5768 26398 5820 26450
rect 5820 26398 6376 26450
rect 5600 26386 6376 26398
rect 5195 26318 5251 26374
rect 5276 26318 5332 26374
rect 5357 26318 5413 26374
rect 5438 26318 5494 26374
rect 5519 26318 5575 26374
rect 5600 26334 5632 26386
rect 5632 26334 5684 26386
rect 5684 26334 5700 26386
rect 5700 26334 5752 26386
rect 5752 26334 5768 26386
rect 5768 26334 5820 26386
rect 5820 26334 6376 26386
rect 5600 26322 6376 26334
rect 5195 26238 5251 26294
rect 5276 26238 5332 26294
rect 5357 26238 5413 26294
rect 5438 26238 5494 26294
rect 5519 26238 5575 26294
rect 5600 26270 5632 26322
rect 5632 26270 5684 26322
rect 5684 26270 5700 26322
rect 5700 26270 5752 26322
rect 5752 26270 5768 26322
rect 5768 26270 5820 26322
rect 5820 26270 6376 26322
rect 5600 26258 6376 26270
rect 5195 26158 5251 26214
rect 5276 26158 5332 26214
rect 5357 26158 5413 26214
rect 5438 26158 5494 26214
rect 5519 26158 5575 26214
rect 5600 26206 5632 26258
rect 5632 26206 5684 26258
rect 5684 26206 5700 26258
rect 5700 26206 5752 26258
rect 5752 26206 5768 26258
rect 5768 26206 5820 26258
rect 5820 26206 6376 26258
rect 5600 26194 6376 26206
rect 5600 26142 5632 26194
rect 5632 26142 5684 26194
rect 5684 26142 5700 26194
rect 5700 26142 5752 26194
rect 5752 26142 5768 26194
rect 5768 26142 5820 26194
rect 5820 26142 6376 26194
rect 5195 26078 5251 26134
rect 5276 26078 5332 26134
rect 5357 26078 5413 26134
rect 5438 26078 5494 26134
rect 5519 26078 5575 26134
rect 5600 26129 6376 26142
rect 5600 26077 5632 26129
rect 5632 26077 5684 26129
rect 5684 26077 5700 26129
rect 5700 26077 5752 26129
rect 5752 26077 5768 26129
rect 5768 26077 5820 26129
rect 5820 26077 6376 26129
rect 5600 26064 6376 26077
rect 5195 25998 5251 26054
rect 5276 25998 5332 26054
rect 5357 25998 5413 26054
rect 5438 25998 5494 26054
rect 5519 25998 5575 26054
rect 5600 26012 5632 26064
rect 5632 26012 5684 26064
rect 5684 26012 5700 26064
rect 5700 26012 5752 26064
rect 5752 26012 5768 26064
rect 5768 26012 5820 26064
rect 5820 26012 6376 26064
rect 5600 25999 6376 26012
rect 5195 25918 5251 25974
rect 5276 25918 5332 25974
rect 5357 25918 5413 25974
rect 5438 25918 5494 25974
rect 5519 25918 5575 25974
rect 5600 25947 5632 25999
rect 5632 25947 5684 25999
rect 5684 25947 5700 25999
rect 5700 25947 5752 25999
rect 5752 25947 5768 25999
rect 5768 25947 5820 25999
rect 5820 25947 6376 25999
rect 5600 25934 6376 25947
rect 5195 25838 5251 25894
rect 5276 25838 5332 25894
rect 5357 25838 5413 25894
rect 5438 25838 5494 25894
rect 5519 25838 5575 25894
rect 5600 25882 5632 25934
rect 5632 25882 5684 25934
rect 5684 25882 5700 25934
rect 5700 25882 5752 25934
rect 5752 25882 5768 25934
rect 5768 25882 5820 25934
rect 5820 25882 6376 25934
rect 5600 25869 6376 25882
rect 5600 25817 5632 25869
rect 5632 25817 5684 25869
rect 5684 25817 5700 25869
rect 5700 25817 5752 25869
rect 5752 25817 5768 25869
rect 5768 25817 5820 25869
rect 5820 25817 6376 25869
rect 5195 25758 5251 25814
rect 5276 25758 5332 25814
rect 5357 25758 5413 25814
rect 5438 25758 5494 25814
rect 5519 25758 5575 25814
rect 5600 25804 6376 25817
rect 5600 25752 5632 25804
rect 5632 25752 5684 25804
rect 5684 25752 5700 25804
rect 5700 25752 5752 25804
rect 5752 25752 5768 25804
rect 5768 25752 5820 25804
rect 5820 25752 6376 25804
rect 5600 25739 6376 25752
rect 5195 25678 5251 25734
rect 5276 25678 5332 25734
rect 5357 25678 5413 25734
rect 5438 25678 5494 25734
rect 5519 25678 5575 25734
rect 5600 25687 5632 25739
rect 5632 25687 5684 25739
rect 5684 25687 5700 25739
rect 5700 25687 5752 25739
rect 5752 25687 5768 25739
rect 5768 25687 5820 25739
rect 5820 25687 6376 25739
rect 5600 25674 6376 25687
rect 5195 25598 5251 25654
rect 5276 25598 5332 25654
rect 5357 25598 5413 25654
rect 5438 25598 5494 25654
rect 5519 25598 5575 25654
rect 5600 25622 5632 25674
rect 5632 25622 5684 25674
rect 5684 25622 5700 25674
rect 5700 25622 5752 25674
rect 5752 25622 5768 25674
rect 5768 25622 5820 25674
rect 5820 25622 6376 25674
rect 5600 25609 6376 25622
rect 5195 25518 5251 25574
rect 5276 25518 5332 25574
rect 5357 25518 5413 25574
rect 5438 25518 5494 25574
rect 5519 25518 5575 25574
rect 5600 25557 5632 25609
rect 5632 25557 5684 25609
rect 5684 25557 5700 25609
rect 5700 25557 5752 25609
rect 5752 25557 5768 25609
rect 5768 25557 5820 25609
rect 5820 25557 6376 25609
rect 5600 25544 6376 25557
rect 5195 25438 5251 25494
rect 5276 25438 5332 25494
rect 5357 25438 5413 25494
rect 5438 25438 5494 25494
rect 5519 25438 5575 25494
rect 5600 25492 5632 25544
rect 5632 25492 5684 25544
rect 5684 25492 5700 25544
rect 5700 25492 5752 25544
rect 5752 25492 5768 25544
rect 5768 25492 5820 25544
rect 5820 25492 6376 25544
rect 5600 25479 6376 25492
rect 5600 25427 5632 25479
rect 5632 25427 5684 25479
rect 5684 25427 5700 25479
rect 5700 25427 5752 25479
rect 5752 25427 5768 25479
rect 5768 25427 5820 25479
rect 5820 25427 6376 25479
rect 5600 25414 6376 25427
rect 5195 25358 5251 25414
rect 5276 25358 5332 25414
rect 5357 25358 5413 25414
rect 5438 25358 5494 25414
rect 5519 25358 5575 25414
rect 5600 25362 5632 25414
rect 5632 25362 5684 25414
rect 5684 25362 5700 25414
rect 5700 25362 5752 25414
rect 5752 25362 5768 25414
rect 5768 25362 5820 25414
rect 5820 25362 6376 25414
rect 5600 25358 6376 25362
rect 8580 24973 8636 25029
rect 8661 24973 8717 25029
rect 8742 24973 8798 25029
rect 8823 24973 8879 25029
rect 8904 25025 8960 25029
rect 8985 25025 9041 25029
rect 8904 24973 8933 25025
rect 8933 24973 8959 25025
rect 8959 24973 8960 25025
rect 8985 24973 9011 25025
rect 9011 24973 9041 25025
rect 8580 24893 8636 24949
rect 8661 24893 8717 24949
rect 8742 24893 8798 24949
rect 8823 24893 8879 24949
rect 8904 24909 8933 24949
rect 8933 24909 8959 24949
rect 8959 24909 8960 24949
rect 8985 24909 9011 24949
rect 9011 24909 9041 24949
rect 8904 24897 8960 24909
rect 8985 24897 9041 24909
rect 8904 24893 8933 24897
rect 8933 24893 8959 24897
rect 8959 24893 8960 24897
rect 8985 24893 9011 24897
rect 9011 24893 9041 24897
rect 8580 24813 8636 24869
rect 8661 24813 8717 24869
rect 8742 24813 8798 24869
rect 8823 24813 8879 24869
rect 8904 24845 8933 24869
rect 8933 24845 8959 24869
rect 8959 24845 8960 24869
rect 8985 24845 9011 24869
rect 9011 24845 9041 24869
rect 8904 24833 8960 24845
rect 8985 24833 9041 24845
rect 8904 24813 8933 24833
rect 8933 24813 8959 24833
rect 8959 24813 8960 24833
rect 8985 24813 9011 24833
rect 9011 24813 9041 24833
rect 8580 24733 8636 24789
rect 8661 24733 8717 24789
rect 8742 24733 8798 24789
rect 8823 24733 8879 24789
rect 8904 24781 8933 24789
rect 8933 24781 8959 24789
rect 8959 24781 8960 24789
rect 8985 24781 9011 24789
rect 9011 24781 9041 24789
rect 8904 24769 8960 24781
rect 8985 24769 9041 24781
rect 8904 24733 8933 24769
rect 8933 24733 8959 24769
rect 8959 24733 8960 24769
rect 8985 24733 9011 24769
rect 9011 24733 9041 24769
rect 8580 24653 8636 24709
rect 8661 24653 8717 24709
rect 8742 24653 8798 24709
rect 8823 24653 8879 24709
rect 8904 24705 8960 24709
rect 8985 24705 9041 24709
rect 8904 24653 8933 24705
rect 8933 24653 8959 24705
rect 8959 24653 8960 24705
rect 8985 24653 9011 24705
rect 9011 24653 9041 24705
rect 8580 24573 8636 24629
rect 8661 24573 8717 24629
rect 8742 24573 8798 24629
rect 8823 24573 8879 24629
rect 8904 24589 8933 24629
rect 8933 24589 8959 24629
rect 8959 24589 8960 24629
rect 8985 24589 9011 24629
rect 9011 24589 9041 24629
rect 8904 24577 8960 24589
rect 8985 24577 9041 24589
rect 8904 24573 8933 24577
rect 8933 24573 8959 24577
rect 8959 24573 8960 24577
rect 8985 24573 9011 24577
rect 9011 24573 9041 24577
rect 8580 24493 8636 24549
rect 8661 24493 8717 24549
rect 8742 24493 8798 24549
rect 8823 24493 8879 24549
rect 8904 24525 8933 24549
rect 8933 24525 8959 24549
rect 8959 24525 8960 24549
rect 8985 24525 9011 24549
rect 9011 24525 9041 24549
rect 8904 24513 8960 24525
rect 8985 24513 9041 24525
rect 8904 24493 8933 24513
rect 8933 24493 8959 24513
rect 8959 24493 8960 24513
rect 8985 24493 9011 24513
rect 9011 24493 9041 24513
rect 8580 24413 8636 24469
rect 8661 24413 8717 24469
rect 8742 24413 8798 24469
rect 8823 24413 8879 24469
rect 8904 24461 8933 24469
rect 8933 24461 8959 24469
rect 8959 24461 8960 24469
rect 8985 24461 9011 24469
rect 9011 24461 9041 24469
rect 8904 24449 8960 24461
rect 8985 24449 9041 24461
rect 8904 24413 8933 24449
rect 8933 24413 8959 24449
rect 8959 24413 8960 24449
rect 8985 24413 9011 24449
rect 9011 24413 9041 24449
rect 8580 24333 8636 24389
rect 8661 24333 8717 24389
rect 8742 24333 8798 24389
rect 8823 24333 8879 24389
rect 8904 24385 8960 24389
rect 8985 24385 9041 24389
rect 8904 24333 8933 24385
rect 8933 24333 8959 24385
rect 8959 24333 8960 24385
rect 8985 24333 9011 24385
rect 9011 24333 9041 24385
rect 8580 24253 8636 24309
rect 8661 24253 8717 24309
rect 8742 24253 8798 24309
rect 8823 24253 8879 24309
rect 8904 24269 8933 24309
rect 8933 24269 8959 24309
rect 8959 24269 8960 24309
rect 8985 24269 9011 24309
rect 9011 24269 9041 24309
rect 8904 24257 8960 24269
rect 8985 24257 9041 24269
rect 8904 24253 8933 24257
rect 8933 24253 8959 24257
rect 8959 24253 8960 24257
rect 8985 24253 9011 24257
rect 9011 24253 9041 24257
rect 8580 24173 8636 24229
rect 8661 24173 8717 24229
rect 8742 24173 8798 24229
rect 8823 24173 8879 24229
rect 8904 24205 8933 24229
rect 8933 24205 8959 24229
rect 8959 24205 8960 24229
rect 8985 24205 9011 24229
rect 9011 24205 9041 24229
rect 8904 24193 8960 24205
rect 8985 24193 9041 24205
rect 8904 24173 8933 24193
rect 8933 24173 8959 24193
rect 8959 24173 8960 24193
rect 8985 24173 9011 24193
rect 9011 24173 9041 24193
rect 8580 24093 8636 24149
rect 8661 24093 8717 24149
rect 8742 24093 8798 24149
rect 8823 24093 8879 24149
rect 8904 24141 8933 24149
rect 8933 24141 8959 24149
rect 8959 24141 8960 24149
rect 8985 24141 9011 24149
rect 9011 24141 9041 24149
rect 8904 24129 8960 24141
rect 8985 24129 9041 24141
rect 8904 24093 8933 24129
rect 8933 24093 8959 24129
rect 8959 24093 8960 24129
rect 8985 24093 9011 24129
rect 9011 24093 9041 24129
rect 8580 24013 8636 24069
rect 8661 24013 8717 24069
rect 8742 24013 8798 24069
rect 8823 24013 8879 24069
rect 8904 24064 8960 24069
rect 8985 24064 9041 24069
rect 8904 24013 8933 24064
rect 8933 24013 8959 24064
rect 8959 24013 8960 24064
rect 8985 24013 9011 24064
rect 9011 24013 9041 24064
rect 8580 23933 8636 23989
rect 8661 23933 8717 23989
rect 8742 23933 8798 23989
rect 8823 23933 8879 23989
rect 8904 23947 8933 23989
rect 8933 23947 8959 23989
rect 8959 23947 8960 23989
rect 8985 23947 9011 23989
rect 9011 23947 9041 23989
rect 8904 23934 8960 23947
rect 8985 23934 9041 23947
rect 8904 23933 8933 23934
rect 8933 23933 8959 23934
rect 8959 23933 8960 23934
rect 8985 23933 9011 23934
rect 9011 23933 9041 23934
rect 8580 23853 8636 23909
rect 8661 23853 8717 23909
rect 8742 23853 8798 23909
rect 8823 23853 8879 23909
rect 8904 23882 8933 23909
rect 8933 23882 8959 23909
rect 8959 23882 8960 23909
rect 8985 23882 9011 23909
rect 9011 23882 9041 23909
rect 8904 23869 8960 23882
rect 8985 23869 9041 23882
rect 8904 23853 8933 23869
rect 8933 23853 8959 23869
rect 8959 23853 8960 23869
rect 8985 23853 9011 23869
rect 9011 23853 9041 23869
rect 8580 23773 8636 23829
rect 8661 23773 8717 23829
rect 8742 23773 8798 23829
rect 8823 23773 8879 23829
rect 8904 23817 8933 23829
rect 8933 23817 8959 23829
rect 8959 23817 8960 23829
rect 8985 23817 9011 23829
rect 9011 23817 9041 23829
rect 8904 23804 8960 23817
rect 8985 23804 9041 23817
rect 8904 23773 8933 23804
rect 8933 23773 8959 23804
rect 8959 23773 8960 23804
rect 8985 23773 9011 23804
rect 9011 23773 9041 23804
rect 8580 23693 8636 23749
rect 8661 23693 8717 23749
rect 8742 23693 8798 23749
rect 8823 23693 8879 23749
rect 8904 23739 8960 23749
rect 8985 23739 9041 23749
rect 8904 23693 8933 23739
rect 8933 23693 8959 23739
rect 8959 23693 8960 23739
rect 8985 23693 9011 23739
rect 9011 23693 9041 23739
rect 8580 23613 8636 23669
rect 8661 23613 8717 23669
rect 8742 23613 8798 23669
rect 8823 23613 8879 23669
rect 8904 23622 8933 23669
rect 8933 23622 8959 23669
rect 8959 23622 8960 23669
rect 8985 23622 9011 23669
rect 9011 23622 9041 23669
rect 8904 23613 8960 23622
rect 8985 23613 9041 23622
rect 8580 23533 8636 23589
rect 8661 23533 8717 23589
rect 8742 23533 8798 23589
rect 8823 23533 8879 23589
rect 8904 23557 8933 23589
rect 8933 23557 8959 23589
rect 8959 23557 8960 23589
rect 8985 23557 9011 23589
rect 9011 23557 9041 23589
rect 8904 23544 8960 23557
rect 8985 23544 9041 23557
rect 8904 23533 8933 23544
rect 8933 23533 8959 23544
rect 8959 23533 8960 23544
rect 8985 23533 9011 23544
rect 9011 23533 9041 23544
rect 8580 23453 8636 23509
rect 8661 23453 8717 23509
rect 8742 23453 8798 23509
rect 8823 23453 8879 23509
rect 8904 23492 8933 23509
rect 8933 23492 8959 23509
rect 8959 23492 8960 23509
rect 8985 23492 9011 23509
rect 9011 23492 9041 23509
rect 8904 23479 8960 23492
rect 8985 23479 9041 23492
rect 8904 23453 8933 23479
rect 8933 23453 8959 23479
rect 8959 23453 8960 23479
rect 8985 23453 9011 23479
rect 9011 23453 9041 23479
rect 8580 23373 8636 23429
rect 8661 23373 8717 23429
rect 8742 23373 8798 23429
rect 8823 23373 8879 23429
rect 8904 23427 8933 23429
rect 8933 23427 8959 23429
rect 8959 23427 8960 23429
rect 8985 23427 9011 23429
rect 9011 23427 9041 23429
rect 8904 23414 8960 23427
rect 8985 23414 9041 23427
rect 8904 23373 8933 23414
rect 8933 23373 8959 23414
rect 8959 23373 8960 23414
rect 8985 23373 9011 23414
rect 9011 23373 9041 23414
rect 8580 23293 8636 23349
rect 8661 23293 8717 23349
rect 8742 23293 8798 23349
rect 8823 23293 8879 23349
rect 8904 23297 8933 23349
rect 8933 23297 8959 23349
rect 8959 23297 8960 23349
rect 8985 23297 9011 23349
rect 9011 23297 9041 23349
rect 8904 23293 8960 23297
rect 8985 23293 9041 23297
rect 9066 23293 9762 25029
rect 10666 25025 10722 25029
rect 10747 25025 10803 25029
rect 10828 25025 10884 25029
rect 10666 24973 10721 25025
rect 10721 24973 10722 25025
rect 10747 24973 10773 25025
rect 10773 24973 10799 25025
rect 10799 24973 10803 25025
rect 10828 24973 10851 25025
rect 10851 24973 10884 25025
rect 10909 24973 10965 25029
rect 10990 24973 11046 25029
rect 11071 24973 11127 25029
rect 11152 25025 11848 25029
rect 11152 24973 11641 25025
rect 11641 24973 11693 25025
rect 11693 24973 11719 25025
rect 11719 24973 11771 25025
rect 11771 24973 11848 25025
rect 11152 24961 11848 24973
rect 10666 24909 10721 24949
rect 10721 24909 10722 24949
rect 10747 24909 10773 24949
rect 10773 24909 10799 24949
rect 10799 24909 10803 24949
rect 10828 24909 10851 24949
rect 10851 24909 10884 24949
rect 10666 24897 10722 24909
rect 10747 24897 10803 24909
rect 10828 24897 10884 24909
rect 10666 24893 10721 24897
rect 10721 24893 10722 24897
rect 10747 24893 10773 24897
rect 10773 24893 10799 24897
rect 10799 24893 10803 24897
rect 10828 24893 10851 24897
rect 10851 24893 10884 24897
rect 10909 24893 10965 24949
rect 10990 24893 11046 24949
rect 11071 24893 11127 24949
rect 11152 24909 11641 24961
rect 11641 24909 11693 24961
rect 11693 24909 11719 24961
rect 11719 24909 11771 24961
rect 11771 24909 11848 24961
rect 11152 24897 11848 24909
rect 10666 24845 10721 24869
rect 10721 24845 10722 24869
rect 10747 24845 10773 24869
rect 10773 24845 10799 24869
rect 10799 24845 10803 24869
rect 10828 24845 10851 24869
rect 10851 24845 10884 24869
rect 10666 24833 10722 24845
rect 10747 24833 10803 24845
rect 10828 24833 10884 24845
rect 10666 24813 10721 24833
rect 10721 24813 10722 24833
rect 10747 24813 10773 24833
rect 10773 24813 10799 24833
rect 10799 24813 10803 24833
rect 10828 24813 10851 24833
rect 10851 24813 10884 24833
rect 10909 24813 10965 24869
rect 10990 24813 11046 24869
rect 11071 24813 11127 24869
rect 11152 24845 11641 24897
rect 11641 24845 11693 24897
rect 11693 24845 11719 24897
rect 11719 24845 11771 24897
rect 11771 24845 11848 24897
rect 11152 24833 11848 24845
rect 10666 24781 10721 24789
rect 10721 24781 10722 24789
rect 10747 24781 10773 24789
rect 10773 24781 10799 24789
rect 10799 24781 10803 24789
rect 10828 24781 10851 24789
rect 10851 24781 10884 24789
rect 10666 24769 10722 24781
rect 10747 24769 10803 24781
rect 10828 24769 10884 24781
rect 10666 24733 10721 24769
rect 10721 24733 10722 24769
rect 10747 24733 10773 24769
rect 10773 24733 10799 24769
rect 10799 24733 10803 24769
rect 10828 24733 10851 24769
rect 10851 24733 10884 24769
rect 10909 24733 10965 24789
rect 10990 24733 11046 24789
rect 11071 24733 11127 24789
rect 11152 24781 11641 24833
rect 11641 24781 11693 24833
rect 11693 24781 11719 24833
rect 11719 24781 11771 24833
rect 11771 24781 11848 24833
rect 11152 24769 11848 24781
rect 11152 24717 11641 24769
rect 11641 24717 11693 24769
rect 11693 24717 11719 24769
rect 11719 24717 11771 24769
rect 11771 24717 11848 24769
rect 10666 24705 10722 24709
rect 10747 24705 10803 24709
rect 10828 24705 10884 24709
rect 10666 24653 10721 24705
rect 10721 24653 10722 24705
rect 10747 24653 10773 24705
rect 10773 24653 10799 24705
rect 10799 24653 10803 24705
rect 10828 24653 10851 24705
rect 10851 24653 10884 24705
rect 10909 24653 10965 24709
rect 10990 24653 11046 24709
rect 11071 24653 11127 24709
rect 11152 24705 11848 24717
rect 11152 24653 11641 24705
rect 11641 24653 11693 24705
rect 11693 24653 11719 24705
rect 11719 24653 11771 24705
rect 11771 24653 11848 24705
rect 11152 24641 11848 24653
rect 10666 24589 10721 24629
rect 10721 24589 10722 24629
rect 10747 24589 10773 24629
rect 10773 24589 10799 24629
rect 10799 24589 10803 24629
rect 10828 24589 10851 24629
rect 10851 24589 10884 24629
rect 10666 24577 10722 24589
rect 10747 24577 10803 24589
rect 10828 24577 10884 24589
rect 10666 24573 10721 24577
rect 10721 24573 10722 24577
rect 10747 24573 10773 24577
rect 10773 24573 10799 24577
rect 10799 24573 10803 24577
rect 10828 24573 10851 24577
rect 10851 24573 10884 24577
rect 10909 24573 10965 24629
rect 10990 24573 11046 24629
rect 11071 24573 11127 24629
rect 11152 24589 11641 24641
rect 11641 24589 11693 24641
rect 11693 24589 11719 24641
rect 11719 24589 11771 24641
rect 11771 24589 11848 24641
rect 11152 24577 11848 24589
rect 10666 24525 10721 24549
rect 10721 24525 10722 24549
rect 10747 24525 10773 24549
rect 10773 24525 10799 24549
rect 10799 24525 10803 24549
rect 10828 24525 10851 24549
rect 10851 24525 10884 24549
rect 10666 24513 10722 24525
rect 10747 24513 10803 24525
rect 10828 24513 10884 24525
rect 10666 24493 10721 24513
rect 10721 24493 10722 24513
rect 10747 24493 10773 24513
rect 10773 24493 10799 24513
rect 10799 24493 10803 24513
rect 10828 24493 10851 24513
rect 10851 24493 10884 24513
rect 10909 24493 10965 24549
rect 10990 24493 11046 24549
rect 11071 24493 11127 24549
rect 11152 24525 11641 24577
rect 11641 24525 11693 24577
rect 11693 24525 11719 24577
rect 11719 24525 11771 24577
rect 11771 24525 11848 24577
rect 11152 24513 11848 24525
rect 10666 24461 10721 24469
rect 10721 24461 10722 24469
rect 10747 24461 10773 24469
rect 10773 24461 10799 24469
rect 10799 24461 10803 24469
rect 10828 24461 10851 24469
rect 10851 24461 10884 24469
rect 10666 24449 10722 24461
rect 10747 24449 10803 24461
rect 10828 24449 10884 24461
rect 10666 24413 10721 24449
rect 10721 24413 10722 24449
rect 10747 24413 10773 24449
rect 10773 24413 10799 24449
rect 10799 24413 10803 24449
rect 10828 24413 10851 24449
rect 10851 24413 10884 24449
rect 10909 24413 10965 24469
rect 10990 24413 11046 24469
rect 11071 24413 11127 24469
rect 11152 24461 11641 24513
rect 11641 24461 11693 24513
rect 11693 24461 11719 24513
rect 11719 24461 11771 24513
rect 11771 24461 11848 24513
rect 11152 24449 11848 24461
rect 11152 24397 11641 24449
rect 11641 24397 11693 24449
rect 11693 24397 11719 24449
rect 11719 24397 11771 24449
rect 11771 24397 11848 24449
rect 10666 24385 10722 24389
rect 10747 24385 10803 24389
rect 10828 24385 10884 24389
rect 10666 24333 10721 24385
rect 10721 24333 10722 24385
rect 10747 24333 10773 24385
rect 10773 24333 10799 24385
rect 10799 24333 10803 24385
rect 10828 24333 10851 24385
rect 10851 24333 10884 24385
rect 10909 24333 10965 24389
rect 10990 24333 11046 24389
rect 11071 24333 11127 24389
rect 11152 24385 11848 24397
rect 11152 24333 11641 24385
rect 11641 24333 11693 24385
rect 11693 24333 11719 24385
rect 11719 24333 11771 24385
rect 11771 24333 11848 24385
rect 11152 24321 11848 24333
rect 10666 24269 10721 24309
rect 10721 24269 10722 24309
rect 10747 24269 10773 24309
rect 10773 24269 10799 24309
rect 10799 24269 10803 24309
rect 10828 24269 10851 24309
rect 10851 24269 10884 24309
rect 10666 24257 10722 24269
rect 10747 24257 10803 24269
rect 10828 24257 10884 24269
rect 10666 24253 10721 24257
rect 10721 24253 10722 24257
rect 10747 24253 10773 24257
rect 10773 24253 10799 24257
rect 10799 24253 10803 24257
rect 10828 24253 10851 24257
rect 10851 24253 10884 24257
rect 10909 24253 10965 24309
rect 10990 24253 11046 24309
rect 11071 24253 11127 24309
rect 11152 24269 11641 24321
rect 11641 24269 11693 24321
rect 11693 24269 11719 24321
rect 11719 24269 11771 24321
rect 11771 24269 11848 24321
rect 11152 24257 11848 24269
rect 10666 24205 10721 24229
rect 10721 24205 10722 24229
rect 10747 24205 10773 24229
rect 10773 24205 10799 24229
rect 10799 24205 10803 24229
rect 10828 24205 10851 24229
rect 10851 24205 10884 24229
rect 10666 24193 10722 24205
rect 10747 24193 10803 24205
rect 10828 24193 10884 24205
rect 10666 24173 10721 24193
rect 10721 24173 10722 24193
rect 10747 24173 10773 24193
rect 10773 24173 10799 24193
rect 10799 24173 10803 24193
rect 10828 24173 10851 24193
rect 10851 24173 10884 24193
rect 10909 24173 10965 24229
rect 10990 24173 11046 24229
rect 11071 24173 11127 24229
rect 11152 24205 11641 24257
rect 11641 24205 11693 24257
rect 11693 24205 11719 24257
rect 11719 24205 11771 24257
rect 11771 24205 11848 24257
rect 11152 24193 11848 24205
rect 10666 24141 10721 24149
rect 10721 24141 10722 24149
rect 10747 24141 10773 24149
rect 10773 24141 10799 24149
rect 10799 24141 10803 24149
rect 10828 24141 10851 24149
rect 10851 24141 10884 24149
rect 10666 24129 10722 24141
rect 10747 24129 10803 24141
rect 10828 24129 10884 24141
rect 10666 24093 10721 24129
rect 10721 24093 10722 24129
rect 10747 24093 10773 24129
rect 10773 24093 10799 24129
rect 10799 24093 10803 24129
rect 10828 24093 10851 24129
rect 10851 24093 10884 24129
rect 10909 24093 10965 24149
rect 10990 24093 11046 24149
rect 11071 24093 11127 24149
rect 11152 24141 11641 24193
rect 11641 24141 11693 24193
rect 11693 24141 11719 24193
rect 11719 24141 11771 24193
rect 11771 24141 11848 24193
rect 11152 24129 11848 24141
rect 11152 24077 11641 24129
rect 11641 24077 11693 24129
rect 11693 24077 11719 24129
rect 11719 24077 11771 24129
rect 11771 24077 11848 24129
rect 10666 24064 10722 24069
rect 10747 24064 10803 24069
rect 10828 24064 10884 24069
rect 10666 24013 10721 24064
rect 10721 24013 10722 24064
rect 10747 24013 10773 24064
rect 10773 24013 10799 24064
rect 10799 24013 10803 24064
rect 10828 24013 10851 24064
rect 10851 24013 10884 24064
rect 10909 24013 10965 24069
rect 10990 24013 11046 24069
rect 11071 24013 11127 24069
rect 11152 24064 11848 24077
rect 11152 24012 11641 24064
rect 11641 24012 11693 24064
rect 11693 24012 11719 24064
rect 11719 24012 11771 24064
rect 11771 24012 11848 24064
rect 11152 23999 11848 24012
rect 10666 23947 10721 23989
rect 10721 23947 10722 23989
rect 10747 23947 10773 23989
rect 10773 23947 10799 23989
rect 10799 23947 10803 23989
rect 10828 23947 10851 23989
rect 10851 23947 10884 23989
rect 10666 23934 10722 23947
rect 10747 23934 10803 23947
rect 10828 23934 10884 23947
rect 10666 23933 10721 23934
rect 10721 23933 10722 23934
rect 10747 23933 10773 23934
rect 10773 23933 10799 23934
rect 10799 23933 10803 23934
rect 10828 23933 10851 23934
rect 10851 23933 10884 23934
rect 10909 23933 10965 23989
rect 10990 23933 11046 23989
rect 11071 23933 11127 23989
rect 11152 23947 11641 23999
rect 11641 23947 11693 23999
rect 11693 23947 11719 23999
rect 11719 23947 11771 23999
rect 11771 23947 11848 23999
rect 11152 23934 11848 23947
rect 10666 23882 10721 23909
rect 10721 23882 10722 23909
rect 10747 23882 10773 23909
rect 10773 23882 10799 23909
rect 10799 23882 10803 23909
rect 10828 23882 10851 23909
rect 10851 23882 10884 23909
rect 10666 23869 10722 23882
rect 10747 23869 10803 23882
rect 10828 23869 10884 23882
rect 10666 23853 10721 23869
rect 10721 23853 10722 23869
rect 10747 23853 10773 23869
rect 10773 23853 10799 23869
rect 10799 23853 10803 23869
rect 10828 23853 10851 23869
rect 10851 23853 10884 23869
rect 10909 23853 10965 23909
rect 10990 23853 11046 23909
rect 11071 23853 11127 23909
rect 11152 23882 11641 23934
rect 11641 23882 11693 23934
rect 11693 23882 11719 23934
rect 11719 23882 11771 23934
rect 11771 23882 11848 23934
rect 11152 23869 11848 23882
rect 10666 23817 10721 23829
rect 10721 23817 10722 23829
rect 10747 23817 10773 23829
rect 10773 23817 10799 23829
rect 10799 23817 10803 23829
rect 10828 23817 10851 23829
rect 10851 23817 10884 23829
rect 10666 23804 10722 23817
rect 10747 23804 10803 23817
rect 10828 23804 10884 23817
rect 10666 23773 10721 23804
rect 10721 23773 10722 23804
rect 10747 23773 10773 23804
rect 10773 23773 10799 23804
rect 10799 23773 10803 23804
rect 10828 23773 10851 23804
rect 10851 23773 10884 23804
rect 10909 23773 10965 23829
rect 10990 23773 11046 23829
rect 11071 23773 11127 23829
rect 11152 23817 11641 23869
rect 11641 23817 11693 23869
rect 11693 23817 11719 23869
rect 11719 23817 11771 23869
rect 11771 23817 11848 23869
rect 11152 23804 11848 23817
rect 11152 23752 11641 23804
rect 11641 23752 11693 23804
rect 11693 23752 11719 23804
rect 11719 23752 11771 23804
rect 11771 23752 11848 23804
rect 10666 23739 10722 23749
rect 10747 23739 10803 23749
rect 10828 23739 10884 23749
rect 10666 23693 10721 23739
rect 10721 23693 10722 23739
rect 10747 23693 10773 23739
rect 10773 23693 10799 23739
rect 10799 23693 10803 23739
rect 10828 23693 10851 23739
rect 10851 23693 10884 23739
rect 10909 23693 10965 23749
rect 10990 23693 11046 23749
rect 11071 23693 11127 23749
rect 11152 23739 11848 23752
rect 11152 23687 11641 23739
rect 11641 23687 11693 23739
rect 11693 23687 11719 23739
rect 11719 23687 11771 23739
rect 11771 23687 11848 23739
rect 11152 23674 11848 23687
rect 10666 23622 10721 23669
rect 10721 23622 10722 23669
rect 10747 23622 10773 23669
rect 10773 23622 10799 23669
rect 10799 23622 10803 23669
rect 10828 23622 10851 23669
rect 10851 23622 10884 23669
rect 10666 23613 10722 23622
rect 10747 23613 10803 23622
rect 10828 23613 10884 23622
rect 10909 23613 10965 23669
rect 10990 23613 11046 23669
rect 11071 23613 11127 23669
rect 11152 23622 11641 23674
rect 11641 23622 11693 23674
rect 11693 23622 11719 23674
rect 11719 23622 11771 23674
rect 11771 23622 11848 23674
rect 11152 23609 11848 23622
rect 10666 23557 10721 23589
rect 10721 23557 10722 23589
rect 10747 23557 10773 23589
rect 10773 23557 10799 23589
rect 10799 23557 10803 23589
rect 10828 23557 10851 23589
rect 10851 23557 10884 23589
rect 10666 23544 10722 23557
rect 10747 23544 10803 23557
rect 10828 23544 10884 23557
rect 10666 23533 10721 23544
rect 10721 23533 10722 23544
rect 10747 23533 10773 23544
rect 10773 23533 10799 23544
rect 10799 23533 10803 23544
rect 10828 23533 10851 23544
rect 10851 23533 10884 23544
rect 10909 23533 10965 23589
rect 10990 23533 11046 23589
rect 11071 23533 11127 23589
rect 11152 23557 11641 23609
rect 11641 23557 11693 23609
rect 11693 23557 11719 23609
rect 11719 23557 11771 23609
rect 11771 23557 11848 23609
rect 11152 23544 11848 23557
rect 10666 23492 10721 23509
rect 10721 23492 10722 23509
rect 10747 23492 10773 23509
rect 10773 23492 10799 23509
rect 10799 23492 10803 23509
rect 10828 23492 10851 23509
rect 10851 23492 10884 23509
rect 10666 23479 10722 23492
rect 10747 23479 10803 23492
rect 10828 23479 10884 23492
rect 10666 23453 10721 23479
rect 10721 23453 10722 23479
rect 10747 23453 10773 23479
rect 10773 23453 10799 23479
rect 10799 23453 10803 23479
rect 10828 23453 10851 23479
rect 10851 23453 10884 23479
rect 10909 23453 10965 23509
rect 10990 23453 11046 23509
rect 11071 23453 11127 23509
rect 11152 23492 11641 23544
rect 11641 23492 11693 23544
rect 11693 23492 11719 23544
rect 11719 23492 11771 23544
rect 11771 23492 11848 23544
rect 11152 23479 11848 23492
rect 10666 23427 10721 23429
rect 10721 23427 10722 23429
rect 10747 23427 10773 23429
rect 10773 23427 10799 23429
rect 10799 23427 10803 23429
rect 10828 23427 10851 23429
rect 10851 23427 10884 23429
rect 10666 23414 10722 23427
rect 10747 23414 10803 23427
rect 10828 23414 10884 23427
rect 10666 23373 10721 23414
rect 10721 23373 10722 23414
rect 10747 23373 10773 23414
rect 10773 23373 10799 23414
rect 10799 23373 10803 23414
rect 10828 23373 10851 23414
rect 10851 23373 10884 23414
rect 10909 23373 10965 23429
rect 10990 23373 11046 23429
rect 11071 23373 11127 23429
rect 11152 23427 11641 23479
rect 11641 23427 11693 23479
rect 11693 23427 11719 23479
rect 11719 23427 11771 23479
rect 11771 23427 11848 23479
rect 11152 23414 11848 23427
rect 11152 23362 11641 23414
rect 11641 23362 11693 23414
rect 11693 23362 11719 23414
rect 11719 23362 11771 23414
rect 11771 23362 11848 23414
rect 11152 23349 11848 23362
rect 10666 23297 10721 23349
rect 10721 23297 10722 23349
rect 10747 23297 10773 23349
rect 10773 23297 10799 23349
rect 10799 23297 10803 23349
rect 10828 23297 10851 23349
rect 10851 23297 10884 23349
rect 10666 23293 10722 23297
rect 10747 23293 10803 23297
rect 10828 23293 10884 23297
rect 10909 23293 10965 23349
rect 10990 23293 11046 23349
rect 11071 23293 11127 23349
rect 11152 23297 11641 23349
rect 11641 23297 11693 23349
rect 11693 23297 11719 23349
rect 11719 23297 11771 23349
rect 11771 23297 11848 23349
rect 11152 23293 11848 23297
rect 3109 22438 3165 22494
rect 3190 22438 3246 22494
rect 3271 22438 3327 22494
rect 3352 22438 3408 22494
rect 3433 22438 3489 22494
rect 3109 22358 3165 22414
rect 3190 22358 3246 22414
rect 3271 22358 3327 22414
rect 3352 22358 3408 22414
rect 3433 22358 3489 22414
rect 3109 22278 3165 22334
rect 3190 22278 3246 22334
rect 3271 22278 3327 22334
rect 3352 22278 3408 22334
rect 3433 22278 3489 22334
rect 3109 22198 3165 22254
rect 3190 22198 3246 22254
rect 3271 22198 3327 22254
rect 3352 22198 3408 22254
rect 3433 22198 3489 22254
rect 3109 22118 3165 22174
rect 3190 22118 3246 22174
rect 3271 22118 3327 22174
rect 3352 22118 3408 22174
rect 3433 22118 3489 22174
rect 3109 22038 3165 22094
rect 3190 22038 3246 22094
rect 3271 22038 3327 22094
rect 3352 22038 3408 22094
rect 3433 22038 3489 22094
rect 3109 21958 3165 22014
rect 3190 21958 3246 22014
rect 3271 21958 3327 22014
rect 3352 21958 3408 22014
rect 3433 21958 3489 22014
rect 3109 21878 3165 21934
rect 3190 21878 3246 21934
rect 3271 21878 3327 21934
rect 3352 21878 3408 21934
rect 3433 21878 3489 21934
rect 3109 21798 3165 21854
rect 3190 21798 3246 21854
rect 3271 21798 3327 21854
rect 3352 21798 3408 21854
rect 3433 21798 3489 21854
rect 3109 21718 3165 21774
rect 3190 21718 3246 21774
rect 3271 21718 3327 21774
rect 3352 21718 3408 21774
rect 3433 21718 3489 21774
rect 3109 21638 3165 21694
rect 3190 21638 3246 21694
rect 3271 21638 3327 21694
rect 3352 21638 3408 21694
rect 3433 21638 3489 21694
rect 3109 21558 3165 21614
rect 3190 21558 3246 21614
rect 3271 21558 3327 21614
rect 3352 21558 3408 21614
rect 3433 21558 3489 21614
rect 3109 21478 3165 21534
rect 3190 21478 3246 21534
rect 3271 21478 3327 21534
rect 3352 21478 3408 21534
rect 3433 21478 3489 21534
rect 3109 21398 3165 21454
rect 3190 21398 3246 21454
rect 3271 21398 3327 21454
rect 3352 21398 3408 21454
rect 3433 21398 3489 21454
rect 3109 21318 3165 21374
rect 3190 21318 3246 21374
rect 3271 21318 3327 21374
rect 3352 21318 3408 21374
rect 3433 21318 3489 21374
rect 3109 21238 3165 21294
rect 3190 21238 3246 21294
rect 3271 21238 3327 21294
rect 3352 21238 3408 21294
rect 3433 21238 3489 21294
rect 3109 21158 3165 21214
rect 3190 21158 3246 21214
rect 3271 21158 3327 21214
rect 3352 21158 3408 21214
rect 3433 21158 3489 21214
rect 3109 21078 3165 21134
rect 3190 21078 3246 21134
rect 3271 21078 3327 21134
rect 3352 21078 3408 21134
rect 3433 21078 3489 21134
rect 3109 20998 3165 21054
rect 3190 20998 3246 21054
rect 3271 20998 3327 21054
rect 3352 20998 3408 21054
rect 3433 20998 3489 21054
rect 3109 20918 3165 20974
rect 3190 20918 3246 20974
rect 3271 20918 3327 20974
rect 3352 20918 3408 20974
rect 3433 20918 3489 20974
rect 3109 20838 3165 20894
rect 3190 20838 3246 20894
rect 3271 20838 3327 20894
rect 3352 20838 3408 20894
rect 3433 20838 3489 20894
rect 3109 20758 3165 20814
rect 3190 20758 3246 20814
rect 3271 20758 3327 20814
rect 3352 20758 3408 20814
rect 3433 20758 3489 20814
rect 3514 20758 4290 22494
rect 5195 22438 5251 22494
rect 5276 22438 5332 22494
rect 5357 22438 5413 22494
rect 5438 22438 5494 22494
rect 5519 22438 5575 22494
rect 5600 22490 6376 22494
rect 5600 22438 5632 22490
rect 5632 22438 5684 22490
rect 5684 22438 5700 22490
rect 5700 22438 5752 22490
rect 5752 22438 5768 22490
rect 5768 22438 5820 22490
rect 5820 22438 6376 22490
rect 5600 22426 6376 22438
rect 5195 22358 5251 22414
rect 5276 22358 5332 22414
rect 5357 22358 5413 22414
rect 5438 22358 5494 22414
rect 5519 22358 5575 22414
rect 5600 22374 5632 22426
rect 5632 22374 5684 22426
rect 5684 22374 5700 22426
rect 5700 22374 5752 22426
rect 5752 22374 5768 22426
rect 5768 22374 5820 22426
rect 5820 22374 6376 22426
rect 5600 22362 6376 22374
rect 5195 22278 5251 22334
rect 5276 22278 5332 22334
rect 5357 22278 5413 22334
rect 5438 22278 5494 22334
rect 5519 22278 5575 22334
rect 5600 22310 5632 22362
rect 5632 22310 5684 22362
rect 5684 22310 5700 22362
rect 5700 22310 5752 22362
rect 5752 22310 5768 22362
rect 5768 22310 5820 22362
rect 5820 22310 6376 22362
rect 5600 22298 6376 22310
rect 5195 22198 5251 22254
rect 5276 22198 5332 22254
rect 5357 22198 5413 22254
rect 5438 22198 5494 22254
rect 5519 22198 5575 22254
rect 5600 22246 5632 22298
rect 5632 22246 5684 22298
rect 5684 22246 5700 22298
rect 5700 22246 5752 22298
rect 5752 22246 5768 22298
rect 5768 22246 5820 22298
rect 5820 22246 6376 22298
rect 5600 22234 6376 22246
rect 5600 22182 5632 22234
rect 5632 22182 5684 22234
rect 5684 22182 5700 22234
rect 5700 22182 5752 22234
rect 5752 22182 5768 22234
rect 5768 22182 5820 22234
rect 5820 22182 6376 22234
rect 5195 22118 5251 22174
rect 5276 22118 5332 22174
rect 5357 22118 5413 22174
rect 5438 22118 5494 22174
rect 5519 22118 5575 22174
rect 5600 22170 6376 22182
rect 5600 22118 5632 22170
rect 5632 22118 5684 22170
rect 5684 22118 5700 22170
rect 5700 22118 5752 22170
rect 5752 22118 5768 22170
rect 5768 22118 5820 22170
rect 5820 22118 6376 22170
rect 5600 22106 6376 22118
rect 5195 22038 5251 22094
rect 5276 22038 5332 22094
rect 5357 22038 5413 22094
rect 5438 22038 5494 22094
rect 5519 22038 5575 22094
rect 5600 22054 5632 22106
rect 5632 22054 5684 22106
rect 5684 22054 5700 22106
rect 5700 22054 5752 22106
rect 5752 22054 5768 22106
rect 5768 22054 5820 22106
rect 5820 22054 6376 22106
rect 5600 22042 6376 22054
rect 5195 21958 5251 22014
rect 5276 21958 5332 22014
rect 5357 21958 5413 22014
rect 5438 21958 5494 22014
rect 5519 21958 5575 22014
rect 5600 21990 5632 22042
rect 5632 21990 5684 22042
rect 5684 21990 5700 22042
rect 5700 21990 5752 22042
rect 5752 21990 5768 22042
rect 5768 21990 5820 22042
rect 5820 21990 6376 22042
rect 5600 21978 6376 21990
rect 5195 21878 5251 21934
rect 5276 21878 5332 21934
rect 5357 21878 5413 21934
rect 5438 21878 5494 21934
rect 5519 21878 5575 21934
rect 5600 21926 5632 21978
rect 5632 21926 5684 21978
rect 5684 21926 5700 21978
rect 5700 21926 5752 21978
rect 5752 21926 5768 21978
rect 5768 21926 5820 21978
rect 5820 21926 6376 21978
rect 5600 21914 6376 21926
rect 5600 21862 5632 21914
rect 5632 21862 5684 21914
rect 5684 21862 5700 21914
rect 5700 21862 5752 21914
rect 5752 21862 5768 21914
rect 5768 21862 5820 21914
rect 5820 21862 6376 21914
rect 5195 21798 5251 21854
rect 5276 21798 5332 21854
rect 5357 21798 5413 21854
rect 5438 21798 5494 21854
rect 5519 21798 5575 21854
rect 5600 21850 6376 21862
rect 5600 21798 5632 21850
rect 5632 21798 5684 21850
rect 5684 21798 5700 21850
rect 5700 21798 5752 21850
rect 5752 21798 5768 21850
rect 5768 21798 5820 21850
rect 5820 21798 6376 21850
rect 5600 21786 6376 21798
rect 5195 21718 5251 21774
rect 5276 21718 5332 21774
rect 5357 21718 5413 21774
rect 5438 21718 5494 21774
rect 5519 21718 5575 21774
rect 5600 21734 5632 21786
rect 5632 21734 5684 21786
rect 5684 21734 5700 21786
rect 5700 21734 5752 21786
rect 5752 21734 5768 21786
rect 5768 21734 5820 21786
rect 5820 21734 6376 21786
rect 5600 21722 6376 21734
rect 5195 21638 5251 21694
rect 5276 21638 5332 21694
rect 5357 21638 5413 21694
rect 5438 21638 5494 21694
rect 5519 21638 5575 21694
rect 5600 21670 5632 21722
rect 5632 21670 5684 21722
rect 5684 21670 5700 21722
rect 5700 21670 5752 21722
rect 5752 21670 5768 21722
rect 5768 21670 5820 21722
rect 5820 21670 6376 21722
rect 5600 21658 6376 21670
rect 5195 21558 5251 21614
rect 5276 21558 5332 21614
rect 5357 21558 5413 21614
rect 5438 21558 5494 21614
rect 5519 21558 5575 21614
rect 5600 21606 5632 21658
rect 5632 21606 5684 21658
rect 5684 21606 5700 21658
rect 5700 21606 5752 21658
rect 5752 21606 5768 21658
rect 5768 21606 5820 21658
rect 5820 21606 6376 21658
rect 5600 21594 6376 21606
rect 5600 21542 5632 21594
rect 5632 21542 5684 21594
rect 5684 21542 5700 21594
rect 5700 21542 5752 21594
rect 5752 21542 5768 21594
rect 5768 21542 5820 21594
rect 5820 21542 6376 21594
rect 5195 21478 5251 21534
rect 5276 21478 5332 21534
rect 5357 21478 5413 21534
rect 5438 21478 5494 21534
rect 5519 21478 5575 21534
rect 5600 21529 6376 21542
rect 5600 21477 5632 21529
rect 5632 21477 5684 21529
rect 5684 21477 5700 21529
rect 5700 21477 5752 21529
rect 5752 21477 5768 21529
rect 5768 21477 5820 21529
rect 5820 21477 6376 21529
rect 5600 21464 6376 21477
rect 5195 21398 5251 21454
rect 5276 21398 5332 21454
rect 5357 21398 5413 21454
rect 5438 21398 5494 21454
rect 5519 21398 5575 21454
rect 5600 21412 5632 21464
rect 5632 21412 5684 21464
rect 5684 21412 5700 21464
rect 5700 21412 5752 21464
rect 5752 21412 5768 21464
rect 5768 21412 5820 21464
rect 5820 21412 6376 21464
rect 5600 21399 6376 21412
rect 5195 21318 5251 21374
rect 5276 21318 5332 21374
rect 5357 21318 5413 21374
rect 5438 21318 5494 21374
rect 5519 21318 5575 21374
rect 5600 21347 5632 21399
rect 5632 21347 5684 21399
rect 5684 21347 5700 21399
rect 5700 21347 5752 21399
rect 5752 21347 5768 21399
rect 5768 21347 5820 21399
rect 5820 21347 6376 21399
rect 5600 21334 6376 21347
rect 5195 21238 5251 21294
rect 5276 21238 5332 21294
rect 5357 21238 5413 21294
rect 5438 21238 5494 21294
rect 5519 21238 5575 21294
rect 5600 21282 5632 21334
rect 5632 21282 5684 21334
rect 5684 21282 5700 21334
rect 5700 21282 5752 21334
rect 5752 21282 5768 21334
rect 5768 21282 5820 21334
rect 5820 21282 6376 21334
rect 5600 21269 6376 21282
rect 5600 21217 5632 21269
rect 5632 21217 5684 21269
rect 5684 21217 5700 21269
rect 5700 21217 5752 21269
rect 5752 21217 5768 21269
rect 5768 21217 5820 21269
rect 5820 21217 6376 21269
rect 5195 21158 5251 21214
rect 5276 21158 5332 21214
rect 5357 21158 5413 21214
rect 5438 21158 5494 21214
rect 5519 21158 5575 21214
rect 5600 21204 6376 21217
rect 5600 21152 5632 21204
rect 5632 21152 5684 21204
rect 5684 21152 5700 21204
rect 5700 21152 5752 21204
rect 5752 21152 5768 21204
rect 5768 21152 5820 21204
rect 5820 21152 6376 21204
rect 5600 21139 6376 21152
rect 5195 21078 5251 21134
rect 5276 21078 5332 21134
rect 5357 21078 5413 21134
rect 5438 21078 5494 21134
rect 5519 21078 5575 21134
rect 5600 21087 5632 21139
rect 5632 21087 5684 21139
rect 5684 21087 5700 21139
rect 5700 21087 5752 21139
rect 5752 21087 5768 21139
rect 5768 21087 5820 21139
rect 5820 21087 6376 21139
rect 5600 21074 6376 21087
rect 5195 20998 5251 21054
rect 5276 20998 5332 21054
rect 5357 20998 5413 21054
rect 5438 20998 5494 21054
rect 5519 20998 5575 21054
rect 5600 21022 5632 21074
rect 5632 21022 5684 21074
rect 5684 21022 5700 21074
rect 5700 21022 5752 21074
rect 5752 21022 5768 21074
rect 5768 21022 5820 21074
rect 5820 21022 6376 21074
rect 5600 21009 6376 21022
rect 5195 20918 5251 20974
rect 5276 20918 5332 20974
rect 5357 20918 5413 20974
rect 5438 20918 5494 20974
rect 5519 20918 5575 20974
rect 5600 20957 5632 21009
rect 5632 20957 5684 21009
rect 5684 20957 5700 21009
rect 5700 20957 5752 21009
rect 5752 20957 5768 21009
rect 5768 20957 5820 21009
rect 5820 20957 6376 21009
rect 5600 20944 6376 20957
rect 5195 20838 5251 20894
rect 5276 20838 5332 20894
rect 5357 20838 5413 20894
rect 5438 20838 5494 20894
rect 5519 20838 5575 20894
rect 5600 20892 5632 20944
rect 5632 20892 5684 20944
rect 5684 20892 5700 20944
rect 5700 20892 5752 20944
rect 5752 20892 5768 20944
rect 5768 20892 5820 20944
rect 5820 20892 6376 20944
rect 5600 20879 6376 20892
rect 5600 20827 5632 20879
rect 5632 20827 5684 20879
rect 5684 20827 5700 20879
rect 5700 20827 5752 20879
rect 5752 20827 5768 20879
rect 5768 20827 5820 20879
rect 5820 20827 6376 20879
rect 5600 20814 6376 20827
rect 5195 20758 5251 20814
rect 5276 20758 5332 20814
rect 5357 20758 5413 20814
rect 5438 20758 5494 20814
rect 5519 20758 5575 20814
rect 5600 20762 5632 20814
rect 5632 20762 5684 20814
rect 5684 20762 5700 20814
rect 5700 20762 5752 20814
rect 5752 20762 5768 20814
rect 5768 20762 5820 20814
rect 5820 20762 6376 20814
rect 5600 20758 6376 20762
rect 7640 20373 7696 20429
rect 7726 20373 7782 20429
rect 7812 20373 7868 20429
rect 7898 20373 7954 20429
rect 7984 20425 8040 20429
rect 8070 20425 8126 20429
rect 7984 20373 8013 20425
rect 8013 20373 8039 20425
rect 8039 20373 8040 20425
rect 8070 20373 8091 20425
rect 8091 20373 8126 20425
rect 8156 20373 8212 20429
rect 8242 20373 8298 20429
rect 8327 20373 8383 20429
rect 8412 20373 8468 20429
rect 8497 20373 8553 20429
rect 9079 20373 9135 20429
rect 9170 20373 9226 20429
rect 9260 20373 9316 20429
rect 9350 20373 9406 20429
rect 9440 20373 9496 20429
rect 9530 20373 9586 20429
rect 9620 20373 9676 20429
rect 9710 20373 9766 20429
rect 7640 20293 7696 20349
rect 7726 20293 7782 20349
rect 7812 20293 7868 20349
rect 7898 20293 7954 20349
rect 7984 20309 8013 20349
rect 8013 20309 8039 20349
rect 8039 20309 8040 20349
rect 8070 20309 8091 20349
rect 8091 20309 8126 20349
rect 7984 20297 8040 20309
rect 8070 20297 8126 20309
rect 7984 20293 8013 20297
rect 8013 20293 8039 20297
rect 8039 20293 8040 20297
rect 8070 20293 8091 20297
rect 8091 20293 8126 20297
rect 8156 20293 8212 20349
rect 8242 20293 8298 20349
rect 8327 20293 8383 20349
rect 8412 20293 8468 20349
rect 8497 20293 8553 20349
rect 7640 20213 7696 20269
rect 7726 20213 7782 20269
rect 7812 20213 7868 20269
rect 7898 20213 7954 20269
rect 7984 20245 8013 20269
rect 8013 20245 8039 20269
rect 8039 20245 8040 20269
rect 8070 20245 8091 20269
rect 8091 20245 8126 20269
rect 7984 20233 8040 20245
rect 8070 20233 8126 20245
rect 7984 20213 8013 20233
rect 8013 20213 8039 20233
rect 8039 20213 8040 20233
rect 8070 20213 8091 20233
rect 8091 20213 8126 20233
rect 8156 20213 8212 20269
rect 8242 20213 8298 20269
rect 8327 20213 8383 20269
rect 8412 20213 8468 20269
rect 8497 20213 8553 20269
rect 9079 20293 9135 20349
rect 9170 20293 9226 20349
rect 9260 20293 9316 20349
rect 9350 20293 9406 20349
rect 9440 20293 9496 20349
rect 9530 20293 9586 20349
rect 9620 20293 9676 20349
rect 9710 20293 9766 20349
rect 7640 20133 7696 20189
rect 7726 20133 7782 20189
rect 7812 20133 7868 20189
rect 7898 20133 7954 20189
rect 7984 20181 8013 20189
rect 8013 20181 8039 20189
rect 8039 20181 8040 20189
rect 8070 20181 8091 20189
rect 8091 20181 8126 20189
rect 7984 20169 8040 20181
rect 8070 20169 8126 20181
rect 7984 20133 8013 20169
rect 8013 20133 8039 20169
rect 8039 20133 8040 20169
rect 8070 20133 8091 20169
rect 8091 20133 8126 20169
rect 8156 20133 8212 20189
rect 8242 20133 8298 20189
rect 8327 20133 8383 20189
rect 8412 20133 8468 20189
rect 8497 20133 8553 20189
rect 9079 20213 9135 20269
rect 9170 20213 9226 20269
rect 9260 20213 9316 20269
rect 9350 20213 9406 20269
rect 9440 20213 9496 20269
rect 9530 20213 9586 20269
rect 9620 20213 9676 20269
rect 9710 20213 9766 20269
rect 9079 20133 9135 20189
rect 9170 20133 9226 20189
rect 9260 20133 9316 20189
rect 9350 20133 9406 20189
rect 9440 20133 9496 20189
rect 9530 20133 9586 20189
rect 9620 20133 9676 20189
rect 9710 20133 9766 20189
rect 7640 20053 7696 20109
rect 7726 20053 7782 20109
rect 7812 20053 7868 20109
rect 7898 20053 7954 20109
rect 7984 20105 8040 20109
rect 8070 20105 8126 20109
rect 7984 20053 8013 20105
rect 8013 20053 8039 20105
rect 8039 20053 8040 20105
rect 8070 20053 8091 20105
rect 8091 20053 8126 20105
rect 8156 20053 8212 20109
rect 8242 20053 8298 20109
rect 8327 20053 8383 20109
rect 8412 20053 8468 20109
rect 8497 20053 8553 20109
rect 9079 20053 9135 20109
rect 9170 20053 9226 20109
rect 9260 20053 9316 20109
rect 9350 20053 9406 20109
rect 9440 20053 9496 20109
rect 9530 20053 9586 20109
rect 9620 20053 9676 20109
rect 9710 20053 9766 20109
rect 7640 19973 7696 20029
rect 7726 19973 7782 20029
rect 7812 19973 7868 20029
rect 7898 19973 7954 20029
rect 7984 19989 8013 20029
rect 8013 19989 8039 20029
rect 8039 19989 8040 20029
rect 8070 19989 8091 20029
rect 8091 19989 8126 20029
rect 7984 19977 8040 19989
rect 8070 19977 8126 19989
rect 7984 19973 8013 19977
rect 8013 19973 8039 19977
rect 8039 19973 8040 19977
rect 8070 19973 8091 19977
rect 8091 19973 8126 19977
rect 8156 19973 8212 20029
rect 8242 19973 8298 20029
rect 8327 19973 8383 20029
rect 8412 19973 8468 20029
rect 8497 19973 8553 20029
rect 7640 19893 7696 19949
rect 7726 19893 7782 19949
rect 7812 19893 7868 19949
rect 7898 19893 7954 19949
rect 7984 19925 8013 19949
rect 8013 19925 8039 19949
rect 8039 19925 8040 19949
rect 8070 19925 8091 19949
rect 8091 19925 8126 19949
rect 7984 19913 8040 19925
rect 8070 19913 8126 19925
rect 7984 19893 8013 19913
rect 8013 19893 8039 19913
rect 8039 19893 8040 19913
rect 8070 19893 8091 19913
rect 8091 19893 8126 19913
rect 8156 19893 8212 19949
rect 8242 19893 8298 19949
rect 8327 19893 8383 19949
rect 8412 19893 8468 19949
rect 8497 19893 8553 19949
rect 9079 19973 9135 20029
rect 9170 19973 9226 20029
rect 9260 19973 9316 20029
rect 9350 19973 9406 20029
rect 9440 19973 9496 20029
rect 9530 19973 9586 20029
rect 9620 19973 9676 20029
rect 9710 19973 9766 20029
rect 7640 19813 7696 19869
rect 7726 19813 7782 19869
rect 7812 19813 7868 19869
rect 7898 19813 7954 19869
rect 7984 19861 8013 19869
rect 8013 19861 8039 19869
rect 8039 19861 8040 19869
rect 8070 19861 8091 19869
rect 8091 19861 8126 19869
rect 7984 19849 8040 19861
rect 8070 19849 8126 19861
rect 7984 19813 8013 19849
rect 8013 19813 8039 19849
rect 8039 19813 8040 19849
rect 8070 19813 8091 19849
rect 8091 19813 8126 19849
rect 8156 19813 8212 19869
rect 8242 19813 8298 19869
rect 8327 19813 8383 19869
rect 8412 19813 8468 19869
rect 8497 19813 8553 19869
rect 9079 19893 9135 19949
rect 9170 19893 9226 19949
rect 9260 19893 9316 19949
rect 9350 19893 9406 19949
rect 9440 19893 9496 19949
rect 9530 19893 9586 19949
rect 9620 19893 9676 19949
rect 9710 19893 9766 19949
rect 9079 19813 9135 19869
rect 9170 19813 9226 19869
rect 9260 19813 9316 19869
rect 9350 19813 9406 19869
rect 9440 19813 9496 19869
rect 9530 19813 9586 19869
rect 9620 19813 9676 19869
rect 9710 19813 9766 19869
rect 7640 19733 7696 19789
rect 7726 19733 7782 19789
rect 7812 19733 7868 19789
rect 7898 19733 7954 19789
rect 7984 19785 8040 19789
rect 8070 19785 8126 19789
rect 7984 19733 8013 19785
rect 8013 19733 8039 19785
rect 8039 19733 8040 19785
rect 8070 19733 8091 19785
rect 8091 19733 8126 19785
rect 8156 19733 8212 19789
rect 8242 19733 8298 19789
rect 8327 19733 8383 19789
rect 8412 19733 8468 19789
rect 8497 19733 8553 19789
rect 9079 19733 9135 19789
rect 9170 19733 9226 19789
rect 9260 19733 9316 19789
rect 9350 19733 9406 19789
rect 9440 19733 9496 19789
rect 9530 19733 9586 19789
rect 9620 19733 9676 19789
rect 9710 19733 9766 19789
rect 7640 19653 7696 19709
rect 7726 19653 7782 19709
rect 7812 19653 7868 19709
rect 7898 19653 7954 19709
rect 7984 19669 8013 19709
rect 8013 19669 8039 19709
rect 8039 19669 8040 19709
rect 8070 19669 8091 19709
rect 8091 19669 8126 19709
rect 7984 19657 8040 19669
rect 8070 19657 8126 19669
rect 7984 19653 8013 19657
rect 8013 19653 8039 19657
rect 8039 19653 8040 19657
rect 8070 19653 8091 19657
rect 8091 19653 8126 19657
rect 8156 19653 8212 19709
rect 8242 19653 8298 19709
rect 8327 19653 8383 19709
rect 8412 19653 8468 19709
rect 8497 19653 8553 19709
rect 7640 19573 7696 19629
rect 7726 19573 7782 19629
rect 7812 19573 7868 19629
rect 7898 19573 7954 19629
rect 7984 19605 8013 19629
rect 8013 19605 8039 19629
rect 8039 19605 8040 19629
rect 8070 19605 8091 19629
rect 8091 19605 8126 19629
rect 7984 19593 8040 19605
rect 8070 19593 8126 19605
rect 7984 19573 8013 19593
rect 8013 19573 8039 19593
rect 8039 19573 8040 19593
rect 8070 19573 8091 19593
rect 8091 19573 8126 19593
rect 8156 19573 8212 19629
rect 8242 19573 8298 19629
rect 8327 19573 8383 19629
rect 8412 19573 8468 19629
rect 8497 19573 8553 19629
rect 9079 19653 9135 19709
rect 9170 19653 9226 19709
rect 9260 19653 9316 19709
rect 9350 19653 9406 19709
rect 9440 19653 9496 19709
rect 9530 19653 9586 19709
rect 9620 19653 9676 19709
rect 9710 19653 9766 19709
rect 7640 19493 7696 19549
rect 7726 19493 7782 19549
rect 7812 19493 7868 19549
rect 7898 19493 7954 19549
rect 7984 19541 8013 19549
rect 8013 19541 8039 19549
rect 8039 19541 8040 19549
rect 8070 19541 8091 19549
rect 8091 19541 8126 19549
rect 7984 19529 8040 19541
rect 8070 19529 8126 19541
rect 7984 19493 8013 19529
rect 8013 19493 8039 19529
rect 8039 19493 8040 19529
rect 8070 19493 8091 19529
rect 8091 19493 8126 19529
rect 8156 19493 8212 19549
rect 8242 19493 8298 19549
rect 8327 19493 8383 19549
rect 8412 19493 8468 19549
rect 8497 19493 8553 19549
rect 9079 19573 9135 19629
rect 9170 19573 9226 19629
rect 9260 19573 9316 19629
rect 9350 19573 9406 19629
rect 9440 19573 9496 19629
rect 9530 19573 9586 19629
rect 9620 19573 9676 19629
rect 9710 19573 9766 19629
rect 9079 19493 9135 19549
rect 9170 19493 9226 19549
rect 9260 19493 9316 19549
rect 9350 19493 9406 19549
rect 9440 19493 9496 19549
rect 9530 19493 9586 19549
rect 9620 19493 9676 19549
rect 9710 19493 9766 19549
rect 7640 19413 7696 19469
rect 7726 19413 7782 19469
rect 7812 19413 7868 19469
rect 7898 19413 7954 19469
rect 7984 19464 8040 19469
rect 8070 19464 8126 19469
rect 7984 19413 8013 19464
rect 8013 19413 8039 19464
rect 8039 19413 8040 19464
rect 8070 19413 8091 19464
rect 8091 19413 8126 19464
rect 8156 19413 8212 19469
rect 8242 19413 8298 19469
rect 8327 19413 8383 19469
rect 8412 19413 8468 19469
rect 8497 19413 8553 19469
rect 9079 19413 9135 19469
rect 9170 19413 9226 19469
rect 9260 19413 9316 19469
rect 9350 19413 9406 19469
rect 9440 19413 9496 19469
rect 9530 19413 9586 19469
rect 9620 19413 9676 19469
rect 9710 19413 9766 19469
rect 7640 19333 7696 19389
rect 7726 19333 7782 19389
rect 7812 19333 7868 19389
rect 7898 19333 7954 19389
rect 7984 19347 8013 19389
rect 8013 19347 8039 19389
rect 8039 19347 8040 19389
rect 8070 19347 8091 19389
rect 8091 19347 8126 19389
rect 7984 19334 8040 19347
rect 8070 19334 8126 19347
rect 7984 19333 8013 19334
rect 8013 19333 8039 19334
rect 8039 19333 8040 19334
rect 8070 19333 8091 19334
rect 8091 19333 8126 19334
rect 8156 19333 8212 19389
rect 8242 19333 8298 19389
rect 8327 19333 8383 19389
rect 8412 19333 8468 19389
rect 8497 19333 8553 19389
rect 7640 19253 7696 19309
rect 7726 19253 7782 19309
rect 7812 19253 7868 19309
rect 7898 19253 7954 19309
rect 7984 19282 8013 19309
rect 8013 19282 8039 19309
rect 8039 19282 8040 19309
rect 8070 19282 8091 19309
rect 8091 19282 8126 19309
rect 7984 19269 8040 19282
rect 8070 19269 8126 19282
rect 7984 19253 8013 19269
rect 8013 19253 8039 19269
rect 8039 19253 8040 19269
rect 8070 19253 8091 19269
rect 8091 19253 8126 19269
rect 8156 19253 8212 19309
rect 8242 19253 8298 19309
rect 8327 19253 8383 19309
rect 8412 19253 8468 19309
rect 8497 19253 8553 19309
rect 9079 19333 9135 19389
rect 9170 19333 9226 19389
rect 9260 19333 9316 19389
rect 9350 19333 9406 19389
rect 9440 19333 9496 19389
rect 9530 19333 9586 19389
rect 9620 19333 9676 19389
rect 9710 19333 9766 19389
rect 7640 19173 7696 19229
rect 7726 19173 7782 19229
rect 7812 19173 7868 19229
rect 7898 19173 7954 19229
rect 7984 19217 8013 19229
rect 8013 19217 8039 19229
rect 8039 19217 8040 19229
rect 8070 19217 8091 19229
rect 8091 19217 8126 19229
rect 7984 19204 8040 19217
rect 8070 19204 8126 19217
rect 7984 19173 8013 19204
rect 8013 19173 8039 19204
rect 8039 19173 8040 19204
rect 8070 19173 8091 19204
rect 8091 19173 8126 19204
rect 8156 19173 8212 19229
rect 8242 19173 8298 19229
rect 8327 19173 8383 19229
rect 8412 19173 8468 19229
rect 8497 19173 8553 19229
rect 9079 19253 9135 19309
rect 9170 19253 9226 19309
rect 9260 19253 9316 19309
rect 9350 19253 9406 19309
rect 9440 19253 9496 19309
rect 9530 19253 9586 19309
rect 9620 19253 9676 19309
rect 9710 19253 9766 19309
rect 9079 19173 9135 19229
rect 9170 19173 9226 19229
rect 9260 19173 9316 19229
rect 9350 19173 9406 19229
rect 9440 19173 9496 19229
rect 9530 19173 9586 19229
rect 9620 19173 9676 19229
rect 9710 19173 9766 19229
rect 7640 19093 7696 19149
rect 7726 19093 7782 19149
rect 7812 19093 7868 19149
rect 7898 19093 7954 19149
rect 7984 19139 8040 19149
rect 8070 19139 8126 19149
rect 7984 19093 8013 19139
rect 8013 19093 8039 19139
rect 8039 19093 8040 19139
rect 8070 19093 8091 19139
rect 8091 19093 8126 19139
rect 8156 19093 8212 19149
rect 8242 19093 8298 19149
rect 8327 19093 8383 19149
rect 8412 19093 8468 19149
rect 8497 19093 8553 19149
rect 9079 19093 9135 19149
rect 9170 19093 9226 19149
rect 9260 19093 9316 19149
rect 9350 19093 9406 19149
rect 9440 19093 9496 19149
rect 9530 19093 9586 19149
rect 9620 19093 9676 19149
rect 9710 19093 9766 19149
rect 7640 19013 7696 19069
rect 7726 19013 7782 19069
rect 7812 19013 7868 19069
rect 7898 19013 7954 19069
rect 7984 19022 8013 19069
rect 8013 19022 8039 19069
rect 8039 19022 8040 19069
rect 8070 19022 8091 19069
rect 8091 19022 8126 19069
rect 7984 19013 8040 19022
rect 8070 19013 8126 19022
rect 8156 19013 8212 19069
rect 8242 19013 8298 19069
rect 8327 19013 8383 19069
rect 8412 19013 8468 19069
rect 8497 19013 8553 19069
rect 9079 19013 9135 19069
rect 9170 19013 9226 19069
rect 9260 19013 9316 19069
rect 9350 19013 9406 19069
rect 9440 19013 9496 19069
rect 9530 19013 9586 19069
rect 9620 19013 9676 19069
rect 9710 19013 9766 19069
rect 7640 18933 7696 18989
rect 7726 18933 7782 18989
rect 7812 18933 7868 18989
rect 7898 18933 7954 18989
rect 7984 18957 8013 18989
rect 8013 18957 8039 18989
rect 8039 18957 8040 18989
rect 8070 18957 8091 18989
rect 8091 18957 8126 18989
rect 7984 18944 8040 18957
rect 8070 18944 8126 18957
rect 7984 18933 8013 18944
rect 8013 18933 8039 18944
rect 8039 18933 8040 18944
rect 8070 18933 8091 18944
rect 8091 18933 8126 18944
rect 8156 18933 8212 18989
rect 8242 18933 8298 18989
rect 8327 18933 8383 18989
rect 8412 18933 8468 18989
rect 8497 18933 8553 18989
rect 7640 18853 7696 18909
rect 7726 18853 7782 18909
rect 7812 18853 7868 18909
rect 7898 18853 7954 18909
rect 7984 18892 8013 18909
rect 8013 18892 8039 18909
rect 8039 18892 8040 18909
rect 8070 18892 8091 18909
rect 8091 18892 8126 18909
rect 7984 18879 8040 18892
rect 8070 18879 8126 18892
rect 7984 18853 8013 18879
rect 8013 18853 8039 18879
rect 8039 18853 8040 18879
rect 8070 18853 8091 18879
rect 8091 18853 8126 18879
rect 8156 18853 8212 18909
rect 8242 18853 8298 18909
rect 8327 18853 8383 18909
rect 8412 18853 8468 18909
rect 8497 18853 8553 18909
rect 9079 18933 9135 18989
rect 9170 18933 9226 18989
rect 9260 18933 9316 18989
rect 9350 18933 9406 18989
rect 9440 18933 9496 18989
rect 9530 18933 9586 18989
rect 9620 18933 9676 18989
rect 9710 18933 9766 18989
rect 7640 18773 7696 18829
rect 7726 18773 7782 18829
rect 7812 18773 7868 18829
rect 7898 18773 7954 18829
rect 7984 18827 8013 18829
rect 8013 18827 8039 18829
rect 8039 18827 8040 18829
rect 8070 18827 8091 18829
rect 8091 18827 8126 18829
rect 7984 18814 8040 18827
rect 8070 18814 8126 18827
rect 7984 18773 8013 18814
rect 8013 18773 8039 18814
rect 8039 18773 8040 18814
rect 8070 18773 8091 18814
rect 8091 18773 8126 18814
rect 8156 18773 8212 18829
rect 8242 18773 8298 18829
rect 8327 18773 8383 18829
rect 8412 18773 8468 18829
rect 8497 18773 8553 18829
rect 9079 18853 9135 18909
rect 9170 18853 9226 18909
rect 9260 18853 9316 18909
rect 9350 18853 9406 18909
rect 9440 18853 9496 18909
rect 9530 18853 9586 18909
rect 9620 18853 9676 18909
rect 9710 18853 9766 18909
rect 9079 18773 9135 18829
rect 9170 18773 9226 18829
rect 9260 18773 9316 18829
rect 9350 18773 9406 18829
rect 9440 18773 9496 18829
rect 9530 18773 9586 18829
rect 9620 18773 9676 18829
rect 9710 18773 9766 18829
rect 7640 18693 7696 18749
rect 7726 18693 7782 18749
rect 7812 18693 7868 18749
rect 7898 18693 7954 18749
rect 7984 18697 8013 18749
rect 8013 18697 8039 18749
rect 8039 18697 8040 18749
rect 8070 18697 8091 18749
rect 8091 18697 8126 18749
rect 7984 18693 8040 18697
rect 8070 18693 8126 18697
rect 8156 18693 8212 18749
rect 8242 18693 8298 18749
rect 8327 18693 8383 18749
rect 8412 18693 8468 18749
rect 8497 18693 8553 18749
rect 9079 18693 9135 18749
rect 9170 18693 9226 18749
rect 9260 18693 9316 18749
rect 9350 18693 9406 18749
rect 9440 18693 9496 18749
rect 9530 18693 9586 18749
rect 9620 18693 9676 18749
rect 9710 18693 9766 18749
rect 5188 17838 5244 17894
rect 5270 17838 5326 17894
rect 5352 17838 5408 17894
rect 5434 17838 5490 17894
rect 5516 17838 5572 17894
rect 5598 17890 5654 17894
rect 5680 17890 5736 17894
rect 5762 17890 5818 17894
rect 5598 17838 5632 17890
rect 5632 17838 5654 17890
rect 5680 17838 5684 17890
rect 5684 17838 5700 17890
rect 5700 17838 5736 17890
rect 5762 17838 5768 17890
rect 5768 17838 5818 17890
rect 5844 17838 5900 17894
rect 5926 17838 5982 17894
rect 6008 17838 6064 17894
rect 6090 17838 6146 17894
rect 6172 17838 6228 17894
rect 6254 17838 6310 17894
rect 6336 17838 6392 17894
rect 6418 17838 6474 17894
rect 6500 17890 6556 17894
rect 6582 17890 6638 17894
rect 6664 17890 6720 17894
rect 6500 17838 6552 17890
rect 6552 17838 6556 17890
rect 6582 17838 6604 17890
rect 6604 17838 6620 17890
rect 6620 17838 6638 17890
rect 6664 17838 6672 17890
rect 6672 17838 6688 17890
rect 6688 17838 6720 17890
rect 6746 17838 6802 17894
rect 6828 17838 6884 17894
rect 6909 17838 6965 17894
rect 6990 17838 7046 17894
rect 7071 17838 7127 17894
rect 7152 17838 7208 17894
rect 7233 17838 7289 17894
rect 7314 17838 7370 17894
rect 5188 17758 5244 17814
rect 5270 17758 5326 17814
rect 5352 17758 5408 17814
rect 5434 17758 5490 17814
rect 5516 17758 5572 17814
rect 5598 17774 5632 17814
rect 5632 17774 5654 17814
rect 5680 17774 5684 17814
rect 5684 17774 5700 17814
rect 5700 17774 5736 17814
rect 5762 17774 5768 17814
rect 5768 17774 5818 17814
rect 5598 17762 5654 17774
rect 5680 17762 5736 17774
rect 5762 17762 5818 17774
rect 5598 17758 5632 17762
rect 5632 17758 5654 17762
rect 5680 17758 5684 17762
rect 5684 17758 5700 17762
rect 5700 17758 5736 17762
rect 5762 17758 5768 17762
rect 5768 17758 5818 17762
rect 5844 17758 5900 17814
rect 5926 17758 5982 17814
rect 6008 17758 6064 17814
rect 6090 17758 6146 17814
rect 6172 17758 6228 17814
rect 6254 17758 6310 17814
rect 6336 17758 6392 17814
rect 6418 17758 6474 17814
rect 6500 17774 6552 17814
rect 6552 17774 6556 17814
rect 6582 17774 6604 17814
rect 6604 17774 6620 17814
rect 6620 17774 6638 17814
rect 6664 17774 6672 17814
rect 6672 17774 6688 17814
rect 6688 17774 6720 17814
rect 6500 17762 6556 17774
rect 6582 17762 6638 17774
rect 6664 17762 6720 17774
rect 6500 17758 6552 17762
rect 6552 17758 6556 17762
rect 6582 17758 6604 17762
rect 6604 17758 6620 17762
rect 6620 17758 6638 17762
rect 6664 17758 6672 17762
rect 6672 17758 6688 17762
rect 6688 17758 6720 17762
rect 6746 17758 6802 17814
rect 6828 17758 6884 17814
rect 6909 17758 6965 17814
rect 6990 17758 7046 17814
rect 7071 17758 7127 17814
rect 7152 17758 7208 17814
rect 7233 17758 7289 17814
rect 7314 17758 7370 17814
rect 5188 17678 5244 17734
rect 5270 17678 5326 17734
rect 5352 17678 5408 17734
rect 5434 17678 5490 17734
rect 5516 17678 5572 17734
rect 5598 17710 5632 17734
rect 5632 17710 5654 17734
rect 5680 17710 5684 17734
rect 5684 17710 5700 17734
rect 5700 17710 5736 17734
rect 5762 17710 5768 17734
rect 5768 17710 5818 17734
rect 5598 17698 5654 17710
rect 5680 17698 5736 17710
rect 5762 17698 5818 17710
rect 5598 17678 5632 17698
rect 5632 17678 5654 17698
rect 5680 17678 5684 17698
rect 5684 17678 5700 17698
rect 5700 17678 5736 17698
rect 5762 17678 5768 17698
rect 5768 17678 5818 17698
rect 5844 17678 5900 17734
rect 5926 17678 5982 17734
rect 6008 17678 6064 17734
rect 6090 17678 6146 17734
rect 6172 17678 6228 17734
rect 6254 17678 6310 17734
rect 6336 17678 6392 17734
rect 6418 17678 6474 17734
rect 6500 17710 6552 17734
rect 6552 17710 6556 17734
rect 6582 17710 6604 17734
rect 6604 17710 6620 17734
rect 6620 17710 6638 17734
rect 6664 17710 6672 17734
rect 6672 17710 6688 17734
rect 6688 17710 6720 17734
rect 6500 17698 6556 17710
rect 6582 17698 6638 17710
rect 6664 17698 6720 17710
rect 6500 17678 6552 17698
rect 6552 17678 6556 17698
rect 6582 17678 6604 17698
rect 6604 17678 6620 17698
rect 6620 17678 6638 17698
rect 6664 17678 6672 17698
rect 6672 17678 6688 17698
rect 6688 17678 6720 17698
rect 6746 17678 6802 17734
rect 6828 17678 6884 17734
rect 6909 17678 6965 17734
rect 6990 17678 7046 17734
rect 7071 17678 7127 17734
rect 7152 17678 7208 17734
rect 7233 17678 7289 17734
rect 7314 17678 7370 17734
rect 5188 17598 5244 17654
rect 5270 17598 5326 17654
rect 5352 17598 5408 17654
rect 5434 17598 5490 17654
rect 5516 17598 5572 17654
rect 5598 17646 5632 17654
rect 5632 17646 5654 17654
rect 5680 17646 5684 17654
rect 5684 17646 5700 17654
rect 5700 17646 5736 17654
rect 5762 17646 5768 17654
rect 5768 17646 5818 17654
rect 5598 17634 5654 17646
rect 5680 17634 5736 17646
rect 5762 17634 5818 17646
rect 5598 17598 5632 17634
rect 5632 17598 5654 17634
rect 5680 17598 5684 17634
rect 5684 17598 5700 17634
rect 5700 17598 5736 17634
rect 5762 17598 5768 17634
rect 5768 17598 5818 17634
rect 5844 17598 5900 17654
rect 5926 17598 5982 17654
rect 6008 17598 6064 17654
rect 6090 17598 6146 17654
rect 6172 17598 6228 17654
rect 6254 17598 6310 17654
rect 6336 17598 6392 17654
rect 6418 17598 6474 17654
rect 6500 17646 6552 17654
rect 6552 17646 6556 17654
rect 6582 17646 6604 17654
rect 6604 17646 6620 17654
rect 6620 17646 6638 17654
rect 6664 17646 6672 17654
rect 6672 17646 6688 17654
rect 6688 17646 6720 17654
rect 6500 17634 6556 17646
rect 6582 17634 6638 17646
rect 6664 17634 6720 17646
rect 6500 17598 6552 17634
rect 6552 17598 6556 17634
rect 6582 17598 6604 17634
rect 6604 17598 6620 17634
rect 6620 17598 6638 17634
rect 6664 17598 6672 17634
rect 6672 17598 6688 17634
rect 6688 17598 6720 17634
rect 6746 17598 6802 17654
rect 6828 17598 6884 17654
rect 6909 17598 6965 17654
rect 6990 17598 7046 17654
rect 7071 17598 7127 17654
rect 7152 17598 7208 17654
rect 7233 17598 7289 17654
rect 7314 17598 7370 17654
rect 5188 17518 5244 17574
rect 5270 17518 5326 17574
rect 5352 17518 5408 17574
rect 5434 17518 5490 17574
rect 5516 17518 5572 17574
rect 5598 17570 5654 17574
rect 5680 17570 5736 17574
rect 5762 17570 5818 17574
rect 5598 17518 5632 17570
rect 5632 17518 5654 17570
rect 5680 17518 5684 17570
rect 5684 17518 5700 17570
rect 5700 17518 5736 17570
rect 5762 17518 5768 17570
rect 5768 17518 5818 17570
rect 5844 17518 5900 17574
rect 5926 17518 5982 17574
rect 6008 17518 6064 17574
rect 6090 17518 6146 17574
rect 6172 17518 6228 17574
rect 6254 17518 6310 17574
rect 6336 17518 6392 17574
rect 6418 17518 6474 17574
rect 6500 17570 6556 17574
rect 6582 17570 6638 17574
rect 6664 17570 6720 17574
rect 6500 17518 6552 17570
rect 6552 17518 6556 17570
rect 6582 17518 6604 17570
rect 6604 17518 6620 17570
rect 6620 17518 6638 17570
rect 6664 17518 6672 17570
rect 6672 17518 6688 17570
rect 6688 17518 6720 17570
rect 6746 17518 6802 17574
rect 6828 17518 6884 17574
rect 6909 17518 6965 17574
rect 6990 17518 7046 17574
rect 7071 17518 7127 17574
rect 7152 17518 7208 17574
rect 7233 17518 7289 17574
rect 7314 17518 7370 17574
rect 5188 17438 5244 17494
rect 5270 17438 5326 17494
rect 5352 17438 5408 17494
rect 5434 17438 5490 17494
rect 5516 17438 5572 17494
rect 5598 17454 5632 17494
rect 5632 17454 5654 17494
rect 5680 17454 5684 17494
rect 5684 17454 5700 17494
rect 5700 17454 5736 17494
rect 5762 17454 5768 17494
rect 5768 17454 5818 17494
rect 5598 17442 5654 17454
rect 5680 17442 5736 17454
rect 5762 17442 5818 17454
rect 5598 17438 5632 17442
rect 5632 17438 5654 17442
rect 5680 17438 5684 17442
rect 5684 17438 5700 17442
rect 5700 17438 5736 17442
rect 5762 17438 5768 17442
rect 5768 17438 5818 17442
rect 5844 17438 5900 17494
rect 5926 17438 5982 17494
rect 6008 17438 6064 17494
rect 6090 17438 6146 17494
rect 6172 17438 6228 17494
rect 6254 17438 6310 17494
rect 6336 17438 6392 17494
rect 6418 17438 6474 17494
rect 6500 17454 6552 17494
rect 6552 17454 6556 17494
rect 6582 17454 6604 17494
rect 6604 17454 6620 17494
rect 6620 17454 6638 17494
rect 6664 17454 6672 17494
rect 6672 17454 6688 17494
rect 6688 17454 6720 17494
rect 6500 17442 6556 17454
rect 6582 17442 6638 17454
rect 6664 17442 6720 17454
rect 6500 17438 6552 17442
rect 6552 17438 6556 17442
rect 6582 17438 6604 17442
rect 6604 17438 6620 17442
rect 6620 17438 6638 17442
rect 6664 17438 6672 17442
rect 6672 17438 6688 17442
rect 6688 17438 6720 17442
rect 6746 17438 6802 17494
rect 6828 17438 6884 17494
rect 6909 17438 6965 17494
rect 6990 17438 7046 17494
rect 7071 17438 7127 17494
rect 7152 17438 7208 17494
rect 7233 17438 7289 17494
rect 7314 17438 7370 17494
rect 5188 17358 5244 17414
rect 5270 17358 5326 17414
rect 5352 17358 5408 17414
rect 5434 17358 5490 17414
rect 5516 17358 5572 17414
rect 5598 17390 5632 17414
rect 5632 17390 5654 17414
rect 5680 17390 5684 17414
rect 5684 17390 5700 17414
rect 5700 17390 5736 17414
rect 5762 17390 5768 17414
rect 5768 17390 5818 17414
rect 5598 17378 5654 17390
rect 5680 17378 5736 17390
rect 5762 17378 5818 17390
rect 5598 17358 5632 17378
rect 5632 17358 5654 17378
rect 5680 17358 5684 17378
rect 5684 17358 5700 17378
rect 5700 17358 5736 17378
rect 5762 17358 5768 17378
rect 5768 17358 5818 17378
rect 5844 17358 5900 17414
rect 5926 17358 5982 17414
rect 6008 17358 6064 17414
rect 6090 17358 6146 17414
rect 6172 17358 6228 17414
rect 6254 17358 6310 17414
rect 6336 17358 6392 17414
rect 6418 17358 6474 17414
rect 6500 17390 6552 17414
rect 6552 17390 6556 17414
rect 6582 17390 6604 17414
rect 6604 17390 6620 17414
rect 6620 17390 6638 17414
rect 6664 17390 6672 17414
rect 6672 17390 6688 17414
rect 6688 17390 6720 17414
rect 6500 17378 6556 17390
rect 6582 17378 6638 17390
rect 6664 17378 6720 17390
rect 6500 17358 6552 17378
rect 6552 17358 6556 17378
rect 6582 17358 6604 17378
rect 6604 17358 6620 17378
rect 6620 17358 6638 17378
rect 6664 17358 6672 17378
rect 6672 17358 6688 17378
rect 6688 17358 6720 17378
rect 6746 17358 6802 17414
rect 6828 17358 6884 17414
rect 6909 17358 6965 17414
rect 6990 17358 7046 17414
rect 7071 17358 7127 17414
rect 7152 17358 7208 17414
rect 7233 17358 7289 17414
rect 7314 17358 7370 17414
rect 5188 17278 5244 17334
rect 5270 17278 5326 17334
rect 5352 17278 5408 17334
rect 5434 17278 5490 17334
rect 5516 17278 5572 17334
rect 5598 17326 5632 17334
rect 5632 17326 5654 17334
rect 5680 17326 5684 17334
rect 5684 17326 5700 17334
rect 5700 17326 5736 17334
rect 5762 17326 5768 17334
rect 5768 17326 5818 17334
rect 5598 17314 5654 17326
rect 5680 17314 5736 17326
rect 5762 17314 5818 17326
rect 5598 17278 5632 17314
rect 5632 17278 5654 17314
rect 5680 17278 5684 17314
rect 5684 17278 5700 17314
rect 5700 17278 5736 17314
rect 5762 17278 5768 17314
rect 5768 17278 5818 17314
rect 5844 17278 5900 17334
rect 5926 17278 5982 17334
rect 6008 17278 6064 17334
rect 6090 17278 6146 17334
rect 6172 17278 6228 17334
rect 6254 17278 6310 17334
rect 6336 17278 6392 17334
rect 6418 17278 6474 17334
rect 6500 17326 6552 17334
rect 6552 17326 6556 17334
rect 6582 17326 6604 17334
rect 6604 17326 6620 17334
rect 6620 17326 6638 17334
rect 6664 17326 6672 17334
rect 6672 17326 6688 17334
rect 6688 17326 6720 17334
rect 6500 17314 6556 17326
rect 6582 17314 6638 17326
rect 6664 17314 6720 17326
rect 6500 17278 6552 17314
rect 6552 17278 6556 17314
rect 6582 17278 6604 17314
rect 6604 17278 6620 17314
rect 6620 17278 6638 17314
rect 6664 17278 6672 17314
rect 6672 17278 6688 17314
rect 6688 17278 6720 17314
rect 6746 17278 6802 17334
rect 6828 17278 6884 17334
rect 6909 17278 6965 17334
rect 6990 17278 7046 17334
rect 7071 17278 7127 17334
rect 7152 17278 7208 17334
rect 7233 17278 7289 17334
rect 7314 17278 7370 17334
rect 5188 17198 5244 17254
rect 5270 17198 5326 17254
rect 5352 17198 5408 17254
rect 5434 17198 5490 17254
rect 5516 17198 5572 17254
rect 5598 17250 5654 17254
rect 5680 17250 5736 17254
rect 5762 17250 5818 17254
rect 5598 17198 5632 17250
rect 5632 17198 5654 17250
rect 5680 17198 5684 17250
rect 5684 17198 5700 17250
rect 5700 17198 5736 17250
rect 5762 17198 5768 17250
rect 5768 17198 5818 17250
rect 5844 17198 5900 17254
rect 5926 17198 5982 17254
rect 6008 17198 6064 17254
rect 6090 17198 6146 17254
rect 6172 17198 6228 17254
rect 6254 17198 6310 17254
rect 6336 17198 6392 17254
rect 6418 17198 6474 17254
rect 6500 17250 6556 17254
rect 6582 17250 6638 17254
rect 6664 17250 6720 17254
rect 6500 17198 6552 17250
rect 6552 17198 6556 17250
rect 6582 17198 6604 17250
rect 6604 17198 6620 17250
rect 6620 17198 6638 17250
rect 6664 17198 6672 17250
rect 6672 17198 6688 17250
rect 6688 17198 6720 17250
rect 6746 17198 6802 17254
rect 6828 17198 6884 17254
rect 6909 17198 6965 17254
rect 6990 17198 7046 17254
rect 7071 17198 7127 17254
rect 7152 17198 7208 17254
rect 7233 17198 7289 17254
rect 7314 17198 7370 17254
rect 5188 17118 5244 17174
rect 5270 17118 5326 17174
rect 5352 17118 5408 17174
rect 5434 17118 5490 17174
rect 5516 17118 5572 17174
rect 5598 17134 5632 17174
rect 5632 17134 5654 17174
rect 5680 17134 5684 17174
rect 5684 17134 5700 17174
rect 5700 17134 5736 17174
rect 5762 17134 5768 17174
rect 5768 17134 5818 17174
rect 5598 17122 5654 17134
rect 5680 17122 5736 17134
rect 5762 17122 5818 17134
rect 5598 17118 5632 17122
rect 5632 17118 5654 17122
rect 5680 17118 5684 17122
rect 5684 17118 5700 17122
rect 5700 17118 5736 17122
rect 5762 17118 5768 17122
rect 5768 17118 5818 17122
rect 5844 17118 5900 17174
rect 5926 17118 5982 17174
rect 6008 17118 6064 17174
rect 6090 17118 6146 17174
rect 6172 17118 6228 17174
rect 6254 17118 6310 17174
rect 6336 17118 6392 17174
rect 6418 17118 6474 17174
rect 6500 17134 6552 17174
rect 6552 17134 6556 17174
rect 6582 17134 6604 17174
rect 6604 17134 6620 17174
rect 6620 17134 6638 17174
rect 6664 17134 6672 17174
rect 6672 17134 6688 17174
rect 6688 17134 6720 17174
rect 6500 17122 6556 17134
rect 6582 17122 6638 17134
rect 6664 17122 6720 17134
rect 6500 17118 6552 17122
rect 6552 17118 6556 17122
rect 6582 17118 6604 17122
rect 6604 17118 6620 17122
rect 6620 17118 6638 17122
rect 6664 17118 6672 17122
rect 6672 17118 6688 17122
rect 6688 17118 6720 17122
rect 6746 17118 6802 17174
rect 6828 17118 6884 17174
rect 6909 17118 6965 17174
rect 6990 17118 7046 17174
rect 7071 17118 7127 17174
rect 7152 17118 7208 17174
rect 7233 17118 7289 17174
rect 7314 17118 7370 17174
rect 5188 17038 5244 17094
rect 5270 17038 5326 17094
rect 5352 17038 5408 17094
rect 5434 17038 5490 17094
rect 5516 17038 5572 17094
rect 5598 17070 5632 17094
rect 5632 17070 5654 17094
rect 5680 17070 5684 17094
rect 5684 17070 5700 17094
rect 5700 17070 5736 17094
rect 5762 17070 5768 17094
rect 5768 17070 5818 17094
rect 5598 17058 5654 17070
rect 5680 17058 5736 17070
rect 5762 17058 5818 17070
rect 5598 17038 5632 17058
rect 5632 17038 5654 17058
rect 5680 17038 5684 17058
rect 5684 17038 5700 17058
rect 5700 17038 5736 17058
rect 5762 17038 5768 17058
rect 5768 17038 5818 17058
rect 5844 17038 5900 17094
rect 5926 17038 5982 17094
rect 6008 17038 6064 17094
rect 6090 17038 6146 17094
rect 6172 17038 6228 17094
rect 6254 17038 6310 17094
rect 6336 17038 6392 17094
rect 6418 17038 6474 17094
rect 6500 17070 6552 17094
rect 6552 17070 6556 17094
rect 6582 17070 6604 17094
rect 6604 17070 6620 17094
rect 6620 17070 6638 17094
rect 6664 17070 6672 17094
rect 6672 17070 6688 17094
rect 6688 17070 6720 17094
rect 6500 17058 6556 17070
rect 6582 17058 6638 17070
rect 6664 17058 6720 17070
rect 6500 17038 6552 17058
rect 6552 17038 6556 17058
rect 6582 17038 6604 17058
rect 6604 17038 6620 17058
rect 6620 17038 6638 17058
rect 6664 17038 6672 17058
rect 6672 17038 6688 17058
rect 6688 17038 6720 17058
rect 6746 17038 6802 17094
rect 6828 17038 6884 17094
rect 6909 17038 6965 17094
rect 6990 17038 7046 17094
rect 7071 17038 7127 17094
rect 7152 17038 7208 17094
rect 7233 17038 7289 17094
rect 7314 17038 7370 17094
rect 5188 16958 5244 17014
rect 5270 16958 5326 17014
rect 5352 16958 5408 17014
rect 5434 16958 5490 17014
rect 5516 16958 5572 17014
rect 5598 17006 5632 17014
rect 5632 17006 5654 17014
rect 5680 17006 5684 17014
rect 5684 17006 5700 17014
rect 5700 17006 5736 17014
rect 5762 17006 5768 17014
rect 5768 17006 5818 17014
rect 5598 16994 5654 17006
rect 5680 16994 5736 17006
rect 5762 16994 5818 17006
rect 5598 16958 5632 16994
rect 5632 16958 5654 16994
rect 5680 16958 5684 16994
rect 5684 16958 5700 16994
rect 5700 16958 5736 16994
rect 5762 16958 5768 16994
rect 5768 16958 5818 16994
rect 5844 16958 5900 17014
rect 5926 16958 5982 17014
rect 6008 16958 6064 17014
rect 6090 16958 6146 17014
rect 6172 16958 6228 17014
rect 6254 16958 6310 17014
rect 6336 16958 6392 17014
rect 6418 16958 6474 17014
rect 6500 17006 6552 17014
rect 6552 17006 6556 17014
rect 6582 17006 6604 17014
rect 6604 17006 6620 17014
rect 6620 17006 6638 17014
rect 6664 17006 6672 17014
rect 6672 17006 6688 17014
rect 6688 17006 6720 17014
rect 6500 16994 6556 17006
rect 6582 16994 6638 17006
rect 6664 16994 6720 17006
rect 6500 16958 6552 16994
rect 6552 16958 6556 16994
rect 6582 16958 6604 16994
rect 6604 16958 6620 16994
rect 6620 16958 6638 16994
rect 6664 16958 6672 16994
rect 6672 16958 6688 16994
rect 6688 16958 6720 16994
rect 6746 16958 6802 17014
rect 6828 16958 6884 17014
rect 6909 16958 6965 17014
rect 6990 16958 7046 17014
rect 7071 16958 7127 17014
rect 7152 16958 7208 17014
rect 7233 16958 7289 17014
rect 7314 16958 7370 17014
rect 5188 16878 5244 16934
rect 5270 16878 5326 16934
rect 5352 16878 5408 16934
rect 5434 16878 5490 16934
rect 5516 16878 5572 16934
rect 5598 16929 5654 16934
rect 5680 16929 5736 16934
rect 5762 16929 5818 16934
rect 5598 16878 5632 16929
rect 5632 16878 5654 16929
rect 5680 16878 5684 16929
rect 5684 16878 5700 16929
rect 5700 16878 5736 16929
rect 5762 16878 5768 16929
rect 5768 16878 5818 16929
rect 5844 16878 5900 16934
rect 5926 16878 5982 16934
rect 6008 16878 6064 16934
rect 6090 16878 6146 16934
rect 6172 16878 6228 16934
rect 6254 16878 6310 16934
rect 6336 16878 6392 16934
rect 6418 16878 6474 16934
rect 6500 16929 6556 16934
rect 6582 16929 6638 16934
rect 6664 16929 6720 16934
rect 6500 16878 6552 16929
rect 6552 16878 6556 16929
rect 6582 16878 6604 16929
rect 6604 16878 6620 16929
rect 6620 16878 6638 16929
rect 6664 16878 6672 16929
rect 6672 16878 6688 16929
rect 6688 16878 6720 16929
rect 6746 16878 6802 16934
rect 6828 16878 6884 16934
rect 6909 16878 6965 16934
rect 6990 16878 7046 16934
rect 7071 16878 7127 16934
rect 7152 16878 7208 16934
rect 7233 16878 7289 16934
rect 7314 16878 7370 16934
rect 5188 16798 5244 16854
rect 5270 16798 5326 16854
rect 5352 16798 5408 16854
rect 5434 16798 5490 16854
rect 5516 16798 5572 16854
rect 5598 16812 5632 16854
rect 5632 16812 5654 16854
rect 5680 16812 5684 16854
rect 5684 16812 5700 16854
rect 5700 16812 5736 16854
rect 5762 16812 5768 16854
rect 5768 16812 5818 16854
rect 5598 16799 5654 16812
rect 5680 16799 5736 16812
rect 5762 16799 5818 16812
rect 5598 16798 5632 16799
rect 5632 16798 5654 16799
rect 5680 16798 5684 16799
rect 5684 16798 5700 16799
rect 5700 16798 5736 16799
rect 5762 16798 5768 16799
rect 5768 16798 5818 16799
rect 5844 16798 5900 16854
rect 5926 16798 5982 16854
rect 6008 16798 6064 16854
rect 6090 16798 6146 16854
rect 6172 16798 6228 16854
rect 6254 16798 6310 16854
rect 6336 16798 6392 16854
rect 6418 16798 6474 16854
rect 6500 16812 6552 16854
rect 6552 16812 6556 16854
rect 6582 16812 6604 16854
rect 6604 16812 6620 16854
rect 6620 16812 6638 16854
rect 6664 16812 6672 16854
rect 6672 16812 6688 16854
rect 6688 16812 6720 16854
rect 6500 16799 6556 16812
rect 6582 16799 6638 16812
rect 6664 16799 6720 16812
rect 6500 16798 6552 16799
rect 6552 16798 6556 16799
rect 6582 16798 6604 16799
rect 6604 16798 6620 16799
rect 6620 16798 6638 16799
rect 6664 16798 6672 16799
rect 6672 16798 6688 16799
rect 6688 16798 6720 16799
rect 6746 16798 6802 16854
rect 6828 16798 6884 16854
rect 6909 16798 6965 16854
rect 6990 16798 7046 16854
rect 7071 16798 7127 16854
rect 7152 16798 7208 16854
rect 7233 16798 7289 16854
rect 7314 16798 7370 16854
rect 5188 16718 5244 16774
rect 5270 16718 5326 16774
rect 5352 16718 5408 16774
rect 5434 16718 5490 16774
rect 5516 16718 5572 16774
rect 5598 16747 5632 16774
rect 5632 16747 5654 16774
rect 5680 16747 5684 16774
rect 5684 16747 5700 16774
rect 5700 16747 5736 16774
rect 5762 16747 5768 16774
rect 5768 16747 5818 16774
rect 5598 16734 5654 16747
rect 5680 16734 5736 16747
rect 5762 16734 5818 16747
rect 5598 16718 5632 16734
rect 5632 16718 5654 16734
rect 5680 16718 5684 16734
rect 5684 16718 5700 16734
rect 5700 16718 5736 16734
rect 5762 16718 5768 16734
rect 5768 16718 5818 16734
rect 5844 16718 5900 16774
rect 5926 16718 5982 16774
rect 6008 16718 6064 16774
rect 6090 16718 6146 16774
rect 6172 16718 6228 16774
rect 6254 16718 6310 16774
rect 6336 16718 6392 16774
rect 6418 16718 6474 16774
rect 6500 16747 6552 16774
rect 6552 16747 6556 16774
rect 6582 16747 6604 16774
rect 6604 16747 6620 16774
rect 6620 16747 6638 16774
rect 6664 16747 6672 16774
rect 6672 16747 6688 16774
rect 6688 16747 6720 16774
rect 6500 16734 6556 16747
rect 6582 16734 6638 16747
rect 6664 16734 6720 16747
rect 6500 16718 6552 16734
rect 6552 16718 6556 16734
rect 6582 16718 6604 16734
rect 6604 16718 6620 16734
rect 6620 16718 6638 16734
rect 6664 16718 6672 16734
rect 6672 16718 6688 16734
rect 6688 16718 6720 16734
rect 6746 16718 6802 16774
rect 6828 16718 6884 16774
rect 6909 16718 6965 16774
rect 6990 16718 7046 16774
rect 7071 16718 7127 16774
rect 7152 16718 7208 16774
rect 7233 16718 7289 16774
rect 7314 16718 7370 16774
rect 5188 16638 5244 16694
rect 5270 16638 5326 16694
rect 5352 16638 5408 16694
rect 5434 16638 5490 16694
rect 5516 16638 5572 16694
rect 5598 16682 5632 16694
rect 5632 16682 5654 16694
rect 5680 16682 5684 16694
rect 5684 16682 5700 16694
rect 5700 16682 5736 16694
rect 5762 16682 5768 16694
rect 5768 16682 5818 16694
rect 5598 16669 5654 16682
rect 5680 16669 5736 16682
rect 5762 16669 5818 16682
rect 5598 16638 5632 16669
rect 5632 16638 5654 16669
rect 5680 16638 5684 16669
rect 5684 16638 5700 16669
rect 5700 16638 5736 16669
rect 5762 16638 5768 16669
rect 5768 16638 5818 16669
rect 5844 16638 5900 16694
rect 5926 16638 5982 16694
rect 6008 16638 6064 16694
rect 6090 16638 6146 16694
rect 6172 16638 6228 16694
rect 6254 16638 6310 16694
rect 6336 16638 6392 16694
rect 6418 16638 6474 16694
rect 6500 16682 6552 16694
rect 6552 16682 6556 16694
rect 6582 16682 6604 16694
rect 6604 16682 6620 16694
rect 6620 16682 6638 16694
rect 6664 16682 6672 16694
rect 6672 16682 6688 16694
rect 6688 16682 6720 16694
rect 6500 16669 6556 16682
rect 6582 16669 6638 16682
rect 6664 16669 6720 16682
rect 6500 16638 6552 16669
rect 6552 16638 6556 16669
rect 6582 16638 6604 16669
rect 6604 16638 6620 16669
rect 6620 16638 6638 16669
rect 6664 16638 6672 16669
rect 6672 16638 6688 16669
rect 6688 16638 6720 16669
rect 6746 16638 6802 16694
rect 6828 16638 6884 16694
rect 6909 16638 6965 16694
rect 6990 16638 7046 16694
rect 7071 16638 7127 16694
rect 7152 16638 7208 16694
rect 7233 16638 7289 16694
rect 7314 16638 7370 16694
rect 5188 16558 5244 16614
rect 5270 16558 5326 16614
rect 5352 16558 5408 16614
rect 5434 16558 5490 16614
rect 5516 16558 5572 16614
rect 5598 16604 5654 16614
rect 5680 16604 5736 16614
rect 5762 16604 5818 16614
rect 5598 16558 5632 16604
rect 5632 16558 5654 16604
rect 5680 16558 5684 16604
rect 5684 16558 5700 16604
rect 5700 16558 5736 16604
rect 5762 16558 5768 16604
rect 5768 16558 5818 16604
rect 5844 16558 5900 16614
rect 5926 16558 5982 16614
rect 6008 16558 6064 16614
rect 6090 16558 6146 16614
rect 6172 16558 6228 16614
rect 6254 16558 6310 16614
rect 6336 16558 6392 16614
rect 6418 16558 6474 16614
rect 6500 16604 6556 16614
rect 6582 16604 6638 16614
rect 6664 16604 6720 16614
rect 6500 16558 6552 16604
rect 6552 16558 6556 16604
rect 6582 16558 6604 16604
rect 6604 16558 6620 16604
rect 6620 16558 6638 16604
rect 6664 16558 6672 16604
rect 6672 16558 6688 16604
rect 6688 16558 6720 16604
rect 6746 16558 6802 16614
rect 6828 16558 6884 16614
rect 6909 16558 6965 16614
rect 6990 16558 7046 16614
rect 7071 16558 7127 16614
rect 7152 16558 7208 16614
rect 7233 16558 7289 16614
rect 7314 16558 7370 16614
rect 5188 16478 5244 16534
rect 5270 16478 5326 16534
rect 5352 16478 5408 16534
rect 5434 16478 5490 16534
rect 5516 16478 5572 16534
rect 5598 16487 5632 16534
rect 5632 16487 5654 16534
rect 5680 16487 5684 16534
rect 5684 16487 5700 16534
rect 5700 16487 5736 16534
rect 5762 16487 5768 16534
rect 5768 16487 5818 16534
rect 5598 16478 5654 16487
rect 5680 16478 5736 16487
rect 5762 16478 5818 16487
rect 5844 16478 5900 16534
rect 5926 16478 5982 16534
rect 6008 16478 6064 16534
rect 6090 16478 6146 16534
rect 6172 16478 6228 16534
rect 6254 16478 6310 16534
rect 6336 16478 6392 16534
rect 6418 16478 6474 16534
rect 6500 16487 6552 16534
rect 6552 16487 6556 16534
rect 6582 16487 6604 16534
rect 6604 16487 6620 16534
rect 6620 16487 6638 16534
rect 6664 16487 6672 16534
rect 6672 16487 6688 16534
rect 6688 16487 6720 16534
rect 6500 16478 6556 16487
rect 6582 16478 6638 16487
rect 6664 16478 6720 16487
rect 6746 16478 6802 16534
rect 6828 16478 6884 16534
rect 6909 16478 6965 16534
rect 6990 16478 7046 16534
rect 7071 16478 7127 16534
rect 7152 16478 7208 16534
rect 7233 16478 7289 16534
rect 7314 16478 7370 16534
rect 5188 16398 5244 16454
rect 5270 16398 5326 16454
rect 5352 16398 5408 16454
rect 5434 16398 5490 16454
rect 5516 16398 5572 16454
rect 5598 16422 5632 16454
rect 5632 16422 5654 16454
rect 5680 16422 5684 16454
rect 5684 16422 5700 16454
rect 5700 16422 5736 16454
rect 5762 16422 5768 16454
rect 5768 16422 5818 16454
rect 5598 16409 5654 16422
rect 5680 16409 5736 16422
rect 5762 16409 5818 16422
rect 5598 16398 5632 16409
rect 5632 16398 5654 16409
rect 5680 16398 5684 16409
rect 5684 16398 5700 16409
rect 5700 16398 5736 16409
rect 5762 16398 5768 16409
rect 5768 16398 5818 16409
rect 5844 16398 5900 16454
rect 5926 16398 5982 16454
rect 6008 16398 6064 16454
rect 6090 16398 6146 16454
rect 6172 16398 6228 16454
rect 6254 16398 6310 16454
rect 6336 16398 6392 16454
rect 6418 16398 6474 16454
rect 6500 16422 6552 16454
rect 6552 16422 6556 16454
rect 6582 16422 6604 16454
rect 6604 16422 6620 16454
rect 6620 16422 6638 16454
rect 6664 16422 6672 16454
rect 6672 16422 6688 16454
rect 6688 16422 6720 16454
rect 6500 16409 6556 16422
rect 6582 16409 6638 16422
rect 6664 16409 6720 16422
rect 6500 16398 6552 16409
rect 6552 16398 6556 16409
rect 6582 16398 6604 16409
rect 6604 16398 6620 16409
rect 6620 16398 6638 16409
rect 6664 16398 6672 16409
rect 6672 16398 6688 16409
rect 6688 16398 6720 16409
rect 6746 16398 6802 16454
rect 6828 16398 6884 16454
rect 6909 16398 6965 16454
rect 6990 16398 7046 16454
rect 7071 16398 7127 16454
rect 7152 16398 7208 16454
rect 7233 16398 7289 16454
rect 7314 16398 7370 16454
rect 5188 16318 5244 16374
rect 5270 16318 5326 16374
rect 5352 16318 5408 16374
rect 5434 16318 5490 16374
rect 5516 16318 5572 16374
rect 5598 16357 5632 16374
rect 5632 16357 5654 16374
rect 5680 16357 5684 16374
rect 5684 16357 5700 16374
rect 5700 16357 5736 16374
rect 5762 16357 5768 16374
rect 5768 16357 5818 16374
rect 5598 16344 5654 16357
rect 5680 16344 5736 16357
rect 5762 16344 5818 16357
rect 5598 16318 5632 16344
rect 5632 16318 5654 16344
rect 5680 16318 5684 16344
rect 5684 16318 5700 16344
rect 5700 16318 5736 16344
rect 5762 16318 5768 16344
rect 5768 16318 5818 16344
rect 5844 16318 5900 16374
rect 5926 16318 5982 16374
rect 6008 16318 6064 16374
rect 6090 16318 6146 16374
rect 6172 16318 6228 16374
rect 6254 16318 6310 16374
rect 6336 16318 6392 16374
rect 6418 16318 6474 16374
rect 6500 16357 6552 16374
rect 6552 16357 6556 16374
rect 6582 16357 6604 16374
rect 6604 16357 6620 16374
rect 6620 16357 6638 16374
rect 6664 16357 6672 16374
rect 6672 16357 6688 16374
rect 6688 16357 6720 16374
rect 6500 16344 6556 16357
rect 6582 16344 6638 16357
rect 6664 16344 6720 16357
rect 6500 16318 6552 16344
rect 6552 16318 6556 16344
rect 6582 16318 6604 16344
rect 6604 16318 6620 16344
rect 6620 16318 6638 16344
rect 6664 16318 6672 16344
rect 6672 16318 6688 16344
rect 6688 16318 6720 16344
rect 6746 16318 6802 16374
rect 6828 16318 6884 16374
rect 6909 16318 6965 16374
rect 6990 16318 7046 16374
rect 7071 16318 7127 16374
rect 7152 16318 7208 16374
rect 7233 16318 7289 16374
rect 7314 16318 7370 16374
rect 5188 16238 5244 16294
rect 5270 16238 5326 16294
rect 5352 16238 5408 16294
rect 5434 16238 5490 16294
rect 5516 16238 5572 16294
rect 5598 16292 5632 16294
rect 5632 16292 5654 16294
rect 5680 16292 5684 16294
rect 5684 16292 5700 16294
rect 5700 16292 5736 16294
rect 5762 16292 5768 16294
rect 5768 16292 5818 16294
rect 5598 16279 5654 16292
rect 5680 16279 5736 16292
rect 5762 16279 5818 16292
rect 5598 16238 5632 16279
rect 5632 16238 5654 16279
rect 5680 16238 5684 16279
rect 5684 16238 5700 16279
rect 5700 16238 5736 16279
rect 5762 16238 5768 16279
rect 5768 16238 5818 16279
rect 5844 16238 5900 16294
rect 5926 16238 5982 16294
rect 6008 16238 6064 16294
rect 6090 16238 6146 16294
rect 6172 16238 6228 16294
rect 6254 16238 6310 16294
rect 6336 16238 6392 16294
rect 6418 16238 6474 16294
rect 6500 16292 6552 16294
rect 6552 16292 6556 16294
rect 6582 16292 6604 16294
rect 6604 16292 6620 16294
rect 6620 16292 6638 16294
rect 6664 16292 6672 16294
rect 6672 16292 6688 16294
rect 6688 16292 6720 16294
rect 6500 16279 6556 16292
rect 6582 16279 6638 16292
rect 6664 16279 6720 16292
rect 6500 16238 6552 16279
rect 6552 16238 6556 16279
rect 6582 16238 6604 16279
rect 6604 16238 6620 16279
rect 6620 16238 6638 16279
rect 6664 16238 6672 16279
rect 6672 16238 6688 16279
rect 6688 16238 6720 16279
rect 6746 16238 6802 16294
rect 6828 16238 6884 16294
rect 6909 16238 6965 16294
rect 6990 16238 7046 16294
rect 7071 16238 7127 16294
rect 7152 16238 7208 16294
rect 7233 16238 7289 16294
rect 7314 16238 7370 16294
rect 5188 16158 5244 16214
rect 5270 16158 5326 16214
rect 5352 16158 5408 16214
rect 5434 16158 5490 16214
rect 5516 16158 5572 16214
rect 5598 16162 5632 16214
rect 5632 16162 5654 16214
rect 5680 16162 5684 16214
rect 5684 16162 5700 16214
rect 5700 16162 5736 16214
rect 5762 16162 5768 16214
rect 5768 16162 5818 16214
rect 5598 16158 5654 16162
rect 5680 16158 5736 16162
rect 5762 16158 5818 16162
rect 5844 16158 5900 16214
rect 5926 16158 5982 16214
rect 6008 16158 6064 16214
rect 6090 16158 6146 16214
rect 6172 16158 6228 16214
rect 6254 16158 6310 16214
rect 6336 16158 6392 16214
rect 6418 16158 6474 16214
rect 6500 16162 6552 16214
rect 6552 16162 6556 16214
rect 6582 16162 6604 16214
rect 6604 16162 6620 16214
rect 6620 16162 6638 16214
rect 6664 16162 6672 16214
rect 6672 16162 6688 16214
rect 6688 16162 6720 16214
rect 6500 16158 6556 16162
rect 6582 16158 6638 16162
rect 6664 16158 6720 16162
rect 6746 16158 6802 16214
rect 6828 16158 6884 16214
rect 6909 16158 6965 16214
rect 6990 16158 7046 16214
rect 7071 16158 7127 16214
rect 7152 16158 7208 16214
rect 7233 16158 7289 16214
rect 7314 16158 7370 16214
rect 7587 15773 7643 15829
rect 7669 15773 7725 15829
rect 7751 15773 7807 15829
rect 7833 15773 7889 15829
rect 7915 15825 7971 15829
rect 7997 15825 8053 15829
rect 8079 15825 8135 15829
rect 7915 15773 7961 15825
rect 7961 15773 7971 15825
rect 7997 15773 8013 15825
rect 8013 15773 8039 15825
rect 8039 15773 8053 15825
rect 8079 15773 8091 15825
rect 8091 15773 8135 15825
rect 8161 15773 8217 15829
rect 8243 15773 8299 15829
rect 8325 15773 8381 15829
rect 8407 15773 8463 15829
rect 8489 15773 8545 15829
rect 8571 15773 8627 15829
rect 8653 15773 8709 15829
rect 8735 15773 8791 15829
rect 8817 15773 8873 15829
rect 8899 15825 8955 15829
rect 8981 15825 9037 15829
rect 8899 15773 8933 15825
rect 8933 15773 8955 15825
rect 8981 15773 9011 15825
rect 9011 15773 9037 15825
rect 9063 15773 9119 15829
rect 9145 15773 9201 15829
rect 9227 15773 9283 15829
rect 9308 15773 9364 15829
rect 9389 15773 9445 15829
rect 9470 15773 9526 15829
rect 9551 15773 9607 15829
rect 9632 15773 9688 15829
rect 9713 15773 9769 15829
rect 7587 15693 7643 15749
rect 7669 15693 7725 15749
rect 7751 15693 7807 15749
rect 7833 15693 7889 15749
rect 7915 15709 7961 15749
rect 7961 15709 7971 15749
rect 7997 15709 8013 15749
rect 8013 15709 8039 15749
rect 8039 15709 8053 15749
rect 8079 15709 8091 15749
rect 8091 15709 8135 15749
rect 7915 15697 7971 15709
rect 7997 15697 8053 15709
rect 8079 15697 8135 15709
rect 7915 15693 7961 15697
rect 7961 15693 7971 15697
rect 7997 15693 8013 15697
rect 8013 15693 8039 15697
rect 8039 15693 8053 15697
rect 8079 15693 8091 15697
rect 8091 15693 8135 15697
rect 8161 15693 8217 15749
rect 8243 15693 8299 15749
rect 8325 15693 8381 15749
rect 8407 15693 8463 15749
rect 8489 15693 8545 15749
rect 8571 15693 8627 15749
rect 8653 15693 8709 15749
rect 8735 15693 8791 15749
rect 8817 15693 8873 15749
rect 8899 15709 8933 15749
rect 8933 15709 8955 15749
rect 8981 15709 9011 15749
rect 9011 15709 9037 15749
rect 8899 15697 8955 15709
rect 8981 15697 9037 15709
rect 8899 15693 8933 15697
rect 8933 15693 8955 15697
rect 8981 15693 9011 15697
rect 9011 15693 9037 15697
rect 9063 15693 9119 15749
rect 9145 15693 9201 15749
rect 9227 15693 9283 15749
rect 9308 15693 9364 15749
rect 9389 15693 9445 15749
rect 9470 15693 9526 15749
rect 9551 15693 9607 15749
rect 9632 15693 9688 15749
rect 9713 15693 9769 15749
rect 7587 15613 7643 15669
rect 7669 15613 7725 15669
rect 7751 15613 7807 15669
rect 7833 15613 7889 15669
rect 7915 15645 7961 15669
rect 7961 15645 7971 15669
rect 7997 15645 8013 15669
rect 8013 15645 8039 15669
rect 8039 15645 8053 15669
rect 8079 15645 8091 15669
rect 8091 15645 8135 15669
rect 7915 15633 7971 15645
rect 7997 15633 8053 15645
rect 8079 15633 8135 15645
rect 7915 15613 7961 15633
rect 7961 15613 7971 15633
rect 7997 15613 8013 15633
rect 8013 15613 8039 15633
rect 8039 15613 8053 15633
rect 8079 15613 8091 15633
rect 8091 15613 8135 15633
rect 8161 15613 8217 15669
rect 8243 15613 8299 15669
rect 8325 15613 8381 15669
rect 8407 15613 8463 15669
rect 8489 15613 8545 15669
rect 8571 15613 8627 15669
rect 8653 15613 8709 15669
rect 8735 15613 8791 15669
rect 8817 15613 8873 15669
rect 8899 15645 8933 15669
rect 8933 15645 8955 15669
rect 8981 15645 9011 15669
rect 9011 15645 9037 15669
rect 8899 15633 8955 15645
rect 8981 15633 9037 15645
rect 8899 15613 8933 15633
rect 8933 15613 8955 15633
rect 8981 15613 9011 15633
rect 9011 15613 9037 15633
rect 9063 15613 9119 15669
rect 9145 15613 9201 15669
rect 9227 15613 9283 15669
rect 9308 15613 9364 15669
rect 9389 15613 9445 15669
rect 9470 15613 9526 15669
rect 9551 15613 9607 15669
rect 9632 15613 9688 15669
rect 9713 15613 9769 15669
rect 7587 15533 7643 15589
rect 7669 15533 7725 15589
rect 7751 15533 7807 15589
rect 7833 15533 7889 15589
rect 7915 15581 7961 15589
rect 7961 15581 7971 15589
rect 7997 15581 8013 15589
rect 8013 15581 8039 15589
rect 8039 15581 8053 15589
rect 8079 15581 8091 15589
rect 8091 15581 8135 15589
rect 7915 15569 7971 15581
rect 7997 15569 8053 15581
rect 8079 15569 8135 15581
rect 7915 15533 7961 15569
rect 7961 15533 7971 15569
rect 7997 15533 8013 15569
rect 8013 15533 8039 15569
rect 8039 15533 8053 15569
rect 8079 15533 8091 15569
rect 8091 15533 8135 15569
rect 8161 15533 8217 15589
rect 8243 15533 8299 15589
rect 8325 15533 8381 15589
rect 8407 15533 8463 15589
rect 8489 15533 8545 15589
rect 8571 15533 8627 15589
rect 8653 15533 8709 15589
rect 8735 15533 8791 15589
rect 8817 15533 8873 15589
rect 8899 15581 8933 15589
rect 8933 15581 8955 15589
rect 8981 15581 9011 15589
rect 9011 15581 9037 15589
rect 8899 15569 8955 15581
rect 8981 15569 9037 15581
rect 8899 15533 8933 15569
rect 8933 15533 8955 15569
rect 8981 15533 9011 15569
rect 9011 15533 9037 15569
rect 9063 15533 9119 15589
rect 9145 15533 9201 15589
rect 9227 15533 9283 15589
rect 9308 15533 9364 15589
rect 9389 15533 9445 15589
rect 9470 15533 9526 15589
rect 9551 15533 9607 15589
rect 9632 15533 9688 15589
rect 9713 15533 9769 15589
rect 7587 15453 7643 15509
rect 7669 15453 7725 15509
rect 7751 15453 7807 15509
rect 7833 15453 7889 15509
rect 7915 15505 7971 15509
rect 7997 15505 8053 15509
rect 8079 15505 8135 15509
rect 7915 15453 7961 15505
rect 7961 15453 7971 15505
rect 7997 15453 8013 15505
rect 8013 15453 8039 15505
rect 8039 15453 8053 15505
rect 8079 15453 8091 15505
rect 8091 15453 8135 15505
rect 8161 15453 8217 15509
rect 8243 15453 8299 15509
rect 8325 15453 8381 15509
rect 8407 15453 8463 15509
rect 8489 15453 8545 15509
rect 8571 15453 8627 15509
rect 8653 15453 8709 15509
rect 8735 15453 8791 15509
rect 8817 15453 8873 15509
rect 8899 15505 8955 15509
rect 8981 15505 9037 15509
rect 8899 15453 8933 15505
rect 8933 15453 8955 15505
rect 8981 15453 9011 15505
rect 9011 15453 9037 15505
rect 9063 15453 9119 15509
rect 9145 15453 9201 15509
rect 9227 15453 9283 15509
rect 9308 15453 9364 15509
rect 9389 15453 9445 15509
rect 9470 15453 9526 15509
rect 9551 15453 9607 15509
rect 9632 15453 9688 15509
rect 9713 15453 9769 15509
rect 7587 15373 7643 15429
rect 7669 15373 7725 15429
rect 7751 15373 7807 15429
rect 7833 15373 7889 15429
rect 7915 15389 7961 15429
rect 7961 15389 7971 15429
rect 7997 15389 8013 15429
rect 8013 15389 8039 15429
rect 8039 15389 8053 15429
rect 8079 15389 8091 15429
rect 8091 15389 8135 15429
rect 7915 15377 7971 15389
rect 7997 15377 8053 15389
rect 8079 15377 8135 15389
rect 7915 15373 7961 15377
rect 7961 15373 7971 15377
rect 7997 15373 8013 15377
rect 8013 15373 8039 15377
rect 8039 15373 8053 15377
rect 8079 15373 8091 15377
rect 8091 15373 8135 15377
rect 8161 15373 8217 15429
rect 8243 15373 8299 15429
rect 8325 15373 8381 15429
rect 8407 15373 8463 15429
rect 8489 15373 8545 15429
rect 8571 15373 8627 15429
rect 8653 15373 8709 15429
rect 8735 15373 8791 15429
rect 8817 15373 8873 15429
rect 8899 15389 8933 15429
rect 8933 15389 8955 15429
rect 8981 15389 9011 15429
rect 9011 15389 9037 15429
rect 8899 15377 8955 15389
rect 8981 15377 9037 15389
rect 8899 15373 8933 15377
rect 8933 15373 8955 15377
rect 8981 15373 9011 15377
rect 9011 15373 9037 15377
rect 9063 15373 9119 15429
rect 9145 15373 9201 15429
rect 9227 15373 9283 15429
rect 9308 15373 9364 15429
rect 9389 15373 9445 15429
rect 9470 15373 9526 15429
rect 9551 15373 9607 15429
rect 9632 15373 9688 15429
rect 9713 15373 9769 15429
rect 7587 15293 7643 15349
rect 7669 15293 7725 15349
rect 7751 15293 7807 15349
rect 7833 15293 7889 15349
rect 7915 15325 7961 15349
rect 7961 15325 7971 15349
rect 7997 15325 8013 15349
rect 8013 15325 8039 15349
rect 8039 15325 8053 15349
rect 8079 15325 8091 15349
rect 8091 15325 8135 15349
rect 7915 15313 7971 15325
rect 7997 15313 8053 15325
rect 8079 15313 8135 15325
rect 7915 15293 7961 15313
rect 7961 15293 7971 15313
rect 7997 15293 8013 15313
rect 8013 15293 8039 15313
rect 8039 15293 8053 15313
rect 8079 15293 8091 15313
rect 8091 15293 8135 15313
rect 8161 15293 8217 15349
rect 8243 15293 8299 15349
rect 8325 15293 8381 15349
rect 8407 15293 8463 15349
rect 8489 15293 8545 15349
rect 8571 15293 8627 15349
rect 8653 15293 8709 15349
rect 8735 15293 8791 15349
rect 8817 15293 8873 15349
rect 8899 15325 8933 15349
rect 8933 15325 8955 15349
rect 8981 15325 9011 15349
rect 9011 15325 9037 15349
rect 8899 15313 8955 15325
rect 8981 15313 9037 15325
rect 8899 15293 8933 15313
rect 8933 15293 8955 15313
rect 8981 15293 9011 15313
rect 9011 15293 9037 15313
rect 9063 15293 9119 15349
rect 9145 15293 9201 15349
rect 9227 15293 9283 15349
rect 9308 15293 9364 15349
rect 9389 15293 9445 15349
rect 9470 15293 9526 15349
rect 9551 15293 9607 15349
rect 9632 15293 9688 15349
rect 9713 15293 9769 15349
rect 7587 15213 7643 15269
rect 7669 15213 7725 15269
rect 7751 15213 7807 15269
rect 7833 15213 7889 15269
rect 7915 15261 7961 15269
rect 7961 15261 7971 15269
rect 7997 15261 8013 15269
rect 8013 15261 8039 15269
rect 8039 15261 8053 15269
rect 8079 15261 8091 15269
rect 8091 15261 8135 15269
rect 7915 15249 7971 15261
rect 7997 15249 8053 15261
rect 8079 15249 8135 15261
rect 7915 15213 7961 15249
rect 7961 15213 7971 15249
rect 7997 15213 8013 15249
rect 8013 15213 8039 15249
rect 8039 15213 8053 15249
rect 8079 15213 8091 15249
rect 8091 15213 8135 15249
rect 8161 15213 8217 15269
rect 8243 15213 8299 15269
rect 8325 15213 8381 15269
rect 8407 15213 8463 15269
rect 8489 15213 8545 15269
rect 8571 15213 8627 15269
rect 8653 15213 8709 15269
rect 8735 15213 8791 15269
rect 8817 15213 8873 15269
rect 8899 15261 8933 15269
rect 8933 15261 8955 15269
rect 8981 15261 9011 15269
rect 9011 15261 9037 15269
rect 8899 15249 8955 15261
rect 8981 15249 9037 15261
rect 8899 15213 8933 15249
rect 8933 15213 8955 15249
rect 8981 15213 9011 15249
rect 9011 15213 9037 15249
rect 9063 15213 9119 15269
rect 9145 15213 9201 15269
rect 9227 15213 9283 15269
rect 9308 15213 9364 15269
rect 9389 15213 9445 15269
rect 9470 15213 9526 15269
rect 9551 15213 9607 15269
rect 9632 15213 9688 15269
rect 9713 15213 9769 15269
rect 7587 15133 7643 15189
rect 7669 15133 7725 15189
rect 7751 15133 7807 15189
rect 7833 15133 7889 15189
rect 7915 15185 7971 15189
rect 7997 15185 8053 15189
rect 8079 15185 8135 15189
rect 7915 15133 7961 15185
rect 7961 15133 7971 15185
rect 7997 15133 8013 15185
rect 8013 15133 8039 15185
rect 8039 15133 8053 15185
rect 8079 15133 8091 15185
rect 8091 15133 8135 15185
rect 8161 15133 8217 15189
rect 8243 15133 8299 15189
rect 8325 15133 8381 15189
rect 8407 15133 8463 15189
rect 8489 15133 8545 15189
rect 8571 15133 8627 15189
rect 8653 15133 8709 15189
rect 8735 15133 8791 15189
rect 8817 15133 8873 15189
rect 8899 15185 8955 15189
rect 8981 15185 9037 15189
rect 8899 15133 8933 15185
rect 8933 15133 8955 15185
rect 8981 15133 9011 15185
rect 9011 15133 9037 15185
rect 9063 15133 9119 15189
rect 9145 15133 9201 15189
rect 9227 15133 9283 15189
rect 9308 15133 9364 15189
rect 9389 15133 9445 15189
rect 9470 15133 9526 15189
rect 9551 15133 9607 15189
rect 9632 15133 9688 15189
rect 9713 15133 9769 15189
rect 7587 15053 7643 15109
rect 7669 15053 7725 15109
rect 7751 15053 7807 15109
rect 7833 15053 7889 15109
rect 7915 15069 7961 15109
rect 7961 15069 7971 15109
rect 7997 15069 8013 15109
rect 8013 15069 8039 15109
rect 8039 15069 8053 15109
rect 8079 15069 8091 15109
rect 8091 15069 8135 15109
rect 7915 15057 7971 15069
rect 7997 15057 8053 15069
rect 8079 15057 8135 15069
rect 7915 15053 7961 15057
rect 7961 15053 7971 15057
rect 7997 15053 8013 15057
rect 8013 15053 8039 15057
rect 8039 15053 8053 15057
rect 8079 15053 8091 15057
rect 8091 15053 8135 15057
rect 8161 15053 8217 15109
rect 8243 15053 8299 15109
rect 8325 15053 8381 15109
rect 8407 15053 8463 15109
rect 8489 15053 8545 15109
rect 8571 15053 8627 15109
rect 8653 15053 8709 15109
rect 8735 15053 8791 15109
rect 8817 15053 8873 15109
rect 8899 15069 8933 15109
rect 8933 15069 8955 15109
rect 8981 15069 9011 15109
rect 9011 15069 9037 15109
rect 8899 15057 8955 15069
rect 8981 15057 9037 15069
rect 8899 15053 8933 15057
rect 8933 15053 8955 15057
rect 8981 15053 9011 15057
rect 9011 15053 9037 15057
rect 9063 15053 9119 15109
rect 9145 15053 9201 15109
rect 9227 15053 9283 15109
rect 9308 15053 9364 15109
rect 9389 15053 9445 15109
rect 9470 15053 9526 15109
rect 9551 15053 9607 15109
rect 9632 15053 9688 15109
rect 9713 15053 9769 15109
rect 7587 14973 7643 15029
rect 7669 14973 7725 15029
rect 7751 14973 7807 15029
rect 7833 14973 7889 15029
rect 7915 15005 7961 15029
rect 7961 15005 7971 15029
rect 7997 15005 8013 15029
rect 8013 15005 8039 15029
rect 8039 15005 8053 15029
rect 8079 15005 8091 15029
rect 8091 15005 8135 15029
rect 7915 14993 7971 15005
rect 7997 14993 8053 15005
rect 8079 14993 8135 15005
rect 7915 14973 7961 14993
rect 7961 14973 7971 14993
rect 7997 14973 8013 14993
rect 8013 14973 8039 14993
rect 8039 14973 8053 14993
rect 8079 14973 8091 14993
rect 8091 14973 8135 14993
rect 8161 14973 8217 15029
rect 8243 14973 8299 15029
rect 8325 14973 8381 15029
rect 8407 14973 8463 15029
rect 8489 14973 8545 15029
rect 8571 14973 8627 15029
rect 8653 14973 8709 15029
rect 8735 14973 8791 15029
rect 8817 14973 8873 15029
rect 8899 15005 8933 15029
rect 8933 15005 8955 15029
rect 8981 15005 9011 15029
rect 9011 15005 9037 15029
rect 8899 14993 8955 15005
rect 8981 14993 9037 15005
rect 8899 14973 8933 14993
rect 8933 14973 8955 14993
rect 8981 14973 9011 14993
rect 9011 14973 9037 14993
rect 9063 14973 9119 15029
rect 9145 14973 9201 15029
rect 9227 14973 9283 15029
rect 9308 14973 9364 15029
rect 9389 14973 9445 15029
rect 9470 14973 9526 15029
rect 9551 14973 9607 15029
rect 9632 14973 9688 15029
rect 9713 14973 9769 15029
rect 7587 14893 7643 14949
rect 7669 14893 7725 14949
rect 7751 14893 7807 14949
rect 7833 14893 7889 14949
rect 7915 14941 7961 14949
rect 7961 14941 7971 14949
rect 7997 14941 8013 14949
rect 8013 14941 8039 14949
rect 8039 14941 8053 14949
rect 8079 14941 8091 14949
rect 8091 14941 8135 14949
rect 7915 14929 7971 14941
rect 7997 14929 8053 14941
rect 8079 14929 8135 14941
rect 7915 14893 7961 14929
rect 7961 14893 7971 14929
rect 7997 14893 8013 14929
rect 8013 14893 8039 14929
rect 8039 14893 8053 14929
rect 8079 14893 8091 14929
rect 8091 14893 8135 14929
rect 8161 14893 8217 14949
rect 8243 14893 8299 14949
rect 8325 14893 8381 14949
rect 8407 14893 8463 14949
rect 8489 14893 8545 14949
rect 8571 14893 8627 14949
rect 8653 14893 8709 14949
rect 8735 14893 8791 14949
rect 8817 14893 8873 14949
rect 8899 14941 8933 14949
rect 8933 14941 8955 14949
rect 8981 14941 9011 14949
rect 9011 14941 9037 14949
rect 8899 14929 8955 14941
rect 8981 14929 9037 14941
rect 8899 14893 8933 14929
rect 8933 14893 8955 14929
rect 8981 14893 9011 14929
rect 9011 14893 9037 14929
rect 9063 14893 9119 14949
rect 9145 14893 9201 14949
rect 9227 14893 9283 14949
rect 9308 14893 9364 14949
rect 9389 14893 9445 14949
rect 9470 14893 9526 14949
rect 9551 14893 9607 14949
rect 9632 14893 9688 14949
rect 9713 14893 9769 14949
rect 7587 14813 7643 14869
rect 7669 14813 7725 14869
rect 7751 14813 7807 14869
rect 7833 14813 7889 14869
rect 7915 14864 7971 14869
rect 7997 14864 8053 14869
rect 8079 14864 8135 14869
rect 7915 14813 7961 14864
rect 7961 14813 7971 14864
rect 7997 14813 8013 14864
rect 8013 14813 8039 14864
rect 8039 14813 8053 14864
rect 8079 14813 8091 14864
rect 8091 14813 8135 14864
rect 8161 14813 8217 14869
rect 8243 14813 8299 14869
rect 8325 14813 8381 14869
rect 8407 14813 8463 14869
rect 8489 14813 8545 14869
rect 8571 14813 8627 14869
rect 8653 14813 8709 14869
rect 8735 14813 8791 14869
rect 8817 14813 8873 14869
rect 8899 14864 8955 14869
rect 8981 14864 9037 14869
rect 8899 14813 8933 14864
rect 8933 14813 8955 14864
rect 8981 14813 9011 14864
rect 9011 14813 9037 14864
rect 9063 14813 9119 14869
rect 9145 14813 9201 14869
rect 9227 14813 9283 14869
rect 9308 14813 9364 14869
rect 9389 14813 9445 14869
rect 9470 14813 9526 14869
rect 9551 14813 9607 14869
rect 9632 14813 9688 14869
rect 9713 14813 9769 14869
rect 7587 14733 7643 14789
rect 7669 14733 7725 14789
rect 7751 14733 7807 14789
rect 7833 14733 7889 14789
rect 7915 14747 7961 14789
rect 7961 14747 7971 14789
rect 7997 14747 8013 14789
rect 8013 14747 8039 14789
rect 8039 14747 8053 14789
rect 8079 14747 8091 14789
rect 8091 14747 8135 14789
rect 7915 14734 7971 14747
rect 7997 14734 8053 14747
rect 8079 14734 8135 14747
rect 7915 14733 7961 14734
rect 7961 14733 7971 14734
rect 7997 14733 8013 14734
rect 8013 14733 8039 14734
rect 8039 14733 8053 14734
rect 8079 14733 8091 14734
rect 8091 14733 8135 14734
rect 8161 14733 8217 14789
rect 8243 14733 8299 14789
rect 8325 14733 8381 14789
rect 8407 14733 8463 14789
rect 8489 14733 8545 14789
rect 8571 14733 8627 14789
rect 8653 14733 8709 14789
rect 8735 14733 8791 14789
rect 8817 14733 8873 14789
rect 8899 14747 8933 14789
rect 8933 14747 8955 14789
rect 8981 14747 9011 14789
rect 9011 14747 9037 14789
rect 8899 14734 8955 14747
rect 8981 14734 9037 14747
rect 8899 14733 8933 14734
rect 8933 14733 8955 14734
rect 8981 14733 9011 14734
rect 9011 14733 9037 14734
rect 9063 14733 9119 14789
rect 9145 14733 9201 14789
rect 9227 14733 9283 14789
rect 9308 14733 9364 14789
rect 9389 14733 9445 14789
rect 9470 14733 9526 14789
rect 9551 14733 9607 14789
rect 9632 14733 9688 14789
rect 9713 14733 9769 14789
rect 7587 14653 7643 14709
rect 7669 14653 7725 14709
rect 7751 14653 7807 14709
rect 7833 14653 7889 14709
rect 7915 14682 7961 14709
rect 7961 14682 7971 14709
rect 7997 14682 8013 14709
rect 8013 14682 8039 14709
rect 8039 14682 8053 14709
rect 8079 14682 8091 14709
rect 8091 14682 8135 14709
rect 7915 14669 7971 14682
rect 7997 14669 8053 14682
rect 8079 14669 8135 14682
rect 7915 14653 7961 14669
rect 7961 14653 7971 14669
rect 7997 14653 8013 14669
rect 8013 14653 8039 14669
rect 8039 14653 8053 14669
rect 8079 14653 8091 14669
rect 8091 14653 8135 14669
rect 8161 14653 8217 14709
rect 8243 14653 8299 14709
rect 8325 14653 8381 14709
rect 8407 14653 8463 14709
rect 8489 14653 8545 14709
rect 8571 14653 8627 14709
rect 8653 14653 8709 14709
rect 8735 14653 8791 14709
rect 8817 14653 8873 14709
rect 8899 14682 8933 14709
rect 8933 14682 8955 14709
rect 8981 14682 9011 14709
rect 9011 14682 9037 14709
rect 8899 14669 8955 14682
rect 8981 14669 9037 14682
rect 8899 14653 8933 14669
rect 8933 14653 8955 14669
rect 8981 14653 9011 14669
rect 9011 14653 9037 14669
rect 9063 14653 9119 14709
rect 9145 14653 9201 14709
rect 9227 14653 9283 14709
rect 9308 14653 9364 14709
rect 9389 14653 9445 14709
rect 9470 14653 9526 14709
rect 9551 14653 9607 14709
rect 9632 14653 9688 14709
rect 9713 14653 9769 14709
rect 7587 14573 7643 14629
rect 7669 14573 7725 14629
rect 7751 14573 7807 14629
rect 7833 14573 7889 14629
rect 7915 14617 7961 14629
rect 7961 14617 7971 14629
rect 7997 14617 8013 14629
rect 8013 14617 8039 14629
rect 8039 14617 8053 14629
rect 8079 14617 8091 14629
rect 8091 14617 8135 14629
rect 7915 14604 7971 14617
rect 7997 14604 8053 14617
rect 8079 14604 8135 14617
rect 7915 14573 7961 14604
rect 7961 14573 7971 14604
rect 7997 14573 8013 14604
rect 8013 14573 8039 14604
rect 8039 14573 8053 14604
rect 8079 14573 8091 14604
rect 8091 14573 8135 14604
rect 8161 14573 8217 14629
rect 8243 14573 8299 14629
rect 8325 14573 8381 14629
rect 8407 14573 8463 14629
rect 8489 14573 8545 14629
rect 8571 14573 8627 14629
rect 8653 14573 8709 14629
rect 8735 14573 8791 14629
rect 8817 14573 8873 14629
rect 8899 14617 8933 14629
rect 8933 14617 8955 14629
rect 8981 14617 9011 14629
rect 9011 14617 9037 14629
rect 8899 14604 8955 14617
rect 8981 14604 9037 14617
rect 8899 14573 8933 14604
rect 8933 14573 8955 14604
rect 8981 14573 9011 14604
rect 9011 14573 9037 14604
rect 9063 14573 9119 14629
rect 9145 14573 9201 14629
rect 9227 14573 9283 14629
rect 9308 14573 9364 14629
rect 9389 14573 9445 14629
rect 9470 14573 9526 14629
rect 9551 14573 9607 14629
rect 9632 14573 9688 14629
rect 9713 14573 9769 14629
rect 7587 14493 7643 14549
rect 7669 14493 7725 14549
rect 7751 14493 7807 14549
rect 7833 14493 7889 14549
rect 7915 14539 7971 14549
rect 7997 14539 8053 14549
rect 8079 14539 8135 14549
rect 7915 14493 7961 14539
rect 7961 14493 7971 14539
rect 7997 14493 8013 14539
rect 8013 14493 8039 14539
rect 8039 14493 8053 14539
rect 8079 14493 8091 14539
rect 8091 14493 8135 14539
rect 8161 14493 8217 14549
rect 8243 14493 8299 14549
rect 8325 14493 8381 14549
rect 8407 14493 8463 14549
rect 8489 14493 8545 14549
rect 8571 14493 8627 14549
rect 8653 14493 8709 14549
rect 8735 14493 8791 14549
rect 8817 14493 8873 14549
rect 8899 14539 8955 14549
rect 8981 14539 9037 14549
rect 8899 14493 8933 14539
rect 8933 14493 8955 14539
rect 8981 14493 9011 14539
rect 9011 14493 9037 14539
rect 9063 14493 9119 14549
rect 9145 14493 9201 14549
rect 9227 14493 9283 14549
rect 9308 14493 9364 14549
rect 9389 14493 9445 14549
rect 9470 14493 9526 14549
rect 9551 14493 9607 14549
rect 9632 14493 9688 14549
rect 9713 14493 9769 14549
rect 7587 14413 7643 14469
rect 7669 14413 7725 14469
rect 7751 14413 7807 14469
rect 7833 14413 7889 14469
rect 7915 14422 7961 14469
rect 7961 14422 7971 14469
rect 7997 14422 8013 14469
rect 8013 14422 8039 14469
rect 8039 14422 8053 14469
rect 8079 14422 8091 14469
rect 8091 14422 8135 14469
rect 7915 14413 7971 14422
rect 7997 14413 8053 14422
rect 8079 14413 8135 14422
rect 8161 14413 8217 14469
rect 8243 14413 8299 14469
rect 8325 14413 8381 14469
rect 8407 14413 8463 14469
rect 8489 14413 8545 14469
rect 8571 14413 8627 14469
rect 8653 14413 8709 14469
rect 8735 14413 8791 14469
rect 8817 14413 8873 14469
rect 8899 14422 8933 14469
rect 8933 14422 8955 14469
rect 8981 14422 9011 14469
rect 9011 14422 9037 14469
rect 8899 14413 8955 14422
rect 8981 14413 9037 14422
rect 9063 14413 9119 14469
rect 9145 14413 9201 14469
rect 9227 14413 9283 14469
rect 9308 14413 9364 14469
rect 9389 14413 9445 14469
rect 9470 14413 9526 14469
rect 9551 14413 9607 14469
rect 9632 14413 9688 14469
rect 9713 14413 9769 14469
rect 7587 14333 7643 14389
rect 7669 14333 7725 14389
rect 7751 14333 7807 14389
rect 7833 14333 7889 14389
rect 7915 14357 7961 14389
rect 7961 14357 7971 14389
rect 7997 14357 8013 14389
rect 8013 14357 8039 14389
rect 8039 14357 8053 14389
rect 8079 14357 8091 14389
rect 8091 14357 8135 14389
rect 7915 14344 7971 14357
rect 7997 14344 8053 14357
rect 8079 14344 8135 14357
rect 7915 14333 7961 14344
rect 7961 14333 7971 14344
rect 7997 14333 8013 14344
rect 8013 14333 8039 14344
rect 8039 14333 8053 14344
rect 8079 14333 8091 14344
rect 8091 14333 8135 14344
rect 8161 14333 8217 14389
rect 8243 14333 8299 14389
rect 8325 14333 8381 14389
rect 8407 14333 8463 14389
rect 8489 14333 8545 14389
rect 8571 14333 8627 14389
rect 8653 14333 8709 14389
rect 8735 14333 8791 14389
rect 8817 14333 8873 14389
rect 8899 14357 8933 14389
rect 8933 14357 8955 14389
rect 8981 14357 9011 14389
rect 9011 14357 9037 14389
rect 8899 14344 8955 14357
rect 8981 14344 9037 14357
rect 8899 14333 8933 14344
rect 8933 14333 8955 14344
rect 8981 14333 9011 14344
rect 9011 14333 9037 14344
rect 9063 14333 9119 14389
rect 9145 14333 9201 14389
rect 9227 14333 9283 14389
rect 9308 14333 9364 14389
rect 9389 14333 9445 14389
rect 9470 14333 9526 14389
rect 9551 14333 9607 14389
rect 9632 14333 9688 14389
rect 9713 14333 9769 14389
rect 7587 14253 7643 14309
rect 7669 14253 7725 14309
rect 7751 14253 7807 14309
rect 7833 14253 7889 14309
rect 7915 14292 7961 14309
rect 7961 14292 7971 14309
rect 7997 14292 8013 14309
rect 8013 14292 8039 14309
rect 8039 14292 8053 14309
rect 8079 14292 8091 14309
rect 8091 14292 8135 14309
rect 7915 14279 7971 14292
rect 7997 14279 8053 14292
rect 8079 14279 8135 14292
rect 7915 14253 7961 14279
rect 7961 14253 7971 14279
rect 7997 14253 8013 14279
rect 8013 14253 8039 14279
rect 8039 14253 8053 14279
rect 8079 14253 8091 14279
rect 8091 14253 8135 14279
rect 8161 14253 8217 14309
rect 8243 14253 8299 14309
rect 8325 14253 8381 14309
rect 8407 14253 8463 14309
rect 8489 14253 8545 14309
rect 8571 14253 8627 14309
rect 8653 14253 8709 14309
rect 8735 14253 8791 14309
rect 8817 14253 8873 14309
rect 8899 14292 8933 14309
rect 8933 14292 8955 14309
rect 8981 14292 9011 14309
rect 9011 14292 9037 14309
rect 8899 14279 8955 14292
rect 8981 14279 9037 14292
rect 8899 14253 8933 14279
rect 8933 14253 8955 14279
rect 8981 14253 9011 14279
rect 9011 14253 9037 14279
rect 9063 14253 9119 14309
rect 9145 14253 9201 14309
rect 9227 14253 9283 14309
rect 9308 14253 9364 14309
rect 9389 14253 9445 14309
rect 9470 14253 9526 14309
rect 9551 14253 9607 14309
rect 9632 14253 9688 14309
rect 9713 14253 9769 14309
rect 7587 14173 7643 14229
rect 7669 14173 7725 14229
rect 7751 14173 7807 14229
rect 7833 14173 7889 14229
rect 7915 14227 7961 14229
rect 7961 14227 7971 14229
rect 7997 14227 8013 14229
rect 8013 14227 8039 14229
rect 8039 14227 8053 14229
rect 8079 14227 8091 14229
rect 8091 14227 8135 14229
rect 7915 14214 7971 14227
rect 7997 14214 8053 14227
rect 8079 14214 8135 14227
rect 7915 14173 7961 14214
rect 7961 14173 7971 14214
rect 7997 14173 8013 14214
rect 8013 14173 8039 14214
rect 8039 14173 8053 14214
rect 8079 14173 8091 14214
rect 8091 14173 8135 14214
rect 8161 14173 8217 14229
rect 8243 14173 8299 14229
rect 8325 14173 8381 14229
rect 8407 14173 8463 14229
rect 8489 14173 8545 14229
rect 8571 14173 8627 14229
rect 8653 14173 8709 14229
rect 8735 14173 8791 14229
rect 8817 14173 8873 14229
rect 8899 14227 8933 14229
rect 8933 14227 8955 14229
rect 8981 14227 9011 14229
rect 9011 14227 9037 14229
rect 8899 14214 8955 14227
rect 8981 14214 9037 14227
rect 8899 14173 8933 14214
rect 8933 14173 8955 14214
rect 8981 14173 9011 14214
rect 9011 14173 9037 14214
rect 9063 14173 9119 14229
rect 9145 14173 9201 14229
rect 9227 14173 9283 14229
rect 9308 14173 9364 14229
rect 9389 14173 9445 14229
rect 9470 14173 9526 14229
rect 9551 14173 9607 14229
rect 9632 14173 9688 14229
rect 9713 14173 9769 14229
rect 7587 14093 7643 14149
rect 7669 14093 7725 14149
rect 7751 14093 7807 14149
rect 7833 14093 7889 14149
rect 7915 14097 7961 14149
rect 7961 14097 7971 14149
rect 7997 14097 8013 14149
rect 8013 14097 8039 14149
rect 8039 14097 8053 14149
rect 8079 14097 8091 14149
rect 8091 14097 8135 14149
rect 7915 14093 7971 14097
rect 7997 14093 8053 14097
rect 8079 14093 8135 14097
rect 8161 14093 8217 14149
rect 8243 14093 8299 14149
rect 8325 14093 8381 14149
rect 8407 14093 8463 14149
rect 8489 14093 8545 14149
rect 8571 14093 8627 14149
rect 8653 14093 8709 14149
rect 8735 14093 8791 14149
rect 8817 14093 8873 14149
rect 8899 14097 8933 14149
rect 8933 14097 8955 14149
rect 8981 14097 9011 14149
rect 9011 14097 9037 14149
rect 8899 14093 8955 14097
rect 8981 14093 9037 14097
rect 9063 14093 9119 14149
rect 9145 14093 9201 14149
rect 9227 14093 9283 14149
rect 9308 14093 9364 14149
rect 9389 14093 9445 14149
rect 9470 14093 9526 14149
rect 9551 14093 9607 14149
rect 9632 14093 9688 14149
rect 9713 14093 9769 14149
rect 5188 13238 5244 13294
rect 5270 13238 5326 13294
rect 5352 13238 5408 13294
rect 5434 13238 5490 13294
rect 5516 13238 5572 13294
rect 5598 13290 5654 13294
rect 5680 13290 5736 13294
rect 5762 13290 5818 13294
rect 5598 13238 5632 13290
rect 5632 13238 5654 13290
rect 5680 13238 5684 13290
rect 5684 13238 5700 13290
rect 5700 13238 5736 13290
rect 5762 13238 5768 13290
rect 5768 13238 5818 13290
rect 5844 13238 5900 13294
rect 5926 13238 5982 13294
rect 6008 13238 6064 13294
rect 6090 13238 6146 13294
rect 6172 13238 6228 13294
rect 6254 13238 6310 13294
rect 6336 13238 6392 13294
rect 6418 13238 6474 13294
rect 6500 13290 6556 13294
rect 6582 13290 6638 13294
rect 6664 13290 6720 13294
rect 6500 13238 6552 13290
rect 6552 13238 6556 13290
rect 6582 13238 6604 13290
rect 6604 13238 6620 13290
rect 6620 13238 6638 13290
rect 6664 13238 6672 13290
rect 6672 13238 6688 13290
rect 6688 13238 6720 13290
rect 6746 13238 6802 13294
rect 6828 13238 6884 13294
rect 6909 13238 6965 13294
rect 6990 13238 7046 13294
rect 7071 13238 7127 13294
rect 7152 13238 7208 13294
rect 7233 13238 7289 13294
rect 7314 13238 7370 13294
rect 5188 13158 5244 13214
rect 5270 13158 5326 13214
rect 5352 13158 5408 13214
rect 5434 13158 5490 13214
rect 5516 13158 5572 13214
rect 5598 13174 5632 13214
rect 5632 13174 5654 13214
rect 5680 13174 5684 13214
rect 5684 13174 5700 13214
rect 5700 13174 5736 13214
rect 5762 13174 5768 13214
rect 5768 13174 5818 13214
rect 5598 13162 5654 13174
rect 5680 13162 5736 13174
rect 5762 13162 5818 13174
rect 5598 13158 5632 13162
rect 5632 13158 5654 13162
rect 5680 13158 5684 13162
rect 5684 13158 5700 13162
rect 5700 13158 5736 13162
rect 5762 13158 5768 13162
rect 5768 13158 5818 13162
rect 5844 13158 5900 13214
rect 5926 13158 5982 13214
rect 6008 13158 6064 13214
rect 6090 13158 6146 13214
rect 6172 13158 6228 13214
rect 6254 13158 6310 13214
rect 6336 13158 6392 13214
rect 6418 13158 6474 13214
rect 6500 13174 6552 13214
rect 6552 13174 6556 13214
rect 6582 13174 6604 13214
rect 6604 13174 6620 13214
rect 6620 13174 6638 13214
rect 6664 13174 6672 13214
rect 6672 13174 6688 13214
rect 6688 13174 6720 13214
rect 6500 13162 6556 13174
rect 6582 13162 6638 13174
rect 6664 13162 6720 13174
rect 6500 13158 6552 13162
rect 6552 13158 6556 13162
rect 6582 13158 6604 13162
rect 6604 13158 6620 13162
rect 6620 13158 6638 13162
rect 6664 13158 6672 13162
rect 6672 13158 6688 13162
rect 6688 13158 6720 13162
rect 6746 13158 6802 13214
rect 6828 13158 6884 13214
rect 6909 13158 6965 13214
rect 6990 13158 7046 13214
rect 7071 13158 7127 13214
rect 7152 13158 7208 13214
rect 7233 13158 7289 13214
rect 7314 13158 7370 13214
rect 5188 13078 5244 13134
rect 5270 13078 5326 13134
rect 5352 13078 5408 13134
rect 5434 13078 5490 13134
rect 5516 13078 5572 13134
rect 5598 13110 5632 13134
rect 5632 13110 5654 13134
rect 5680 13110 5684 13134
rect 5684 13110 5700 13134
rect 5700 13110 5736 13134
rect 5762 13110 5768 13134
rect 5768 13110 5818 13134
rect 5598 13098 5654 13110
rect 5680 13098 5736 13110
rect 5762 13098 5818 13110
rect 5598 13078 5632 13098
rect 5632 13078 5654 13098
rect 5680 13078 5684 13098
rect 5684 13078 5700 13098
rect 5700 13078 5736 13098
rect 5762 13078 5768 13098
rect 5768 13078 5818 13098
rect 5844 13078 5900 13134
rect 5926 13078 5982 13134
rect 6008 13078 6064 13134
rect 6090 13078 6146 13134
rect 6172 13078 6228 13134
rect 6254 13078 6310 13134
rect 6336 13078 6392 13134
rect 6418 13078 6474 13134
rect 6500 13110 6552 13134
rect 6552 13110 6556 13134
rect 6582 13110 6604 13134
rect 6604 13110 6620 13134
rect 6620 13110 6638 13134
rect 6664 13110 6672 13134
rect 6672 13110 6688 13134
rect 6688 13110 6720 13134
rect 6500 13098 6556 13110
rect 6582 13098 6638 13110
rect 6664 13098 6720 13110
rect 6500 13078 6552 13098
rect 6552 13078 6556 13098
rect 6582 13078 6604 13098
rect 6604 13078 6620 13098
rect 6620 13078 6638 13098
rect 6664 13078 6672 13098
rect 6672 13078 6688 13098
rect 6688 13078 6720 13098
rect 6746 13078 6802 13134
rect 6828 13078 6884 13134
rect 6909 13078 6965 13134
rect 6990 13078 7046 13134
rect 7071 13078 7127 13134
rect 7152 13078 7208 13134
rect 7233 13078 7289 13134
rect 7314 13078 7370 13134
rect 5188 12998 5244 13054
rect 5270 12998 5326 13054
rect 5352 12998 5408 13054
rect 5434 12998 5490 13054
rect 5516 12998 5572 13054
rect 5598 13046 5632 13054
rect 5632 13046 5654 13054
rect 5680 13046 5684 13054
rect 5684 13046 5700 13054
rect 5700 13046 5736 13054
rect 5762 13046 5768 13054
rect 5768 13046 5818 13054
rect 5598 13034 5654 13046
rect 5680 13034 5736 13046
rect 5762 13034 5818 13046
rect 5598 12998 5632 13034
rect 5632 12998 5654 13034
rect 5680 12998 5684 13034
rect 5684 12998 5700 13034
rect 5700 12998 5736 13034
rect 5762 12998 5768 13034
rect 5768 12998 5818 13034
rect 5844 12998 5900 13054
rect 5926 12998 5982 13054
rect 6008 12998 6064 13054
rect 6090 12998 6146 13054
rect 6172 12998 6228 13054
rect 6254 12998 6310 13054
rect 6336 12998 6392 13054
rect 6418 12998 6474 13054
rect 6500 13046 6552 13054
rect 6552 13046 6556 13054
rect 6582 13046 6604 13054
rect 6604 13046 6620 13054
rect 6620 13046 6638 13054
rect 6664 13046 6672 13054
rect 6672 13046 6688 13054
rect 6688 13046 6720 13054
rect 6500 13034 6556 13046
rect 6582 13034 6638 13046
rect 6664 13034 6720 13046
rect 6500 12998 6552 13034
rect 6552 12998 6556 13034
rect 6582 12998 6604 13034
rect 6604 12998 6620 13034
rect 6620 12998 6638 13034
rect 6664 12998 6672 13034
rect 6672 12998 6688 13034
rect 6688 12998 6720 13034
rect 6746 12998 6802 13054
rect 6828 12998 6884 13054
rect 6909 12998 6965 13054
rect 6990 12998 7046 13054
rect 7071 12998 7127 13054
rect 7152 12998 7208 13054
rect 7233 12998 7289 13054
rect 7314 12998 7370 13054
rect 5188 12918 5244 12974
rect 5270 12918 5326 12974
rect 5352 12918 5408 12974
rect 5434 12918 5490 12974
rect 5516 12918 5572 12974
rect 5598 12970 5654 12974
rect 5680 12970 5736 12974
rect 5762 12970 5818 12974
rect 5598 12918 5632 12970
rect 5632 12918 5654 12970
rect 5680 12918 5684 12970
rect 5684 12918 5700 12970
rect 5700 12918 5736 12970
rect 5762 12918 5768 12970
rect 5768 12918 5818 12970
rect 5844 12918 5900 12974
rect 5926 12918 5982 12974
rect 6008 12918 6064 12974
rect 6090 12918 6146 12974
rect 6172 12918 6228 12974
rect 6254 12918 6310 12974
rect 6336 12918 6392 12974
rect 6418 12918 6474 12974
rect 6500 12970 6556 12974
rect 6582 12970 6638 12974
rect 6664 12970 6720 12974
rect 6500 12918 6552 12970
rect 6552 12918 6556 12970
rect 6582 12918 6604 12970
rect 6604 12918 6620 12970
rect 6620 12918 6638 12970
rect 6664 12918 6672 12970
rect 6672 12918 6688 12970
rect 6688 12918 6720 12970
rect 6746 12918 6802 12974
rect 6828 12918 6884 12974
rect 6909 12918 6965 12974
rect 6990 12918 7046 12974
rect 7071 12918 7127 12974
rect 7152 12918 7208 12974
rect 7233 12918 7289 12974
rect 7314 12918 7370 12974
rect 5188 12838 5244 12894
rect 5270 12838 5326 12894
rect 5352 12838 5408 12894
rect 5434 12838 5490 12894
rect 5516 12838 5572 12894
rect 5598 12854 5632 12894
rect 5632 12854 5654 12894
rect 5680 12854 5684 12894
rect 5684 12854 5700 12894
rect 5700 12854 5736 12894
rect 5762 12854 5768 12894
rect 5768 12854 5818 12894
rect 5598 12842 5654 12854
rect 5680 12842 5736 12854
rect 5762 12842 5818 12854
rect 5598 12838 5632 12842
rect 5632 12838 5654 12842
rect 5680 12838 5684 12842
rect 5684 12838 5700 12842
rect 5700 12838 5736 12842
rect 5762 12838 5768 12842
rect 5768 12838 5818 12842
rect 5844 12838 5900 12894
rect 5926 12838 5982 12894
rect 6008 12838 6064 12894
rect 6090 12838 6146 12894
rect 6172 12838 6228 12894
rect 6254 12838 6310 12894
rect 6336 12838 6392 12894
rect 6418 12838 6474 12894
rect 6500 12854 6552 12894
rect 6552 12854 6556 12894
rect 6582 12854 6604 12894
rect 6604 12854 6620 12894
rect 6620 12854 6638 12894
rect 6664 12854 6672 12894
rect 6672 12854 6688 12894
rect 6688 12854 6720 12894
rect 6500 12842 6556 12854
rect 6582 12842 6638 12854
rect 6664 12842 6720 12854
rect 6500 12838 6552 12842
rect 6552 12838 6556 12842
rect 6582 12838 6604 12842
rect 6604 12838 6620 12842
rect 6620 12838 6638 12842
rect 6664 12838 6672 12842
rect 6672 12838 6688 12842
rect 6688 12838 6720 12842
rect 6746 12838 6802 12894
rect 6828 12838 6884 12894
rect 6909 12838 6965 12894
rect 6990 12838 7046 12894
rect 7071 12838 7127 12894
rect 7152 12838 7208 12894
rect 7233 12838 7289 12894
rect 7314 12838 7370 12894
rect 5188 12758 5244 12814
rect 5270 12758 5326 12814
rect 5352 12758 5408 12814
rect 5434 12758 5490 12814
rect 5516 12758 5572 12814
rect 5598 12790 5632 12814
rect 5632 12790 5654 12814
rect 5680 12790 5684 12814
rect 5684 12790 5700 12814
rect 5700 12790 5736 12814
rect 5762 12790 5768 12814
rect 5768 12790 5818 12814
rect 5598 12778 5654 12790
rect 5680 12778 5736 12790
rect 5762 12778 5818 12790
rect 5598 12758 5632 12778
rect 5632 12758 5654 12778
rect 5680 12758 5684 12778
rect 5684 12758 5700 12778
rect 5700 12758 5736 12778
rect 5762 12758 5768 12778
rect 5768 12758 5818 12778
rect 5844 12758 5900 12814
rect 5926 12758 5982 12814
rect 6008 12758 6064 12814
rect 6090 12758 6146 12814
rect 6172 12758 6228 12814
rect 6254 12758 6310 12814
rect 6336 12758 6392 12814
rect 6418 12758 6474 12814
rect 6500 12790 6552 12814
rect 6552 12790 6556 12814
rect 6582 12790 6604 12814
rect 6604 12790 6620 12814
rect 6620 12790 6638 12814
rect 6664 12790 6672 12814
rect 6672 12790 6688 12814
rect 6688 12790 6720 12814
rect 6500 12778 6556 12790
rect 6582 12778 6638 12790
rect 6664 12778 6720 12790
rect 6500 12758 6552 12778
rect 6552 12758 6556 12778
rect 6582 12758 6604 12778
rect 6604 12758 6620 12778
rect 6620 12758 6638 12778
rect 6664 12758 6672 12778
rect 6672 12758 6688 12778
rect 6688 12758 6720 12778
rect 6746 12758 6802 12814
rect 6828 12758 6884 12814
rect 6909 12758 6965 12814
rect 6990 12758 7046 12814
rect 7071 12758 7127 12814
rect 7152 12758 7208 12814
rect 7233 12758 7289 12814
rect 7314 12758 7370 12814
rect 5188 12678 5244 12734
rect 5270 12678 5326 12734
rect 5352 12678 5408 12734
rect 5434 12678 5490 12734
rect 5516 12678 5572 12734
rect 5598 12726 5632 12734
rect 5632 12726 5654 12734
rect 5680 12726 5684 12734
rect 5684 12726 5700 12734
rect 5700 12726 5736 12734
rect 5762 12726 5768 12734
rect 5768 12726 5818 12734
rect 5598 12714 5654 12726
rect 5680 12714 5736 12726
rect 5762 12714 5818 12726
rect 5598 12678 5632 12714
rect 5632 12678 5654 12714
rect 5680 12678 5684 12714
rect 5684 12678 5700 12714
rect 5700 12678 5736 12714
rect 5762 12678 5768 12714
rect 5768 12678 5818 12714
rect 5844 12678 5900 12734
rect 5926 12678 5982 12734
rect 6008 12678 6064 12734
rect 6090 12678 6146 12734
rect 6172 12678 6228 12734
rect 6254 12678 6310 12734
rect 6336 12678 6392 12734
rect 6418 12678 6474 12734
rect 6500 12726 6552 12734
rect 6552 12726 6556 12734
rect 6582 12726 6604 12734
rect 6604 12726 6620 12734
rect 6620 12726 6638 12734
rect 6664 12726 6672 12734
rect 6672 12726 6688 12734
rect 6688 12726 6720 12734
rect 6500 12714 6556 12726
rect 6582 12714 6638 12726
rect 6664 12714 6720 12726
rect 6500 12678 6552 12714
rect 6552 12678 6556 12714
rect 6582 12678 6604 12714
rect 6604 12678 6620 12714
rect 6620 12678 6638 12714
rect 6664 12678 6672 12714
rect 6672 12678 6688 12714
rect 6688 12678 6720 12714
rect 6746 12678 6802 12734
rect 6828 12678 6884 12734
rect 6909 12678 6965 12734
rect 6990 12678 7046 12734
rect 7071 12678 7127 12734
rect 7152 12678 7208 12734
rect 7233 12678 7289 12734
rect 7314 12678 7370 12734
rect 5188 12598 5244 12654
rect 5270 12598 5326 12654
rect 5352 12598 5408 12654
rect 5434 12598 5490 12654
rect 5516 12598 5572 12654
rect 5598 12650 5654 12654
rect 5680 12650 5736 12654
rect 5762 12650 5818 12654
rect 5598 12598 5632 12650
rect 5632 12598 5654 12650
rect 5680 12598 5684 12650
rect 5684 12598 5700 12650
rect 5700 12598 5736 12650
rect 5762 12598 5768 12650
rect 5768 12598 5818 12650
rect 5844 12598 5900 12654
rect 5926 12598 5982 12654
rect 6008 12598 6064 12654
rect 6090 12598 6146 12654
rect 6172 12598 6228 12654
rect 6254 12598 6310 12654
rect 6336 12598 6392 12654
rect 6418 12598 6474 12654
rect 6500 12650 6556 12654
rect 6582 12650 6638 12654
rect 6664 12650 6720 12654
rect 6500 12598 6552 12650
rect 6552 12598 6556 12650
rect 6582 12598 6604 12650
rect 6604 12598 6620 12650
rect 6620 12598 6638 12650
rect 6664 12598 6672 12650
rect 6672 12598 6688 12650
rect 6688 12598 6720 12650
rect 6746 12598 6802 12654
rect 6828 12598 6884 12654
rect 6909 12598 6965 12654
rect 6990 12598 7046 12654
rect 7071 12598 7127 12654
rect 7152 12598 7208 12654
rect 7233 12598 7289 12654
rect 7314 12598 7370 12654
rect 5188 12518 5244 12574
rect 5270 12518 5326 12574
rect 5352 12518 5408 12574
rect 5434 12518 5490 12574
rect 5516 12518 5572 12574
rect 5598 12534 5632 12574
rect 5632 12534 5654 12574
rect 5680 12534 5684 12574
rect 5684 12534 5700 12574
rect 5700 12534 5736 12574
rect 5762 12534 5768 12574
rect 5768 12534 5818 12574
rect 5598 12522 5654 12534
rect 5680 12522 5736 12534
rect 5762 12522 5818 12534
rect 5598 12518 5632 12522
rect 5632 12518 5654 12522
rect 5680 12518 5684 12522
rect 5684 12518 5700 12522
rect 5700 12518 5736 12522
rect 5762 12518 5768 12522
rect 5768 12518 5818 12522
rect 5844 12518 5900 12574
rect 5926 12518 5982 12574
rect 6008 12518 6064 12574
rect 6090 12518 6146 12574
rect 6172 12518 6228 12574
rect 6254 12518 6310 12574
rect 6336 12518 6392 12574
rect 6418 12518 6474 12574
rect 6500 12534 6552 12574
rect 6552 12534 6556 12574
rect 6582 12534 6604 12574
rect 6604 12534 6620 12574
rect 6620 12534 6638 12574
rect 6664 12534 6672 12574
rect 6672 12534 6688 12574
rect 6688 12534 6720 12574
rect 6500 12522 6556 12534
rect 6582 12522 6638 12534
rect 6664 12522 6720 12534
rect 6500 12518 6552 12522
rect 6552 12518 6556 12522
rect 6582 12518 6604 12522
rect 6604 12518 6620 12522
rect 6620 12518 6638 12522
rect 6664 12518 6672 12522
rect 6672 12518 6688 12522
rect 6688 12518 6720 12522
rect 6746 12518 6802 12574
rect 6828 12518 6884 12574
rect 6909 12518 6965 12574
rect 6990 12518 7046 12574
rect 7071 12518 7127 12574
rect 7152 12518 7208 12574
rect 7233 12518 7289 12574
rect 7314 12518 7370 12574
rect 5188 12438 5244 12494
rect 5270 12438 5326 12494
rect 5352 12438 5408 12494
rect 5434 12438 5490 12494
rect 5516 12438 5572 12494
rect 5598 12470 5632 12494
rect 5632 12470 5654 12494
rect 5680 12470 5684 12494
rect 5684 12470 5700 12494
rect 5700 12470 5736 12494
rect 5762 12470 5768 12494
rect 5768 12470 5818 12494
rect 5598 12458 5654 12470
rect 5680 12458 5736 12470
rect 5762 12458 5818 12470
rect 5598 12438 5632 12458
rect 5632 12438 5654 12458
rect 5680 12438 5684 12458
rect 5684 12438 5700 12458
rect 5700 12438 5736 12458
rect 5762 12438 5768 12458
rect 5768 12438 5818 12458
rect 5844 12438 5900 12494
rect 5926 12438 5982 12494
rect 6008 12438 6064 12494
rect 6090 12438 6146 12494
rect 6172 12438 6228 12494
rect 6254 12438 6310 12494
rect 6336 12438 6392 12494
rect 6418 12438 6474 12494
rect 6500 12470 6552 12494
rect 6552 12470 6556 12494
rect 6582 12470 6604 12494
rect 6604 12470 6620 12494
rect 6620 12470 6638 12494
rect 6664 12470 6672 12494
rect 6672 12470 6688 12494
rect 6688 12470 6720 12494
rect 6500 12458 6556 12470
rect 6582 12458 6638 12470
rect 6664 12458 6720 12470
rect 6500 12438 6552 12458
rect 6552 12438 6556 12458
rect 6582 12438 6604 12458
rect 6604 12438 6620 12458
rect 6620 12438 6638 12458
rect 6664 12438 6672 12458
rect 6672 12438 6688 12458
rect 6688 12438 6720 12458
rect 6746 12438 6802 12494
rect 6828 12438 6884 12494
rect 6909 12438 6965 12494
rect 6990 12438 7046 12494
rect 7071 12438 7127 12494
rect 7152 12438 7208 12494
rect 7233 12438 7289 12494
rect 7314 12438 7370 12494
rect 5188 12358 5244 12414
rect 5270 12358 5326 12414
rect 5352 12358 5408 12414
rect 5434 12358 5490 12414
rect 5516 12358 5572 12414
rect 5598 12406 5632 12414
rect 5632 12406 5654 12414
rect 5680 12406 5684 12414
rect 5684 12406 5700 12414
rect 5700 12406 5736 12414
rect 5762 12406 5768 12414
rect 5768 12406 5818 12414
rect 5598 12394 5654 12406
rect 5680 12394 5736 12406
rect 5762 12394 5818 12406
rect 5598 12358 5632 12394
rect 5632 12358 5654 12394
rect 5680 12358 5684 12394
rect 5684 12358 5700 12394
rect 5700 12358 5736 12394
rect 5762 12358 5768 12394
rect 5768 12358 5818 12394
rect 5844 12358 5900 12414
rect 5926 12358 5982 12414
rect 6008 12358 6064 12414
rect 6090 12358 6146 12414
rect 6172 12358 6228 12414
rect 6254 12358 6310 12414
rect 6336 12358 6392 12414
rect 6418 12358 6474 12414
rect 6500 12406 6552 12414
rect 6552 12406 6556 12414
rect 6582 12406 6604 12414
rect 6604 12406 6620 12414
rect 6620 12406 6638 12414
rect 6664 12406 6672 12414
rect 6672 12406 6688 12414
rect 6688 12406 6720 12414
rect 6500 12394 6556 12406
rect 6582 12394 6638 12406
rect 6664 12394 6720 12406
rect 6500 12358 6552 12394
rect 6552 12358 6556 12394
rect 6582 12358 6604 12394
rect 6604 12358 6620 12394
rect 6620 12358 6638 12394
rect 6664 12358 6672 12394
rect 6672 12358 6688 12394
rect 6688 12358 6720 12394
rect 6746 12358 6802 12414
rect 6828 12358 6884 12414
rect 6909 12358 6965 12414
rect 6990 12358 7046 12414
rect 7071 12358 7127 12414
rect 7152 12358 7208 12414
rect 7233 12358 7289 12414
rect 7314 12358 7370 12414
rect 5188 12278 5244 12334
rect 5270 12278 5326 12334
rect 5352 12278 5408 12334
rect 5434 12278 5490 12334
rect 5516 12278 5572 12334
rect 5598 12329 5654 12334
rect 5680 12329 5736 12334
rect 5762 12329 5818 12334
rect 5598 12278 5632 12329
rect 5632 12278 5654 12329
rect 5680 12278 5684 12329
rect 5684 12278 5700 12329
rect 5700 12278 5736 12329
rect 5762 12278 5768 12329
rect 5768 12278 5818 12329
rect 5844 12278 5900 12334
rect 5926 12278 5982 12334
rect 6008 12278 6064 12334
rect 6090 12278 6146 12334
rect 6172 12278 6228 12334
rect 6254 12278 6310 12334
rect 6336 12278 6392 12334
rect 6418 12278 6474 12334
rect 6500 12329 6556 12334
rect 6582 12329 6638 12334
rect 6664 12329 6720 12334
rect 6500 12278 6552 12329
rect 6552 12278 6556 12329
rect 6582 12278 6604 12329
rect 6604 12278 6620 12329
rect 6620 12278 6638 12329
rect 6664 12278 6672 12329
rect 6672 12278 6688 12329
rect 6688 12278 6720 12329
rect 6746 12278 6802 12334
rect 6828 12278 6884 12334
rect 6909 12278 6965 12334
rect 6990 12278 7046 12334
rect 7071 12278 7127 12334
rect 7152 12278 7208 12334
rect 7233 12278 7289 12334
rect 7314 12278 7370 12334
rect 5188 12198 5244 12254
rect 5270 12198 5326 12254
rect 5352 12198 5408 12254
rect 5434 12198 5490 12254
rect 5516 12198 5572 12254
rect 5598 12212 5632 12254
rect 5632 12212 5654 12254
rect 5680 12212 5684 12254
rect 5684 12212 5700 12254
rect 5700 12212 5736 12254
rect 5762 12212 5768 12254
rect 5768 12212 5818 12254
rect 5598 12199 5654 12212
rect 5680 12199 5736 12212
rect 5762 12199 5818 12212
rect 5598 12198 5632 12199
rect 5632 12198 5654 12199
rect 5680 12198 5684 12199
rect 5684 12198 5700 12199
rect 5700 12198 5736 12199
rect 5762 12198 5768 12199
rect 5768 12198 5818 12199
rect 5844 12198 5900 12254
rect 5926 12198 5982 12254
rect 6008 12198 6064 12254
rect 6090 12198 6146 12254
rect 6172 12198 6228 12254
rect 6254 12198 6310 12254
rect 6336 12198 6392 12254
rect 6418 12198 6474 12254
rect 6500 12212 6552 12254
rect 6552 12212 6556 12254
rect 6582 12212 6604 12254
rect 6604 12212 6620 12254
rect 6620 12212 6638 12254
rect 6664 12212 6672 12254
rect 6672 12212 6688 12254
rect 6688 12212 6720 12254
rect 6500 12199 6556 12212
rect 6582 12199 6638 12212
rect 6664 12199 6720 12212
rect 6500 12198 6552 12199
rect 6552 12198 6556 12199
rect 6582 12198 6604 12199
rect 6604 12198 6620 12199
rect 6620 12198 6638 12199
rect 6664 12198 6672 12199
rect 6672 12198 6688 12199
rect 6688 12198 6720 12199
rect 6746 12198 6802 12254
rect 6828 12198 6884 12254
rect 6909 12198 6965 12254
rect 6990 12198 7046 12254
rect 7071 12198 7127 12254
rect 7152 12198 7208 12254
rect 7233 12198 7289 12254
rect 7314 12198 7370 12254
rect 5188 12118 5244 12174
rect 5270 12118 5326 12174
rect 5352 12118 5408 12174
rect 5434 12118 5490 12174
rect 5516 12118 5572 12174
rect 5598 12147 5632 12174
rect 5632 12147 5654 12174
rect 5680 12147 5684 12174
rect 5684 12147 5700 12174
rect 5700 12147 5736 12174
rect 5762 12147 5768 12174
rect 5768 12147 5818 12174
rect 5598 12134 5654 12147
rect 5680 12134 5736 12147
rect 5762 12134 5818 12147
rect 5598 12118 5632 12134
rect 5632 12118 5654 12134
rect 5680 12118 5684 12134
rect 5684 12118 5700 12134
rect 5700 12118 5736 12134
rect 5762 12118 5768 12134
rect 5768 12118 5818 12134
rect 5844 12118 5900 12174
rect 5926 12118 5982 12174
rect 6008 12118 6064 12174
rect 6090 12118 6146 12174
rect 6172 12118 6228 12174
rect 6254 12118 6310 12174
rect 6336 12118 6392 12174
rect 6418 12118 6474 12174
rect 6500 12147 6552 12174
rect 6552 12147 6556 12174
rect 6582 12147 6604 12174
rect 6604 12147 6620 12174
rect 6620 12147 6638 12174
rect 6664 12147 6672 12174
rect 6672 12147 6688 12174
rect 6688 12147 6720 12174
rect 6500 12134 6556 12147
rect 6582 12134 6638 12147
rect 6664 12134 6720 12147
rect 6500 12118 6552 12134
rect 6552 12118 6556 12134
rect 6582 12118 6604 12134
rect 6604 12118 6620 12134
rect 6620 12118 6638 12134
rect 6664 12118 6672 12134
rect 6672 12118 6688 12134
rect 6688 12118 6720 12134
rect 6746 12118 6802 12174
rect 6828 12118 6884 12174
rect 6909 12118 6965 12174
rect 6990 12118 7046 12174
rect 7071 12118 7127 12174
rect 7152 12118 7208 12174
rect 7233 12118 7289 12174
rect 7314 12118 7370 12174
rect 5188 12038 5244 12094
rect 5270 12038 5326 12094
rect 5352 12038 5408 12094
rect 5434 12038 5490 12094
rect 5516 12038 5572 12094
rect 5598 12082 5632 12094
rect 5632 12082 5654 12094
rect 5680 12082 5684 12094
rect 5684 12082 5700 12094
rect 5700 12082 5736 12094
rect 5762 12082 5768 12094
rect 5768 12082 5818 12094
rect 5598 12069 5654 12082
rect 5680 12069 5736 12082
rect 5762 12069 5818 12082
rect 5598 12038 5632 12069
rect 5632 12038 5654 12069
rect 5680 12038 5684 12069
rect 5684 12038 5700 12069
rect 5700 12038 5736 12069
rect 5762 12038 5768 12069
rect 5768 12038 5818 12069
rect 5844 12038 5900 12094
rect 5926 12038 5982 12094
rect 6008 12038 6064 12094
rect 6090 12038 6146 12094
rect 6172 12038 6228 12094
rect 6254 12038 6310 12094
rect 6336 12038 6392 12094
rect 6418 12038 6474 12094
rect 6500 12082 6552 12094
rect 6552 12082 6556 12094
rect 6582 12082 6604 12094
rect 6604 12082 6620 12094
rect 6620 12082 6638 12094
rect 6664 12082 6672 12094
rect 6672 12082 6688 12094
rect 6688 12082 6720 12094
rect 6500 12069 6556 12082
rect 6582 12069 6638 12082
rect 6664 12069 6720 12082
rect 6500 12038 6552 12069
rect 6552 12038 6556 12069
rect 6582 12038 6604 12069
rect 6604 12038 6620 12069
rect 6620 12038 6638 12069
rect 6664 12038 6672 12069
rect 6672 12038 6688 12069
rect 6688 12038 6720 12069
rect 6746 12038 6802 12094
rect 6828 12038 6884 12094
rect 6909 12038 6965 12094
rect 6990 12038 7046 12094
rect 7071 12038 7127 12094
rect 7152 12038 7208 12094
rect 7233 12038 7289 12094
rect 7314 12038 7370 12094
rect 5188 11958 5244 12014
rect 5270 11958 5326 12014
rect 5352 11958 5408 12014
rect 5434 11958 5490 12014
rect 5516 11958 5572 12014
rect 5598 12004 5654 12014
rect 5680 12004 5736 12014
rect 5762 12004 5818 12014
rect 5598 11958 5632 12004
rect 5632 11958 5654 12004
rect 5680 11958 5684 12004
rect 5684 11958 5700 12004
rect 5700 11958 5736 12004
rect 5762 11958 5768 12004
rect 5768 11958 5818 12004
rect 5844 11958 5900 12014
rect 5926 11958 5982 12014
rect 6008 11958 6064 12014
rect 6090 11958 6146 12014
rect 6172 11958 6228 12014
rect 6254 11958 6310 12014
rect 6336 11958 6392 12014
rect 6418 11958 6474 12014
rect 6500 12004 6556 12014
rect 6582 12004 6638 12014
rect 6664 12004 6720 12014
rect 6500 11958 6552 12004
rect 6552 11958 6556 12004
rect 6582 11958 6604 12004
rect 6604 11958 6620 12004
rect 6620 11958 6638 12004
rect 6664 11958 6672 12004
rect 6672 11958 6688 12004
rect 6688 11958 6720 12004
rect 6746 11958 6802 12014
rect 6828 11958 6884 12014
rect 6909 11958 6965 12014
rect 6990 11958 7046 12014
rect 7071 11958 7127 12014
rect 7152 11958 7208 12014
rect 7233 11958 7289 12014
rect 7314 11958 7370 12014
rect 5188 11878 5244 11934
rect 5270 11878 5326 11934
rect 5352 11878 5408 11934
rect 5434 11878 5490 11934
rect 5516 11878 5572 11934
rect 5598 11887 5632 11934
rect 5632 11887 5654 11934
rect 5680 11887 5684 11934
rect 5684 11887 5700 11934
rect 5700 11887 5736 11934
rect 5762 11887 5768 11934
rect 5768 11887 5818 11934
rect 5598 11878 5654 11887
rect 5680 11878 5736 11887
rect 5762 11878 5818 11887
rect 5844 11878 5900 11934
rect 5926 11878 5982 11934
rect 6008 11878 6064 11934
rect 6090 11878 6146 11934
rect 6172 11878 6228 11934
rect 6254 11878 6310 11934
rect 6336 11878 6392 11934
rect 6418 11878 6474 11934
rect 6500 11887 6552 11934
rect 6552 11887 6556 11934
rect 6582 11887 6604 11934
rect 6604 11887 6620 11934
rect 6620 11887 6638 11934
rect 6664 11887 6672 11934
rect 6672 11887 6688 11934
rect 6688 11887 6720 11934
rect 6500 11878 6556 11887
rect 6582 11878 6638 11887
rect 6664 11878 6720 11887
rect 6746 11878 6802 11934
rect 6828 11878 6884 11934
rect 6909 11878 6965 11934
rect 6990 11878 7046 11934
rect 7071 11878 7127 11934
rect 7152 11878 7208 11934
rect 7233 11878 7289 11934
rect 7314 11878 7370 11934
rect 5188 11798 5244 11854
rect 5270 11798 5326 11854
rect 5352 11798 5408 11854
rect 5434 11798 5490 11854
rect 5516 11798 5572 11854
rect 5598 11822 5632 11854
rect 5632 11822 5654 11854
rect 5680 11822 5684 11854
rect 5684 11822 5700 11854
rect 5700 11822 5736 11854
rect 5762 11822 5768 11854
rect 5768 11822 5818 11854
rect 5598 11809 5654 11822
rect 5680 11809 5736 11822
rect 5762 11809 5818 11822
rect 5598 11798 5632 11809
rect 5632 11798 5654 11809
rect 5680 11798 5684 11809
rect 5684 11798 5700 11809
rect 5700 11798 5736 11809
rect 5762 11798 5768 11809
rect 5768 11798 5818 11809
rect 5844 11798 5900 11854
rect 5926 11798 5982 11854
rect 6008 11798 6064 11854
rect 6090 11798 6146 11854
rect 6172 11798 6228 11854
rect 6254 11798 6310 11854
rect 6336 11798 6392 11854
rect 6418 11798 6474 11854
rect 6500 11822 6552 11854
rect 6552 11822 6556 11854
rect 6582 11822 6604 11854
rect 6604 11822 6620 11854
rect 6620 11822 6638 11854
rect 6664 11822 6672 11854
rect 6672 11822 6688 11854
rect 6688 11822 6720 11854
rect 6500 11809 6556 11822
rect 6582 11809 6638 11822
rect 6664 11809 6720 11822
rect 6500 11798 6552 11809
rect 6552 11798 6556 11809
rect 6582 11798 6604 11809
rect 6604 11798 6620 11809
rect 6620 11798 6638 11809
rect 6664 11798 6672 11809
rect 6672 11798 6688 11809
rect 6688 11798 6720 11809
rect 6746 11798 6802 11854
rect 6828 11798 6884 11854
rect 6909 11798 6965 11854
rect 6990 11798 7046 11854
rect 7071 11798 7127 11854
rect 7152 11798 7208 11854
rect 7233 11798 7289 11854
rect 7314 11798 7370 11854
rect 5188 11718 5244 11774
rect 5270 11718 5326 11774
rect 5352 11718 5408 11774
rect 5434 11718 5490 11774
rect 5516 11718 5572 11774
rect 5598 11757 5632 11774
rect 5632 11757 5654 11774
rect 5680 11757 5684 11774
rect 5684 11757 5700 11774
rect 5700 11757 5736 11774
rect 5762 11757 5768 11774
rect 5768 11757 5818 11774
rect 5598 11744 5654 11757
rect 5680 11744 5736 11757
rect 5762 11744 5818 11757
rect 5598 11718 5632 11744
rect 5632 11718 5654 11744
rect 5680 11718 5684 11744
rect 5684 11718 5700 11744
rect 5700 11718 5736 11744
rect 5762 11718 5768 11744
rect 5768 11718 5818 11744
rect 5844 11718 5900 11774
rect 5926 11718 5982 11774
rect 6008 11718 6064 11774
rect 6090 11718 6146 11774
rect 6172 11718 6228 11774
rect 6254 11718 6310 11774
rect 6336 11718 6392 11774
rect 6418 11718 6474 11774
rect 6500 11757 6552 11774
rect 6552 11757 6556 11774
rect 6582 11757 6604 11774
rect 6604 11757 6620 11774
rect 6620 11757 6638 11774
rect 6664 11757 6672 11774
rect 6672 11757 6688 11774
rect 6688 11757 6720 11774
rect 6500 11744 6556 11757
rect 6582 11744 6638 11757
rect 6664 11744 6720 11757
rect 6500 11718 6552 11744
rect 6552 11718 6556 11744
rect 6582 11718 6604 11744
rect 6604 11718 6620 11744
rect 6620 11718 6638 11744
rect 6664 11718 6672 11744
rect 6672 11718 6688 11744
rect 6688 11718 6720 11744
rect 6746 11718 6802 11774
rect 6828 11718 6884 11774
rect 6909 11718 6965 11774
rect 6990 11718 7046 11774
rect 7071 11718 7127 11774
rect 7152 11718 7208 11774
rect 7233 11718 7289 11774
rect 7314 11718 7370 11774
rect 5188 11638 5244 11694
rect 5270 11638 5326 11694
rect 5352 11638 5408 11694
rect 5434 11638 5490 11694
rect 5516 11638 5572 11694
rect 5598 11692 5632 11694
rect 5632 11692 5654 11694
rect 5680 11692 5684 11694
rect 5684 11692 5700 11694
rect 5700 11692 5736 11694
rect 5762 11692 5768 11694
rect 5768 11692 5818 11694
rect 5598 11679 5654 11692
rect 5680 11679 5736 11692
rect 5762 11679 5818 11692
rect 5598 11638 5632 11679
rect 5632 11638 5654 11679
rect 5680 11638 5684 11679
rect 5684 11638 5700 11679
rect 5700 11638 5736 11679
rect 5762 11638 5768 11679
rect 5768 11638 5818 11679
rect 5844 11638 5900 11694
rect 5926 11638 5982 11694
rect 6008 11638 6064 11694
rect 6090 11638 6146 11694
rect 6172 11638 6228 11694
rect 6254 11638 6310 11694
rect 6336 11638 6392 11694
rect 6418 11638 6474 11694
rect 6500 11692 6552 11694
rect 6552 11692 6556 11694
rect 6582 11692 6604 11694
rect 6604 11692 6620 11694
rect 6620 11692 6638 11694
rect 6664 11692 6672 11694
rect 6672 11692 6688 11694
rect 6688 11692 6720 11694
rect 6500 11679 6556 11692
rect 6582 11679 6638 11692
rect 6664 11679 6720 11692
rect 6500 11638 6552 11679
rect 6552 11638 6556 11679
rect 6582 11638 6604 11679
rect 6604 11638 6620 11679
rect 6620 11638 6638 11679
rect 6664 11638 6672 11679
rect 6672 11638 6688 11679
rect 6688 11638 6720 11679
rect 6746 11638 6802 11694
rect 6828 11638 6884 11694
rect 6909 11638 6965 11694
rect 6990 11638 7046 11694
rect 7071 11638 7127 11694
rect 7152 11638 7208 11694
rect 7233 11638 7289 11694
rect 7314 11638 7370 11694
rect 5188 11558 5244 11614
rect 5270 11558 5326 11614
rect 5352 11558 5408 11614
rect 5434 11558 5490 11614
rect 5516 11558 5572 11614
rect 5598 11562 5632 11614
rect 5632 11562 5654 11614
rect 5680 11562 5684 11614
rect 5684 11562 5700 11614
rect 5700 11562 5736 11614
rect 5762 11562 5768 11614
rect 5768 11562 5818 11614
rect 5598 11558 5654 11562
rect 5680 11558 5736 11562
rect 5762 11558 5818 11562
rect 5844 11558 5900 11614
rect 5926 11558 5982 11614
rect 6008 11558 6064 11614
rect 6090 11558 6146 11614
rect 6172 11558 6228 11614
rect 6254 11558 6310 11614
rect 6336 11558 6392 11614
rect 6418 11558 6474 11614
rect 6500 11562 6552 11614
rect 6552 11562 6556 11614
rect 6582 11562 6604 11614
rect 6604 11562 6620 11614
rect 6620 11562 6638 11614
rect 6664 11562 6672 11614
rect 6672 11562 6688 11614
rect 6688 11562 6720 11614
rect 6500 11558 6556 11562
rect 6582 11558 6638 11562
rect 6664 11558 6720 11562
rect 6746 11558 6802 11614
rect 6828 11558 6884 11614
rect 6909 11558 6965 11614
rect 6990 11558 7046 11614
rect 7071 11558 7127 11614
rect 7152 11558 7208 11614
rect 7233 11558 7289 11614
rect 7314 11558 7370 11614
rect 7587 11173 7643 11229
rect 7669 11173 7725 11229
rect 7751 11173 7807 11229
rect 7833 11173 7889 11229
rect 7915 11225 7971 11229
rect 7997 11225 8053 11229
rect 8079 11225 8135 11229
rect 7915 11173 7961 11225
rect 7961 11173 7971 11225
rect 7997 11173 8013 11225
rect 8013 11173 8039 11225
rect 8039 11173 8053 11225
rect 8079 11173 8091 11225
rect 8091 11173 8135 11225
rect 8161 11173 8217 11229
rect 8243 11173 8299 11229
rect 8325 11173 8381 11229
rect 8407 11173 8463 11229
rect 8489 11173 8545 11229
rect 8571 11173 8627 11229
rect 8653 11173 8709 11229
rect 8735 11173 8791 11229
rect 8817 11173 8873 11229
rect 8899 11225 8955 11229
rect 8981 11225 9037 11229
rect 8899 11173 8933 11225
rect 8933 11173 8955 11225
rect 8981 11173 9011 11225
rect 9011 11173 9037 11225
rect 9063 11173 9119 11229
rect 9145 11173 9201 11229
rect 9227 11173 9283 11229
rect 9308 11173 9364 11229
rect 9389 11173 9445 11229
rect 9470 11173 9526 11229
rect 9551 11173 9607 11229
rect 9632 11173 9688 11229
rect 9713 11173 9769 11229
rect 7587 11093 7643 11149
rect 7669 11093 7725 11149
rect 7751 11093 7807 11149
rect 7833 11093 7889 11149
rect 7915 11109 7961 11149
rect 7961 11109 7971 11149
rect 7997 11109 8013 11149
rect 8013 11109 8039 11149
rect 8039 11109 8053 11149
rect 8079 11109 8091 11149
rect 8091 11109 8135 11149
rect 7915 11097 7971 11109
rect 7997 11097 8053 11109
rect 8079 11097 8135 11109
rect 7915 11093 7961 11097
rect 7961 11093 7971 11097
rect 7997 11093 8013 11097
rect 8013 11093 8039 11097
rect 8039 11093 8053 11097
rect 8079 11093 8091 11097
rect 8091 11093 8135 11097
rect 8161 11093 8217 11149
rect 8243 11093 8299 11149
rect 8325 11093 8381 11149
rect 8407 11093 8463 11149
rect 8489 11093 8545 11149
rect 8571 11093 8627 11149
rect 8653 11093 8709 11149
rect 8735 11093 8791 11149
rect 8817 11093 8873 11149
rect 8899 11109 8933 11149
rect 8933 11109 8955 11149
rect 8981 11109 9011 11149
rect 9011 11109 9037 11149
rect 8899 11097 8955 11109
rect 8981 11097 9037 11109
rect 8899 11093 8933 11097
rect 8933 11093 8955 11097
rect 8981 11093 9011 11097
rect 9011 11093 9037 11097
rect 9063 11093 9119 11149
rect 9145 11093 9201 11149
rect 9227 11093 9283 11149
rect 9308 11093 9364 11149
rect 9389 11093 9445 11149
rect 9470 11093 9526 11149
rect 9551 11093 9607 11149
rect 9632 11093 9688 11149
rect 9713 11093 9769 11149
rect 7587 11013 7643 11069
rect 7669 11013 7725 11069
rect 7751 11013 7807 11069
rect 7833 11013 7889 11069
rect 7915 11045 7961 11069
rect 7961 11045 7971 11069
rect 7997 11045 8013 11069
rect 8013 11045 8039 11069
rect 8039 11045 8053 11069
rect 8079 11045 8091 11069
rect 8091 11045 8135 11069
rect 7915 11033 7971 11045
rect 7997 11033 8053 11045
rect 8079 11033 8135 11045
rect 7915 11013 7961 11033
rect 7961 11013 7971 11033
rect 7997 11013 8013 11033
rect 8013 11013 8039 11033
rect 8039 11013 8053 11033
rect 8079 11013 8091 11033
rect 8091 11013 8135 11033
rect 8161 11013 8217 11069
rect 8243 11013 8299 11069
rect 8325 11013 8381 11069
rect 8407 11013 8463 11069
rect 8489 11013 8545 11069
rect 8571 11013 8627 11069
rect 8653 11013 8709 11069
rect 8735 11013 8791 11069
rect 8817 11013 8873 11069
rect 8899 11045 8933 11069
rect 8933 11045 8955 11069
rect 8981 11045 9011 11069
rect 9011 11045 9037 11069
rect 8899 11033 8955 11045
rect 8981 11033 9037 11045
rect 8899 11013 8933 11033
rect 8933 11013 8955 11033
rect 8981 11013 9011 11033
rect 9011 11013 9037 11033
rect 9063 11013 9119 11069
rect 9145 11013 9201 11069
rect 9227 11013 9283 11069
rect 9308 11013 9364 11069
rect 9389 11013 9445 11069
rect 9470 11013 9526 11069
rect 9551 11013 9607 11069
rect 9632 11013 9688 11069
rect 9713 11013 9769 11069
rect 7587 10933 7643 10989
rect 7669 10933 7725 10989
rect 7751 10933 7807 10989
rect 7833 10933 7889 10989
rect 7915 10981 7961 10989
rect 7961 10981 7971 10989
rect 7997 10981 8013 10989
rect 8013 10981 8039 10989
rect 8039 10981 8053 10989
rect 8079 10981 8091 10989
rect 8091 10981 8135 10989
rect 7915 10969 7971 10981
rect 7997 10969 8053 10981
rect 8079 10969 8135 10981
rect 7915 10933 7961 10969
rect 7961 10933 7971 10969
rect 7997 10933 8013 10969
rect 8013 10933 8039 10969
rect 8039 10933 8053 10969
rect 8079 10933 8091 10969
rect 8091 10933 8135 10969
rect 8161 10933 8217 10989
rect 8243 10933 8299 10989
rect 8325 10933 8381 10989
rect 8407 10933 8463 10989
rect 8489 10933 8545 10989
rect 8571 10933 8627 10989
rect 8653 10933 8709 10989
rect 8735 10933 8791 10989
rect 8817 10933 8873 10989
rect 8899 10981 8933 10989
rect 8933 10981 8955 10989
rect 8981 10981 9011 10989
rect 9011 10981 9037 10989
rect 8899 10969 8955 10981
rect 8981 10969 9037 10981
rect 8899 10933 8933 10969
rect 8933 10933 8955 10969
rect 8981 10933 9011 10969
rect 9011 10933 9037 10969
rect 9063 10933 9119 10989
rect 9145 10933 9201 10989
rect 9227 10933 9283 10989
rect 9308 10933 9364 10989
rect 9389 10933 9445 10989
rect 9470 10933 9526 10989
rect 9551 10933 9607 10989
rect 9632 10933 9688 10989
rect 9713 10933 9769 10989
rect 7587 10853 7643 10909
rect 7669 10853 7725 10909
rect 7751 10853 7807 10909
rect 7833 10853 7889 10909
rect 7915 10905 7971 10909
rect 7997 10905 8053 10909
rect 8079 10905 8135 10909
rect 7915 10853 7961 10905
rect 7961 10853 7971 10905
rect 7997 10853 8013 10905
rect 8013 10853 8039 10905
rect 8039 10853 8053 10905
rect 8079 10853 8091 10905
rect 8091 10853 8135 10905
rect 8161 10853 8217 10909
rect 8243 10853 8299 10909
rect 8325 10853 8381 10909
rect 8407 10853 8463 10909
rect 8489 10853 8545 10909
rect 8571 10853 8627 10909
rect 8653 10853 8709 10909
rect 8735 10853 8791 10909
rect 8817 10853 8873 10909
rect 8899 10905 8955 10909
rect 8981 10905 9037 10909
rect 8899 10853 8933 10905
rect 8933 10853 8955 10905
rect 8981 10853 9011 10905
rect 9011 10853 9037 10905
rect 9063 10853 9119 10909
rect 9145 10853 9201 10909
rect 9227 10853 9283 10909
rect 9308 10853 9364 10909
rect 9389 10853 9445 10909
rect 9470 10853 9526 10909
rect 9551 10853 9607 10909
rect 9632 10853 9688 10909
rect 9713 10853 9769 10909
rect 7587 10773 7643 10829
rect 7669 10773 7725 10829
rect 7751 10773 7807 10829
rect 7833 10773 7889 10829
rect 7915 10789 7961 10829
rect 7961 10789 7971 10829
rect 7997 10789 8013 10829
rect 8013 10789 8039 10829
rect 8039 10789 8053 10829
rect 8079 10789 8091 10829
rect 8091 10789 8135 10829
rect 7915 10777 7971 10789
rect 7997 10777 8053 10789
rect 8079 10777 8135 10789
rect 7915 10773 7961 10777
rect 7961 10773 7971 10777
rect 7997 10773 8013 10777
rect 8013 10773 8039 10777
rect 8039 10773 8053 10777
rect 8079 10773 8091 10777
rect 8091 10773 8135 10777
rect 8161 10773 8217 10829
rect 8243 10773 8299 10829
rect 8325 10773 8381 10829
rect 8407 10773 8463 10829
rect 8489 10773 8545 10829
rect 8571 10773 8627 10829
rect 8653 10773 8709 10829
rect 8735 10773 8791 10829
rect 8817 10773 8873 10829
rect 8899 10789 8933 10829
rect 8933 10789 8955 10829
rect 8981 10789 9011 10829
rect 9011 10789 9037 10829
rect 8899 10777 8955 10789
rect 8981 10777 9037 10789
rect 8899 10773 8933 10777
rect 8933 10773 8955 10777
rect 8981 10773 9011 10777
rect 9011 10773 9037 10777
rect 9063 10773 9119 10829
rect 9145 10773 9201 10829
rect 9227 10773 9283 10829
rect 9308 10773 9364 10829
rect 9389 10773 9445 10829
rect 9470 10773 9526 10829
rect 9551 10773 9607 10829
rect 9632 10773 9688 10829
rect 9713 10773 9769 10829
rect 7587 10693 7643 10749
rect 7669 10693 7725 10749
rect 7751 10693 7807 10749
rect 7833 10693 7889 10749
rect 7915 10725 7961 10749
rect 7961 10725 7971 10749
rect 7997 10725 8013 10749
rect 8013 10725 8039 10749
rect 8039 10725 8053 10749
rect 8079 10725 8091 10749
rect 8091 10725 8135 10749
rect 7915 10713 7971 10725
rect 7997 10713 8053 10725
rect 8079 10713 8135 10725
rect 7915 10693 7961 10713
rect 7961 10693 7971 10713
rect 7997 10693 8013 10713
rect 8013 10693 8039 10713
rect 8039 10693 8053 10713
rect 8079 10693 8091 10713
rect 8091 10693 8135 10713
rect 8161 10693 8217 10749
rect 8243 10693 8299 10749
rect 8325 10693 8381 10749
rect 8407 10693 8463 10749
rect 8489 10693 8545 10749
rect 8571 10693 8627 10749
rect 8653 10693 8709 10749
rect 8735 10693 8791 10749
rect 8817 10693 8873 10749
rect 8899 10725 8933 10749
rect 8933 10725 8955 10749
rect 8981 10725 9011 10749
rect 9011 10725 9037 10749
rect 8899 10713 8955 10725
rect 8981 10713 9037 10725
rect 8899 10693 8933 10713
rect 8933 10693 8955 10713
rect 8981 10693 9011 10713
rect 9011 10693 9037 10713
rect 9063 10693 9119 10749
rect 9145 10693 9201 10749
rect 9227 10693 9283 10749
rect 9308 10693 9364 10749
rect 9389 10693 9445 10749
rect 9470 10693 9526 10749
rect 9551 10693 9607 10749
rect 9632 10693 9688 10749
rect 9713 10693 9769 10749
rect 7587 10613 7643 10669
rect 7669 10613 7725 10669
rect 7751 10613 7807 10669
rect 7833 10613 7889 10669
rect 7915 10661 7961 10669
rect 7961 10661 7971 10669
rect 7997 10661 8013 10669
rect 8013 10661 8039 10669
rect 8039 10661 8053 10669
rect 8079 10661 8091 10669
rect 8091 10661 8135 10669
rect 7915 10649 7971 10661
rect 7997 10649 8053 10661
rect 8079 10649 8135 10661
rect 7915 10613 7961 10649
rect 7961 10613 7971 10649
rect 7997 10613 8013 10649
rect 8013 10613 8039 10649
rect 8039 10613 8053 10649
rect 8079 10613 8091 10649
rect 8091 10613 8135 10649
rect 8161 10613 8217 10669
rect 8243 10613 8299 10669
rect 8325 10613 8381 10669
rect 8407 10613 8463 10669
rect 8489 10613 8545 10669
rect 8571 10613 8627 10669
rect 8653 10613 8709 10669
rect 8735 10613 8791 10669
rect 8817 10613 8873 10669
rect 8899 10661 8933 10669
rect 8933 10661 8955 10669
rect 8981 10661 9011 10669
rect 9011 10661 9037 10669
rect 8899 10649 8955 10661
rect 8981 10649 9037 10661
rect 8899 10613 8933 10649
rect 8933 10613 8955 10649
rect 8981 10613 9011 10649
rect 9011 10613 9037 10649
rect 9063 10613 9119 10669
rect 9145 10613 9201 10669
rect 9227 10613 9283 10669
rect 9308 10613 9364 10669
rect 9389 10613 9445 10669
rect 9470 10613 9526 10669
rect 9551 10613 9607 10669
rect 9632 10613 9688 10669
rect 9713 10613 9769 10669
rect 7587 10533 7643 10589
rect 7669 10533 7725 10589
rect 7751 10533 7807 10589
rect 7833 10533 7889 10589
rect 7915 10585 7971 10589
rect 7997 10585 8053 10589
rect 8079 10585 8135 10589
rect 7915 10533 7961 10585
rect 7961 10533 7971 10585
rect 7997 10533 8013 10585
rect 8013 10533 8039 10585
rect 8039 10533 8053 10585
rect 8079 10533 8091 10585
rect 8091 10533 8135 10585
rect 8161 10533 8217 10589
rect 8243 10533 8299 10589
rect 8325 10533 8381 10589
rect 8407 10533 8463 10589
rect 8489 10533 8545 10589
rect 8571 10533 8627 10589
rect 8653 10533 8709 10589
rect 8735 10533 8791 10589
rect 8817 10533 8873 10589
rect 8899 10585 8955 10589
rect 8981 10585 9037 10589
rect 8899 10533 8933 10585
rect 8933 10533 8955 10585
rect 8981 10533 9011 10585
rect 9011 10533 9037 10585
rect 9063 10533 9119 10589
rect 9145 10533 9201 10589
rect 9227 10533 9283 10589
rect 9308 10533 9364 10589
rect 9389 10533 9445 10589
rect 9470 10533 9526 10589
rect 9551 10533 9607 10589
rect 9632 10533 9688 10589
rect 9713 10533 9769 10589
rect 7587 10453 7643 10509
rect 7669 10453 7725 10509
rect 7751 10453 7807 10509
rect 7833 10453 7889 10509
rect 7915 10469 7961 10509
rect 7961 10469 7971 10509
rect 7997 10469 8013 10509
rect 8013 10469 8039 10509
rect 8039 10469 8053 10509
rect 8079 10469 8091 10509
rect 8091 10469 8135 10509
rect 7915 10457 7971 10469
rect 7997 10457 8053 10469
rect 8079 10457 8135 10469
rect 7915 10453 7961 10457
rect 7961 10453 7971 10457
rect 7997 10453 8013 10457
rect 8013 10453 8039 10457
rect 8039 10453 8053 10457
rect 8079 10453 8091 10457
rect 8091 10453 8135 10457
rect 8161 10453 8217 10509
rect 8243 10453 8299 10509
rect 8325 10453 8381 10509
rect 8407 10453 8463 10509
rect 8489 10453 8545 10509
rect 8571 10453 8627 10509
rect 8653 10453 8709 10509
rect 8735 10453 8791 10509
rect 8817 10453 8873 10509
rect 8899 10469 8933 10509
rect 8933 10469 8955 10509
rect 8981 10469 9011 10509
rect 9011 10469 9037 10509
rect 8899 10457 8955 10469
rect 8981 10457 9037 10469
rect 8899 10453 8933 10457
rect 8933 10453 8955 10457
rect 8981 10453 9011 10457
rect 9011 10453 9037 10457
rect 9063 10453 9119 10509
rect 9145 10453 9201 10509
rect 9227 10453 9283 10509
rect 9308 10453 9364 10509
rect 9389 10453 9445 10509
rect 9470 10453 9526 10509
rect 9551 10453 9607 10509
rect 9632 10453 9688 10509
rect 9713 10453 9769 10509
rect 7587 10373 7643 10429
rect 7669 10373 7725 10429
rect 7751 10373 7807 10429
rect 7833 10373 7889 10429
rect 7915 10405 7961 10429
rect 7961 10405 7971 10429
rect 7997 10405 8013 10429
rect 8013 10405 8039 10429
rect 8039 10405 8053 10429
rect 8079 10405 8091 10429
rect 8091 10405 8135 10429
rect 7915 10393 7971 10405
rect 7997 10393 8053 10405
rect 8079 10393 8135 10405
rect 7915 10373 7961 10393
rect 7961 10373 7971 10393
rect 7997 10373 8013 10393
rect 8013 10373 8039 10393
rect 8039 10373 8053 10393
rect 8079 10373 8091 10393
rect 8091 10373 8135 10393
rect 8161 10373 8217 10429
rect 8243 10373 8299 10429
rect 8325 10373 8381 10429
rect 8407 10373 8463 10429
rect 8489 10373 8545 10429
rect 8571 10373 8627 10429
rect 8653 10373 8709 10429
rect 8735 10373 8791 10429
rect 8817 10373 8873 10429
rect 8899 10405 8933 10429
rect 8933 10405 8955 10429
rect 8981 10405 9011 10429
rect 9011 10405 9037 10429
rect 8899 10393 8955 10405
rect 8981 10393 9037 10405
rect 8899 10373 8933 10393
rect 8933 10373 8955 10393
rect 8981 10373 9011 10393
rect 9011 10373 9037 10393
rect 9063 10373 9119 10429
rect 9145 10373 9201 10429
rect 9227 10373 9283 10429
rect 9308 10373 9364 10429
rect 9389 10373 9445 10429
rect 9470 10373 9526 10429
rect 9551 10373 9607 10429
rect 9632 10373 9688 10429
rect 9713 10373 9769 10429
rect 7587 10293 7643 10349
rect 7669 10293 7725 10349
rect 7751 10293 7807 10349
rect 7833 10293 7889 10349
rect 7915 10341 7961 10349
rect 7961 10341 7971 10349
rect 7997 10341 8013 10349
rect 8013 10341 8039 10349
rect 8039 10341 8053 10349
rect 8079 10341 8091 10349
rect 8091 10341 8135 10349
rect 7915 10329 7971 10341
rect 7997 10329 8053 10341
rect 8079 10329 8135 10341
rect 7915 10293 7961 10329
rect 7961 10293 7971 10329
rect 7997 10293 8013 10329
rect 8013 10293 8039 10329
rect 8039 10293 8053 10329
rect 8079 10293 8091 10329
rect 8091 10293 8135 10329
rect 8161 10293 8217 10349
rect 8243 10293 8299 10349
rect 8325 10293 8381 10349
rect 8407 10293 8463 10349
rect 8489 10293 8545 10349
rect 8571 10293 8627 10349
rect 8653 10293 8709 10349
rect 8735 10293 8791 10349
rect 8817 10293 8873 10349
rect 8899 10341 8933 10349
rect 8933 10341 8955 10349
rect 8981 10341 9011 10349
rect 9011 10341 9037 10349
rect 8899 10329 8955 10341
rect 8981 10329 9037 10341
rect 8899 10293 8933 10329
rect 8933 10293 8955 10329
rect 8981 10293 9011 10329
rect 9011 10293 9037 10329
rect 9063 10293 9119 10349
rect 9145 10293 9201 10349
rect 9227 10293 9283 10349
rect 9308 10293 9364 10349
rect 9389 10293 9445 10349
rect 9470 10293 9526 10349
rect 9551 10293 9607 10349
rect 9632 10293 9688 10349
rect 9713 10293 9769 10349
rect 7587 10213 7643 10269
rect 7669 10213 7725 10269
rect 7751 10213 7807 10269
rect 7833 10213 7889 10269
rect 7915 10264 7971 10269
rect 7997 10264 8053 10269
rect 8079 10264 8135 10269
rect 7915 10213 7961 10264
rect 7961 10213 7971 10264
rect 7997 10213 8013 10264
rect 8013 10213 8039 10264
rect 8039 10213 8053 10264
rect 8079 10213 8091 10264
rect 8091 10213 8135 10264
rect 8161 10213 8217 10269
rect 8243 10213 8299 10269
rect 8325 10213 8381 10269
rect 8407 10213 8463 10269
rect 8489 10213 8545 10269
rect 8571 10213 8627 10269
rect 8653 10213 8709 10269
rect 8735 10213 8791 10269
rect 8817 10213 8873 10269
rect 8899 10264 8955 10269
rect 8981 10264 9037 10269
rect 8899 10213 8933 10264
rect 8933 10213 8955 10264
rect 8981 10213 9011 10264
rect 9011 10213 9037 10264
rect 9063 10213 9119 10269
rect 9145 10213 9201 10269
rect 9227 10213 9283 10269
rect 9308 10213 9364 10269
rect 9389 10213 9445 10269
rect 9470 10213 9526 10269
rect 9551 10213 9607 10269
rect 9632 10213 9688 10269
rect 9713 10213 9769 10269
rect 7587 10133 7643 10189
rect 7669 10133 7725 10189
rect 7751 10133 7807 10189
rect 7833 10133 7889 10189
rect 7915 10147 7961 10189
rect 7961 10147 7971 10189
rect 7997 10147 8013 10189
rect 8013 10147 8039 10189
rect 8039 10147 8053 10189
rect 8079 10147 8091 10189
rect 8091 10147 8135 10189
rect 7915 10134 7971 10147
rect 7997 10134 8053 10147
rect 8079 10134 8135 10147
rect 7915 10133 7961 10134
rect 7961 10133 7971 10134
rect 7997 10133 8013 10134
rect 8013 10133 8039 10134
rect 8039 10133 8053 10134
rect 8079 10133 8091 10134
rect 8091 10133 8135 10134
rect 8161 10133 8217 10189
rect 8243 10133 8299 10189
rect 8325 10133 8381 10189
rect 8407 10133 8463 10189
rect 8489 10133 8545 10189
rect 8571 10133 8627 10189
rect 8653 10133 8709 10189
rect 8735 10133 8791 10189
rect 8817 10133 8873 10189
rect 8899 10147 8933 10189
rect 8933 10147 8955 10189
rect 8981 10147 9011 10189
rect 9011 10147 9037 10189
rect 8899 10134 8955 10147
rect 8981 10134 9037 10147
rect 8899 10133 8933 10134
rect 8933 10133 8955 10134
rect 8981 10133 9011 10134
rect 9011 10133 9037 10134
rect 9063 10133 9119 10189
rect 9145 10133 9201 10189
rect 9227 10133 9283 10189
rect 9308 10133 9364 10189
rect 9389 10133 9445 10189
rect 9470 10133 9526 10189
rect 9551 10133 9607 10189
rect 9632 10133 9688 10189
rect 9713 10133 9769 10189
rect 7587 10053 7643 10109
rect 7669 10053 7725 10109
rect 7751 10053 7807 10109
rect 7833 10053 7889 10109
rect 7915 10082 7961 10109
rect 7961 10082 7971 10109
rect 7997 10082 8013 10109
rect 8013 10082 8039 10109
rect 8039 10082 8053 10109
rect 8079 10082 8091 10109
rect 8091 10082 8135 10109
rect 7915 10069 7971 10082
rect 7997 10069 8053 10082
rect 8079 10069 8135 10082
rect 7915 10053 7961 10069
rect 7961 10053 7971 10069
rect 7997 10053 8013 10069
rect 8013 10053 8039 10069
rect 8039 10053 8053 10069
rect 8079 10053 8091 10069
rect 8091 10053 8135 10069
rect 8161 10053 8217 10109
rect 8243 10053 8299 10109
rect 8325 10053 8381 10109
rect 8407 10053 8463 10109
rect 8489 10053 8545 10109
rect 8571 10053 8627 10109
rect 8653 10053 8709 10109
rect 8735 10053 8791 10109
rect 8817 10053 8873 10109
rect 8899 10082 8933 10109
rect 8933 10082 8955 10109
rect 8981 10082 9011 10109
rect 9011 10082 9037 10109
rect 8899 10069 8955 10082
rect 8981 10069 9037 10082
rect 8899 10053 8933 10069
rect 8933 10053 8955 10069
rect 8981 10053 9011 10069
rect 9011 10053 9037 10069
rect 9063 10053 9119 10109
rect 9145 10053 9201 10109
rect 9227 10053 9283 10109
rect 9308 10053 9364 10109
rect 9389 10053 9445 10109
rect 9470 10053 9526 10109
rect 9551 10053 9607 10109
rect 9632 10053 9688 10109
rect 9713 10053 9769 10109
rect 7587 9973 7643 10029
rect 7669 9973 7725 10029
rect 7751 9973 7807 10029
rect 7833 9973 7889 10029
rect 7915 10017 7961 10029
rect 7961 10017 7971 10029
rect 7997 10017 8013 10029
rect 8013 10017 8039 10029
rect 8039 10017 8053 10029
rect 8079 10017 8091 10029
rect 8091 10017 8135 10029
rect 7915 10004 7971 10017
rect 7997 10004 8053 10017
rect 8079 10004 8135 10017
rect 7915 9973 7961 10004
rect 7961 9973 7971 10004
rect 7997 9973 8013 10004
rect 8013 9973 8039 10004
rect 8039 9973 8053 10004
rect 8079 9973 8091 10004
rect 8091 9973 8135 10004
rect 8161 9973 8217 10029
rect 8243 9973 8299 10029
rect 8325 9973 8381 10029
rect 8407 9973 8463 10029
rect 8489 9973 8545 10029
rect 8571 9973 8627 10029
rect 8653 9973 8709 10029
rect 8735 9973 8791 10029
rect 8817 9973 8873 10029
rect 8899 10017 8933 10029
rect 8933 10017 8955 10029
rect 8981 10017 9011 10029
rect 9011 10017 9037 10029
rect 8899 10004 8955 10017
rect 8981 10004 9037 10017
rect 8899 9973 8933 10004
rect 8933 9973 8955 10004
rect 8981 9973 9011 10004
rect 9011 9973 9037 10004
rect 9063 9973 9119 10029
rect 9145 9973 9201 10029
rect 9227 9973 9283 10029
rect 9308 9973 9364 10029
rect 9389 9973 9445 10029
rect 9470 9973 9526 10029
rect 9551 9973 9607 10029
rect 9632 9973 9688 10029
rect 9713 9973 9769 10029
rect 7587 9893 7643 9949
rect 7669 9893 7725 9949
rect 7751 9893 7807 9949
rect 7833 9893 7889 9949
rect 7915 9939 7971 9949
rect 7997 9939 8053 9949
rect 8079 9939 8135 9949
rect 7915 9893 7961 9939
rect 7961 9893 7971 9939
rect 7997 9893 8013 9939
rect 8013 9893 8039 9939
rect 8039 9893 8053 9939
rect 8079 9893 8091 9939
rect 8091 9893 8135 9939
rect 8161 9893 8217 9949
rect 8243 9893 8299 9949
rect 8325 9893 8381 9949
rect 8407 9893 8463 9949
rect 8489 9893 8545 9949
rect 8571 9893 8627 9949
rect 8653 9893 8709 9949
rect 8735 9893 8791 9949
rect 8817 9893 8873 9949
rect 8899 9939 8955 9949
rect 8981 9939 9037 9949
rect 8899 9893 8933 9939
rect 8933 9893 8955 9939
rect 8981 9893 9011 9939
rect 9011 9893 9037 9939
rect 9063 9893 9119 9949
rect 9145 9893 9201 9949
rect 9227 9893 9283 9949
rect 9308 9893 9364 9949
rect 9389 9893 9445 9949
rect 9470 9893 9526 9949
rect 9551 9893 9607 9949
rect 9632 9893 9688 9949
rect 9713 9893 9769 9949
rect 7587 9813 7643 9869
rect 7669 9813 7725 9869
rect 7751 9813 7807 9869
rect 7833 9813 7889 9869
rect 7915 9822 7961 9869
rect 7961 9822 7971 9869
rect 7997 9822 8013 9869
rect 8013 9822 8039 9869
rect 8039 9822 8053 9869
rect 8079 9822 8091 9869
rect 8091 9822 8135 9869
rect 7915 9813 7971 9822
rect 7997 9813 8053 9822
rect 8079 9813 8135 9822
rect 8161 9813 8217 9869
rect 8243 9813 8299 9869
rect 8325 9813 8381 9869
rect 8407 9813 8463 9869
rect 8489 9813 8545 9869
rect 8571 9813 8627 9869
rect 8653 9813 8709 9869
rect 8735 9813 8791 9869
rect 8817 9813 8873 9869
rect 8899 9822 8933 9869
rect 8933 9822 8955 9869
rect 8981 9822 9011 9869
rect 9011 9822 9037 9869
rect 8899 9813 8955 9822
rect 8981 9813 9037 9822
rect 9063 9813 9119 9869
rect 9145 9813 9201 9869
rect 9227 9813 9283 9869
rect 9308 9813 9364 9869
rect 9389 9813 9445 9869
rect 9470 9813 9526 9869
rect 9551 9813 9607 9869
rect 9632 9813 9688 9869
rect 9713 9813 9769 9869
rect 7587 9733 7643 9789
rect 7669 9733 7725 9789
rect 7751 9733 7807 9789
rect 7833 9733 7889 9789
rect 7915 9757 7961 9789
rect 7961 9757 7971 9789
rect 7997 9757 8013 9789
rect 8013 9757 8039 9789
rect 8039 9757 8053 9789
rect 8079 9757 8091 9789
rect 8091 9757 8135 9789
rect 7915 9744 7971 9757
rect 7997 9744 8053 9757
rect 8079 9744 8135 9757
rect 7915 9733 7961 9744
rect 7961 9733 7971 9744
rect 7997 9733 8013 9744
rect 8013 9733 8039 9744
rect 8039 9733 8053 9744
rect 8079 9733 8091 9744
rect 8091 9733 8135 9744
rect 8161 9733 8217 9789
rect 8243 9733 8299 9789
rect 8325 9733 8381 9789
rect 8407 9733 8463 9789
rect 8489 9733 8545 9789
rect 8571 9733 8627 9789
rect 8653 9733 8709 9789
rect 8735 9733 8791 9789
rect 8817 9733 8873 9789
rect 8899 9757 8933 9789
rect 8933 9757 8955 9789
rect 8981 9757 9011 9789
rect 9011 9757 9037 9789
rect 8899 9744 8955 9757
rect 8981 9744 9037 9757
rect 8899 9733 8933 9744
rect 8933 9733 8955 9744
rect 8981 9733 9011 9744
rect 9011 9733 9037 9744
rect 9063 9733 9119 9789
rect 9145 9733 9201 9789
rect 9227 9733 9283 9789
rect 9308 9733 9364 9789
rect 9389 9733 9445 9789
rect 9470 9733 9526 9789
rect 9551 9733 9607 9789
rect 9632 9733 9688 9789
rect 9713 9733 9769 9789
rect 7587 9653 7643 9709
rect 7669 9653 7725 9709
rect 7751 9653 7807 9709
rect 7833 9653 7889 9709
rect 7915 9692 7961 9709
rect 7961 9692 7971 9709
rect 7997 9692 8013 9709
rect 8013 9692 8039 9709
rect 8039 9692 8053 9709
rect 8079 9692 8091 9709
rect 8091 9692 8135 9709
rect 7915 9679 7971 9692
rect 7997 9679 8053 9692
rect 8079 9679 8135 9692
rect 7915 9653 7961 9679
rect 7961 9653 7971 9679
rect 7997 9653 8013 9679
rect 8013 9653 8039 9679
rect 8039 9653 8053 9679
rect 8079 9653 8091 9679
rect 8091 9653 8135 9679
rect 8161 9653 8217 9709
rect 8243 9653 8299 9709
rect 8325 9653 8381 9709
rect 8407 9653 8463 9709
rect 8489 9653 8545 9709
rect 8571 9653 8627 9709
rect 8653 9653 8709 9709
rect 8735 9653 8791 9709
rect 8817 9653 8873 9709
rect 8899 9692 8933 9709
rect 8933 9692 8955 9709
rect 8981 9692 9011 9709
rect 9011 9692 9037 9709
rect 8899 9679 8955 9692
rect 8981 9679 9037 9692
rect 8899 9653 8933 9679
rect 8933 9653 8955 9679
rect 8981 9653 9011 9679
rect 9011 9653 9037 9679
rect 9063 9653 9119 9709
rect 9145 9653 9201 9709
rect 9227 9653 9283 9709
rect 9308 9653 9364 9709
rect 9389 9653 9445 9709
rect 9470 9653 9526 9709
rect 9551 9653 9607 9709
rect 9632 9653 9688 9709
rect 9713 9653 9769 9709
rect 7587 9573 7643 9629
rect 7669 9573 7725 9629
rect 7751 9573 7807 9629
rect 7833 9573 7889 9629
rect 7915 9627 7961 9629
rect 7961 9627 7971 9629
rect 7997 9627 8013 9629
rect 8013 9627 8039 9629
rect 8039 9627 8053 9629
rect 8079 9627 8091 9629
rect 8091 9627 8135 9629
rect 7915 9614 7971 9627
rect 7997 9614 8053 9627
rect 8079 9614 8135 9627
rect 7915 9573 7961 9614
rect 7961 9573 7971 9614
rect 7997 9573 8013 9614
rect 8013 9573 8039 9614
rect 8039 9573 8053 9614
rect 8079 9573 8091 9614
rect 8091 9573 8135 9614
rect 8161 9573 8217 9629
rect 8243 9573 8299 9629
rect 8325 9573 8381 9629
rect 8407 9573 8463 9629
rect 8489 9573 8545 9629
rect 8571 9573 8627 9629
rect 8653 9573 8709 9629
rect 8735 9573 8791 9629
rect 8817 9573 8873 9629
rect 8899 9627 8933 9629
rect 8933 9627 8955 9629
rect 8981 9627 9011 9629
rect 9011 9627 9037 9629
rect 8899 9614 8955 9627
rect 8981 9614 9037 9627
rect 8899 9573 8933 9614
rect 8933 9573 8955 9614
rect 8981 9573 9011 9614
rect 9011 9573 9037 9614
rect 9063 9573 9119 9629
rect 9145 9573 9201 9629
rect 9227 9573 9283 9629
rect 9308 9573 9364 9629
rect 9389 9573 9445 9629
rect 9470 9573 9526 9629
rect 9551 9573 9607 9629
rect 9632 9573 9688 9629
rect 9713 9573 9769 9629
rect 7587 9493 7643 9549
rect 7669 9493 7725 9549
rect 7751 9493 7807 9549
rect 7833 9493 7889 9549
rect 7915 9497 7961 9549
rect 7961 9497 7971 9549
rect 7997 9497 8013 9549
rect 8013 9497 8039 9549
rect 8039 9497 8053 9549
rect 8079 9497 8091 9549
rect 8091 9497 8135 9549
rect 7915 9493 7971 9497
rect 7997 9493 8053 9497
rect 8079 9493 8135 9497
rect 8161 9493 8217 9549
rect 8243 9493 8299 9549
rect 8325 9493 8381 9549
rect 8407 9493 8463 9549
rect 8489 9493 8545 9549
rect 8571 9493 8627 9549
rect 8653 9493 8709 9549
rect 8735 9493 8791 9549
rect 8817 9493 8873 9549
rect 8899 9497 8933 9549
rect 8933 9497 8955 9549
rect 8981 9497 9011 9549
rect 9011 9497 9037 9549
rect 8899 9493 8955 9497
rect 8981 9493 9037 9497
rect 9063 9493 9119 9549
rect 9145 9493 9201 9549
rect 9227 9493 9283 9549
rect 9308 9493 9364 9549
rect 9389 9493 9445 9549
rect 9470 9493 9526 9549
rect 9551 9493 9607 9549
rect 9632 9493 9688 9549
rect 9713 9493 9769 9549
rect 7588 7295 7644 7296
rect 7670 7295 7726 7296
rect 7751 7295 7807 7296
rect 7832 7295 7888 7296
rect 7913 7295 7969 7296
rect 7994 7295 8050 7296
rect 8075 7295 8131 7296
rect 8156 7295 8212 7296
rect 8237 7295 8293 7296
rect 8318 7295 8374 7296
rect 8399 7295 8455 7296
rect 8480 7295 8536 7296
rect 8561 7295 8617 7296
rect 8642 7295 8698 7296
rect 8723 7295 8779 7296
rect 8804 7295 8860 7296
rect 8885 7295 8941 7296
rect 8966 7295 9022 7296
rect 9047 7295 9103 7296
rect 7588 7240 7644 7295
rect 7670 7240 7726 7295
rect 7751 7240 7807 7295
rect 7832 7240 7888 7295
rect 7913 7240 7969 7295
rect 7994 7240 8050 7295
rect 8075 7240 8131 7295
rect 8156 7240 8212 7295
rect 8237 7240 8293 7295
rect 8318 7240 8374 7295
rect 8399 7240 8455 7295
rect 8480 7240 8536 7295
rect 8561 7240 8617 7295
rect 8642 7240 8698 7295
rect 8723 7240 8779 7295
rect 8804 7240 8860 7295
rect 8885 7240 8941 7295
rect 8966 7240 9022 7295
rect 9047 7240 9099 7295
rect 9099 7240 9103 7295
rect 7588 7158 7644 7214
rect 7670 7158 7726 7214
rect 7751 7158 7807 7214
rect 7832 7158 7888 7214
rect 7913 7158 7969 7214
rect 7994 7158 8050 7214
rect 8075 7158 8131 7214
rect 8156 7158 8212 7214
rect 8237 7158 8293 7214
rect 8318 7158 8374 7214
rect 8399 7158 8455 7214
rect 8480 7158 8536 7214
rect 8561 7158 8617 7214
rect 8642 7158 8698 7214
rect 8723 7158 8779 7214
rect 8804 7158 8860 7214
rect 8885 7158 8941 7214
rect 8966 7158 9022 7214
rect 9047 7158 9099 7214
rect 9099 7158 9103 7214
rect 7588 7076 7644 7132
rect 7670 7076 7726 7132
rect 7751 7076 7807 7132
rect 7832 7076 7888 7132
rect 7913 7076 7969 7132
rect 7994 7076 8050 7132
rect 8075 7076 8131 7132
rect 8156 7076 8212 7132
rect 8237 7076 8293 7132
rect 8318 7076 8374 7132
rect 8399 7076 8455 7132
rect 8480 7076 8536 7132
rect 8561 7076 8617 7132
rect 8642 7076 8698 7132
rect 8723 7076 8779 7132
rect 8804 7076 8860 7132
rect 8885 7076 8941 7132
rect 8966 7076 9022 7132
rect 9047 7076 9099 7132
rect 9099 7076 9103 7132
rect 7588 6994 7644 7050
rect 7670 6994 7726 7050
rect 7751 6994 7807 7050
rect 7832 6994 7888 7050
rect 7913 6994 7969 7050
rect 7994 6994 8050 7050
rect 8075 6994 8131 7050
rect 8156 6994 8212 7050
rect 8237 6994 8293 7050
rect 8318 6994 8374 7050
rect 8399 6994 8455 7050
rect 8480 6994 8536 7050
rect 8561 6994 8617 7050
rect 8642 6994 8698 7050
rect 8723 6994 8779 7050
rect 8804 6994 8860 7050
rect 8885 6994 8941 7050
rect 8966 6994 9022 7050
rect 9047 6994 9099 7050
rect 9099 6994 9103 7050
rect 7588 6912 7644 6968
rect 7670 6912 7726 6968
rect 7751 6912 7807 6968
rect 7832 6912 7888 6968
rect 7913 6912 7969 6968
rect 7994 6912 8050 6968
rect 8075 6912 8131 6968
rect 8156 6912 8212 6968
rect 8237 6912 8293 6968
rect 8318 6912 8374 6968
rect 8399 6912 8455 6968
rect 8480 6912 8536 6968
rect 8561 6912 8617 6968
rect 8642 6912 8698 6968
rect 8723 6912 8779 6968
rect 8804 6912 8860 6968
rect 8885 6912 8941 6968
rect 8966 6912 9022 6968
rect 9047 6912 9099 6968
rect 9099 6912 9103 6968
rect 7588 6830 7644 6886
rect 7670 6830 7726 6886
rect 7751 6830 7807 6886
rect 7832 6830 7888 6886
rect 7913 6830 7969 6886
rect 7994 6830 8050 6886
rect 8075 6830 8131 6886
rect 8156 6830 8212 6886
rect 8237 6830 8293 6886
rect 8318 6830 8374 6886
rect 8399 6830 8455 6886
rect 8480 6830 8536 6886
rect 8561 6830 8617 6886
rect 8642 6830 8698 6886
rect 8723 6830 8779 6886
rect 8804 6830 8860 6886
rect 8885 6830 8941 6886
rect 8966 6830 9022 6886
rect 9047 6830 9099 6886
rect 9099 6830 9103 6886
rect 7588 6748 7644 6804
rect 7670 6748 7726 6804
rect 7751 6748 7807 6804
rect 7832 6748 7888 6804
rect 7913 6748 7969 6804
rect 7994 6748 8050 6804
rect 8075 6748 8131 6804
rect 8156 6748 8212 6804
rect 8237 6748 8293 6804
rect 8318 6748 8374 6804
rect 8399 6748 8455 6804
rect 8480 6748 8536 6804
rect 8561 6748 8617 6804
rect 8642 6748 8698 6804
rect 8723 6748 8779 6804
rect 8804 6748 8860 6804
rect 8885 6748 8941 6804
rect 8966 6748 9022 6804
rect 9047 6748 9099 6804
rect 9099 6748 9103 6804
rect 7588 6667 7644 6722
rect 7670 6667 7726 6722
rect 7751 6667 7807 6722
rect 7832 6667 7888 6722
rect 7913 6667 7969 6722
rect 7994 6667 8050 6722
rect 8075 6667 8131 6722
rect 8156 6667 8212 6722
rect 8237 6667 8293 6722
rect 8318 6667 8374 6722
rect 8399 6667 8455 6722
rect 8480 6667 8536 6722
rect 8561 6667 8617 6722
rect 8642 6667 8698 6722
rect 8723 6667 8779 6722
rect 8804 6667 8860 6722
rect 8885 6667 8941 6722
rect 8966 6667 9022 6722
rect 9047 6667 9099 6722
rect 9099 6667 9103 6722
rect 7588 6666 7644 6667
rect 7670 6666 7726 6667
rect 7751 6666 7807 6667
rect 7832 6666 7888 6667
rect 7913 6666 7969 6667
rect 7994 6666 8050 6667
rect 8075 6666 8131 6667
rect 8156 6666 8212 6667
rect 8237 6666 8293 6667
rect 8318 6666 8374 6667
rect 8399 6666 8455 6667
rect 8480 6666 8536 6667
rect 8561 6666 8617 6667
rect 8642 6666 8698 6667
rect 8723 6666 8779 6667
rect 8804 6666 8860 6667
rect 8885 6666 8941 6667
rect 8966 6666 9022 6667
rect 9047 6666 9103 6667
rect 5191 5045 5247 5101
rect 5273 5045 5329 5101
rect 5355 5045 5411 5101
rect 5437 5045 5493 5101
rect 5519 5045 5575 5101
rect 5601 5045 5657 5101
rect 5683 5045 5739 5101
rect 5765 5045 5821 5101
rect 5847 5045 5903 5101
rect 5929 5045 5985 5101
rect 6011 5045 6067 5101
rect 6093 5045 6149 5101
rect 6175 5045 6231 5101
rect 6257 5045 6313 5101
rect 6339 5045 6395 5101
rect 6421 5045 6477 5101
rect 6503 5045 6559 5101
rect 6585 5045 6641 5101
rect 6666 5045 6722 5101
rect 6747 5045 6803 5101
rect 6828 5045 6884 5101
rect 6909 5045 6965 5101
rect 6990 5045 7046 5101
rect 7071 5045 7127 5101
rect 7152 5045 7208 5101
rect 7233 5045 7289 5101
rect 7314 5045 7370 5101
rect 5191 4965 5247 5021
rect 5273 4965 5329 5021
rect 5355 4965 5411 5021
rect 5437 4965 5493 5021
rect 5519 4965 5575 5021
rect 5601 4965 5657 5021
rect 5683 4965 5739 5021
rect 5765 4965 5821 5021
rect 5847 4965 5903 5021
rect 5929 4965 5985 5021
rect 6011 4965 6067 5021
rect 6093 4965 6149 5021
rect 6175 4965 6231 5021
rect 6257 4965 6313 5021
rect 6339 4965 6395 5021
rect 6421 4965 6477 5021
rect 6503 4965 6559 5021
rect 6585 4965 6641 5021
rect 6666 4965 6722 5021
rect 6747 4965 6803 5021
rect 6828 4965 6884 5021
rect 6909 4965 6965 5021
rect 6990 4965 7046 5021
rect 7071 4965 7127 5021
rect 7152 4965 7208 5021
rect 7233 4965 7289 5021
rect 7314 4965 7370 5021
rect 5191 4885 5247 4941
rect 5273 4885 5329 4941
rect 5355 4885 5411 4941
rect 5437 4885 5493 4941
rect 5519 4885 5575 4941
rect 5601 4885 5657 4941
rect 5683 4885 5739 4941
rect 5765 4885 5821 4941
rect 5847 4885 5903 4941
rect 5929 4885 5985 4941
rect 6011 4885 6067 4941
rect 6093 4885 6149 4941
rect 6175 4885 6231 4941
rect 6257 4885 6313 4941
rect 6339 4885 6395 4941
rect 6421 4885 6477 4941
rect 6503 4885 6559 4941
rect 6585 4885 6641 4941
rect 6666 4885 6722 4941
rect 6747 4885 6803 4941
rect 6828 4885 6884 4941
rect 6909 4885 6965 4941
rect 6990 4885 7046 4941
rect 7071 4885 7127 4941
rect 7152 4885 7208 4941
rect 7233 4885 7289 4941
rect 7314 4885 7370 4941
rect 5191 4805 5247 4861
rect 5273 4805 5329 4861
rect 5355 4805 5411 4861
rect 5437 4805 5493 4861
rect 5519 4805 5575 4861
rect 5601 4805 5657 4861
rect 5683 4805 5739 4861
rect 5765 4805 5821 4861
rect 5847 4805 5903 4861
rect 5929 4805 5985 4861
rect 6011 4805 6067 4861
rect 6093 4805 6149 4861
rect 6175 4805 6231 4861
rect 6257 4805 6313 4861
rect 6339 4805 6395 4861
rect 6421 4805 6477 4861
rect 6503 4805 6559 4861
rect 6585 4805 6641 4861
rect 6666 4805 6722 4861
rect 6747 4805 6803 4861
rect 6828 4805 6884 4861
rect 6909 4805 6965 4861
rect 6990 4805 7046 4861
rect 7071 4805 7127 4861
rect 7152 4805 7208 4861
rect 7233 4805 7289 4861
rect 7314 4805 7370 4861
rect 5191 4725 5247 4781
rect 5273 4725 5329 4781
rect 5355 4725 5411 4781
rect 5437 4725 5493 4781
rect 5519 4725 5575 4781
rect 5601 4725 5657 4781
rect 5683 4725 5739 4781
rect 5765 4725 5821 4781
rect 5847 4725 5903 4781
rect 5929 4725 5985 4781
rect 6011 4725 6067 4781
rect 6093 4725 6149 4781
rect 6175 4725 6231 4781
rect 6257 4725 6313 4781
rect 6339 4725 6395 4781
rect 6421 4725 6477 4781
rect 6503 4725 6559 4781
rect 6585 4725 6641 4781
rect 6666 4725 6722 4781
rect 6747 4725 6803 4781
rect 6828 4725 6884 4781
rect 6909 4725 6965 4781
rect 6990 4725 7046 4781
rect 7071 4725 7127 4781
rect 7152 4725 7208 4781
rect 7233 4725 7289 4781
rect 7314 4725 7370 4781
rect 5191 4645 5247 4701
rect 5273 4645 5329 4701
rect 5355 4645 5411 4701
rect 5437 4645 5493 4701
rect 5519 4645 5575 4701
rect 5601 4645 5657 4701
rect 5683 4645 5739 4701
rect 5765 4645 5821 4701
rect 5847 4645 5903 4701
rect 5929 4645 5985 4701
rect 6011 4645 6067 4701
rect 6093 4645 6149 4701
rect 6175 4645 6231 4701
rect 6257 4645 6313 4701
rect 6339 4645 6395 4701
rect 6421 4645 6477 4701
rect 6503 4645 6559 4701
rect 6585 4645 6641 4701
rect 6666 4645 6722 4701
rect 6747 4645 6803 4701
rect 6828 4645 6884 4701
rect 6909 4645 6965 4701
rect 6990 4645 7046 4701
rect 7071 4645 7127 4701
rect 7152 4645 7208 4701
rect 7233 4645 7289 4701
rect 7314 4645 7370 4701
rect 5191 4565 5247 4621
rect 5273 4565 5329 4621
rect 5355 4565 5411 4621
rect 5437 4565 5493 4621
rect 5519 4565 5575 4621
rect 5601 4565 5657 4621
rect 5683 4565 5739 4621
rect 5765 4565 5821 4621
rect 5847 4565 5903 4621
rect 5929 4565 5985 4621
rect 6011 4565 6067 4621
rect 6093 4565 6149 4621
rect 6175 4565 6231 4621
rect 6257 4565 6313 4621
rect 6339 4565 6395 4621
rect 6421 4565 6477 4621
rect 6503 4565 6559 4621
rect 6585 4565 6641 4621
rect 6666 4565 6722 4621
rect 6747 4565 6803 4621
rect 6828 4565 6884 4621
rect 6909 4565 6965 4621
rect 6990 4565 7046 4621
rect 7071 4565 7127 4621
rect 7152 4565 7208 4621
rect 7233 4565 7289 4621
rect 7314 4565 7370 4621
rect 5191 4485 5247 4541
rect 5273 4485 5329 4541
rect 5355 4485 5411 4541
rect 5437 4485 5493 4541
rect 5519 4485 5575 4541
rect 5601 4485 5657 4541
rect 5683 4485 5739 4541
rect 5765 4485 5821 4541
rect 5847 4485 5903 4541
rect 5929 4485 5985 4541
rect 6011 4485 6067 4541
rect 6093 4485 6149 4541
rect 6175 4485 6231 4541
rect 6257 4485 6313 4541
rect 6339 4485 6395 4541
rect 6421 4485 6477 4541
rect 6503 4485 6559 4541
rect 6585 4485 6641 4541
rect 6666 4485 6722 4541
rect 6747 4485 6803 4541
rect 6828 4485 6884 4541
rect 6909 4485 6965 4541
rect 6990 4485 7046 4541
rect 7071 4485 7127 4541
rect 7152 4485 7208 4541
rect 7233 4485 7289 4541
rect 7314 4485 7370 4541
rect 5191 4405 5247 4461
rect 5273 4405 5329 4461
rect 5355 4405 5411 4461
rect 5437 4405 5493 4461
rect 5519 4405 5575 4461
rect 5601 4405 5657 4461
rect 5683 4405 5739 4461
rect 5765 4405 5821 4461
rect 5847 4405 5903 4461
rect 5929 4405 5985 4461
rect 6011 4405 6067 4461
rect 6093 4405 6149 4461
rect 6175 4405 6231 4461
rect 6257 4405 6313 4461
rect 6339 4405 6395 4461
rect 6421 4405 6477 4461
rect 6503 4405 6559 4461
rect 6585 4405 6641 4461
rect 6666 4405 6722 4461
rect 6747 4405 6803 4461
rect 6828 4405 6884 4461
rect 6909 4405 6965 4461
rect 6990 4405 7046 4461
rect 7071 4405 7127 4461
rect 7152 4405 7208 4461
rect 7233 4405 7289 4461
rect 7314 4405 7370 4461
rect 5191 4325 5247 4381
rect 5273 4325 5329 4381
rect 5355 4325 5411 4381
rect 5437 4325 5493 4381
rect 5519 4325 5575 4381
rect 5601 4325 5657 4381
rect 5683 4325 5739 4381
rect 5765 4325 5821 4381
rect 5847 4325 5903 4381
rect 5929 4325 5985 4381
rect 6011 4325 6067 4381
rect 6093 4325 6149 4381
rect 6175 4325 6231 4381
rect 6257 4325 6313 4381
rect 6339 4325 6395 4381
rect 6421 4325 6477 4381
rect 6503 4325 6559 4381
rect 6585 4325 6641 4381
rect 6666 4325 6722 4381
rect 6747 4325 6803 4381
rect 6828 4325 6884 4381
rect 6909 4325 6965 4381
rect 6990 4325 7046 4381
rect 7071 4325 7127 4381
rect 7152 4325 7208 4381
rect 7233 4325 7289 4381
rect 7314 4325 7370 4381
rect 5191 4245 5247 4301
rect 5273 4245 5329 4301
rect 5355 4245 5411 4301
rect 5437 4245 5493 4301
rect 5519 4245 5575 4301
rect 5601 4245 5657 4301
rect 5683 4245 5739 4301
rect 5765 4245 5821 4301
rect 5847 4245 5903 4301
rect 5929 4245 5985 4301
rect 6011 4245 6067 4301
rect 6093 4245 6149 4301
rect 6175 4245 6231 4301
rect 6257 4245 6313 4301
rect 6339 4245 6395 4301
rect 6421 4245 6477 4301
rect 6503 4245 6559 4301
rect 6585 4245 6641 4301
rect 6666 4245 6722 4301
rect 6747 4245 6803 4301
rect 6828 4245 6884 4301
rect 6909 4245 6965 4301
rect 6990 4245 7046 4301
rect 7071 4245 7127 4301
rect 7152 4245 7208 4301
rect 7233 4245 7289 4301
rect 7314 4245 7370 4301
rect 5191 4165 5247 4221
rect 5273 4165 5329 4221
rect 5355 4165 5411 4221
rect 5437 4165 5493 4221
rect 5519 4165 5575 4221
rect 5601 4165 5657 4221
rect 5683 4165 5739 4221
rect 5765 4165 5821 4221
rect 5847 4165 5903 4221
rect 5929 4165 5985 4221
rect 6011 4165 6067 4221
rect 6093 4165 6149 4221
rect 6175 4165 6231 4221
rect 6257 4165 6313 4221
rect 6339 4165 6395 4221
rect 6421 4165 6477 4221
rect 6503 4165 6559 4221
rect 6585 4165 6641 4221
rect 6666 4165 6722 4221
rect 6747 4165 6803 4221
rect 6828 4165 6884 4221
rect 6909 4165 6965 4221
rect 6990 4165 7046 4221
rect 7071 4165 7127 4221
rect 7152 4165 7208 4221
rect 7233 4165 7289 4221
rect 7314 4165 7370 4221
rect 5191 4085 5247 4141
rect 5273 4085 5329 4141
rect 5355 4085 5411 4141
rect 5437 4085 5493 4141
rect 5519 4085 5575 4141
rect 5601 4085 5657 4141
rect 5683 4085 5739 4141
rect 5765 4085 5821 4141
rect 5847 4085 5903 4141
rect 5929 4085 5985 4141
rect 6011 4085 6067 4141
rect 6093 4085 6149 4141
rect 6175 4085 6231 4141
rect 6257 4085 6313 4141
rect 6339 4085 6395 4141
rect 6421 4085 6477 4141
rect 6503 4085 6559 4141
rect 6585 4085 6641 4141
rect 6666 4085 6722 4141
rect 6747 4085 6803 4141
rect 6828 4085 6884 4141
rect 6909 4085 6965 4141
rect 6990 4085 7046 4141
rect 7071 4085 7127 4141
rect 7152 4085 7208 4141
rect 7233 4085 7289 4141
rect 7314 4085 7370 4141
rect 5191 4005 5247 4061
rect 5273 4005 5329 4061
rect 5355 4005 5411 4061
rect 5437 4005 5493 4061
rect 5519 4005 5575 4061
rect 5601 4005 5657 4061
rect 5683 4005 5739 4061
rect 5765 4005 5821 4061
rect 5847 4005 5903 4061
rect 5929 4005 5985 4061
rect 6011 4005 6067 4061
rect 6093 4005 6149 4061
rect 6175 4005 6231 4061
rect 6257 4005 6313 4061
rect 6339 4005 6395 4061
rect 6421 4005 6477 4061
rect 6503 4005 6559 4061
rect 6585 4005 6641 4061
rect 6666 4005 6722 4061
rect 6747 4005 6803 4061
rect 6828 4005 6884 4061
rect 6909 4005 6965 4061
rect 6990 4005 7046 4061
rect 7071 4005 7127 4061
rect 7152 4005 7208 4061
rect 7233 4005 7289 4061
rect 7314 4005 7370 4061
rect 5191 3925 5247 3981
rect 5273 3925 5329 3981
rect 5355 3925 5411 3981
rect 5437 3925 5493 3981
rect 5519 3925 5575 3981
rect 5601 3925 5657 3981
rect 5683 3925 5739 3981
rect 5765 3925 5821 3981
rect 5847 3925 5903 3981
rect 5929 3925 5985 3981
rect 6011 3925 6067 3981
rect 6093 3925 6149 3981
rect 6175 3925 6231 3981
rect 6257 3925 6313 3981
rect 6339 3925 6395 3981
rect 6421 3925 6477 3981
rect 6503 3925 6559 3981
rect 6585 3925 6641 3981
rect 6666 3925 6722 3981
rect 6747 3925 6803 3981
rect 6828 3925 6884 3981
rect 6909 3925 6965 3981
rect 6990 3925 7046 3981
rect 7071 3925 7127 3981
rect 7152 3925 7208 3981
rect 7233 3925 7289 3981
rect 7314 3925 7370 3981
rect 5191 3845 5247 3901
rect 5273 3845 5329 3901
rect 5355 3845 5411 3901
rect 5437 3845 5493 3901
rect 5519 3845 5575 3901
rect 5601 3845 5657 3901
rect 5683 3845 5739 3901
rect 5765 3845 5821 3901
rect 5847 3845 5903 3901
rect 5929 3845 5985 3901
rect 6011 3845 6067 3901
rect 6093 3845 6149 3901
rect 6175 3845 6231 3901
rect 6257 3845 6313 3901
rect 6339 3845 6395 3901
rect 6421 3845 6477 3901
rect 6503 3845 6559 3901
rect 6585 3845 6641 3901
rect 6666 3845 6722 3901
rect 6747 3845 6803 3901
rect 6828 3845 6884 3901
rect 6909 3845 6965 3901
rect 6990 3845 7046 3901
rect 7071 3845 7127 3901
rect 7152 3845 7208 3901
rect 7233 3845 7289 3901
rect 7314 3845 7370 3901
rect 5191 3765 5247 3821
rect 5273 3765 5329 3821
rect 5355 3765 5411 3821
rect 5437 3765 5493 3821
rect 5519 3765 5575 3821
rect 5601 3765 5657 3821
rect 5683 3765 5739 3821
rect 5765 3765 5821 3821
rect 5847 3765 5903 3821
rect 5929 3765 5985 3821
rect 6011 3765 6067 3821
rect 6093 3765 6149 3821
rect 6175 3765 6231 3821
rect 6257 3765 6313 3821
rect 6339 3765 6395 3821
rect 6421 3765 6477 3821
rect 6503 3765 6559 3821
rect 6585 3765 6641 3821
rect 6666 3765 6722 3821
rect 6747 3765 6803 3821
rect 6828 3765 6884 3821
rect 6909 3765 6965 3821
rect 6990 3765 7046 3821
rect 7071 3765 7127 3821
rect 7152 3765 7208 3821
rect 7233 3765 7289 3821
rect 7314 3765 7370 3821
rect 5191 3685 5247 3741
rect 5273 3685 5329 3741
rect 5355 3685 5411 3741
rect 5437 3685 5493 3741
rect 5519 3685 5575 3741
rect 5601 3685 5657 3741
rect 5683 3685 5739 3741
rect 5765 3685 5821 3741
rect 5847 3685 5903 3741
rect 5929 3685 5985 3741
rect 6011 3685 6067 3741
rect 6093 3685 6149 3741
rect 6175 3685 6231 3741
rect 6257 3685 6313 3741
rect 6339 3685 6395 3741
rect 6421 3685 6477 3741
rect 6503 3685 6559 3741
rect 6585 3685 6641 3741
rect 6666 3685 6722 3741
rect 6747 3685 6803 3741
rect 6828 3685 6884 3741
rect 6909 3685 6965 3741
rect 6990 3685 7046 3741
rect 7071 3685 7127 3741
rect 7152 3685 7208 3741
rect 7233 3685 7289 3741
rect 7314 3685 7370 3741
rect 5191 3605 5247 3661
rect 5273 3605 5329 3661
rect 5355 3605 5411 3661
rect 5437 3605 5493 3661
rect 5519 3605 5575 3661
rect 5601 3605 5657 3661
rect 5683 3605 5739 3661
rect 5765 3605 5821 3661
rect 5847 3605 5903 3661
rect 5929 3605 5985 3661
rect 6011 3605 6067 3661
rect 6093 3605 6149 3661
rect 6175 3605 6231 3661
rect 6257 3605 6313 3661
rect 6339 3605 6395 3661
rect 6421 3605 6477 3661
rect 6503 3605 6559 3661
rect 6585 3605 6641 3661
rect 6666 3605 6722 3661
rect 6747 3605 6803 3661
rect 6828 3605 6884 3661
rect 6909 3605 6965 3661
rect 6990 3605 7046 3661
rect 7071 3605 7127 3661
rect 7152 3605 7208 3661
rect 7233 3605 7289 3661
rect 7314 3605 7370 3661
rect 5191 3525 5247 3581
rect 5273 3525 5329 3581
rect 5355 3525 5411 3581
rect 5437 3525 5493 3581
rect 5519 3525 5575 3581
rect 5601 3525 5657 3581
rect 5683 3525 5739 3581
rect 5765 3525 5821 3581
rect 5847 3525 5903 3581
rect 5929 3525 5985 3581
rect 6011 3525 6067 3581
rect 6093 3525 6149 3581
rect 6175 3525 6231 3581
rect 6257 3525 6313 3581
rect 6339 3525 6395 3581
rect 6421 3525 6477 3581
rect 6503 3525 6559 3581
rect 6585 3525 6641 3581
rect 6666 3525 6722 3581
rect 6747 3525 6803 3581
rect 6828 3525 6884 3581
rect 6909 3525 6965 3581
rect 6990 3525 7046 3581
rect 7071 3525 7127 3581
rect 7152 3525 7208 3581
rect 7233 3525 7289 3581
rect 7314 3525 7370 3581
rect 5191 3445 5247 3501
rect 5273 3445 5329 3501
rect 5355 3445 5411 3501
rect 5437 3445 5493 3501
rect 5519 3445 5575 3501
rect 5601 3445 5657 3501
rect 5683 3445 5739 3501
rect 5765 3445 5821 3501
rect 5847 3445 5903 3501
rect 5929 3445 5985 3501
rect 6011 3445 6067 3501
rect 6093 3445 6149 3501
rect 6175 3445 6231 3501
rect 6257 3445 6313 3501
rect 6339 3445 6395 3501
rect 6421 3445 6477 3501
rect 6503 3445 6559 3501
rect 6585 3445 6641 3501
rect 6666 3445 6722 3501
rect 6747 3445 6803 3501
rect 6828 3445 6884 3501
rect 6909 3445 6965 3501
rect 6990 3445 7046 3501
rect 7071 3445 7127 3501
rect 7152 3445 7208 3501
rect 7233 3445 7289 3501
rect 7314 3445 7370 3501
rect 5191 3365 5247 3421
rect 5273 3365 5329 3421
rect 5355 3365 5411 3421
rect 5437 3365 5493 3421
rect 5519 3365 5575 3421
rect 5601 3365 5657 3421
rect 5683 3365 5739 3421
rect 5765 3365 5821 3421
rect 5847 3365 5903 3421
rect 5929 3365 5985 3421
rect 6011 3365 6067 3421
rect 6093 3365 6149 3421
rect 6175 3365 6231 3421
rect 6257 3365 6313 3421
rect 6339 3365 6395 3421
rect 6421 3365 6477 3421
rect 6503 3365 6559 3421
rect 6585 3365 6641 3421
rect 6666 3365 6722 3421
rect 6747 3365 6803 3421
rect 6828 3365 6884 3421
rect 6909 3365 6965 3421
rect 6990 3365 7046 3421
rect 7071 3365 7127 3421
rect 7152 3365 7208 3421
rect 7233 3365 7289 3421
rect 7314 3365 7370 3421
rect 5191 3285 5247 3341
rect 5273 3285 5329 3341
rect 5355 3285 5411 3341
rect 5437 3285 5493 3341
rect 5519 3285 5575 3341
rect 5601 3285 5657 3341
rect 5683 3285 5739 3341
rect 5765 3285 5821 3341
rect 5847 3285 5903 3341
rect 5929 3285 5985 3341
rect 6011 3285 6067 3341
rect 6093 3285 6149 3341
rect 6175 3285 6231 3341
rect 6257 3285 6313 3341
rect 6339 3285 6395 3341
rect 6421 3285 6477 3341
rect 6503 3285 6559 3341
rect 6585 3285 6641 3341
rect 6666 3285 6722 3341
rect 6747 3285 6803 3341
rect 6828 3285 6884 3341
rect 6909 3285 6965 3341
rect 6990 3285 7046 3341
rect 7071 3285 7127 3341
rect 7152 3285 7208 3341
rect 7233 3285 7289 3341
rect 7314 3285 7370 3341
rect 5191 3205 5247 3261
rect 5273 3205 5329 3261
rect 5355 3205 5411 3261
rect 5437 3205 5493 3261
rect 5519 3205 5575 3261
rect 5601 3205 5657 3261
rect 5683 3205 5739 3261
rect 5765 3205 5821 3261
rect 5847 3205 5903 3261
rect 5929 3205 5985 3261
rect 6011 3205 6067 3261
rect 6093 3205 6149 3261
rect 6175 3205 6231 3261
rect 6257 3205 6313 3261
rect 6339 3205 6395 3261
rect 6421 3205 6477 3261
rect 6503 3205 6559 3261
rect 6585 3205 6641 3261
rect 6666 3205 6722 3261
rect 6747 3205 6803 3261
rect 6828 3205 6884 3261
rect 6909 3205 6965 3261
rect 6990 3205 7046 3261
rect 7071 3205 7127 3261
rect 7152 3205 7208 3261
rect 7233 3205 7289 3261
rect 7314 3205 7370 3261
rect 5191 3125 5247 3181
rect 5273 3125 5329 3181
rect 5355 3125 5411 3181
rect 5437 3125 5493 3181
rect 5519 3125 5575 3181
rect 5601 3125 5657 3181
rect 5683 3125 5739 3181
rect 5765 3125 5821 3181
rect 5847 3125 5903 3181
rect 5929 3125 5985 3181
rect 6011 3125 6067 3181
rect 6093 3125 6149 3181
rect 6175 3125 6231 3181
rect 6257 3125 6313 3181
rect 6339 3125 6395 3181
rect 6421 3125 6477 3181
rect 6503 3125 6559 3181
rect 6585 3125 6641 3181
rect 6666 3125 6722 3181
rect 6747 3125 6803 3181
rect 6828 3125 6884 3181
rect 6909 3125 6965 3181
rect 6990 3125 7046 3181
rect 7071 3125 7127 3181
rect 7152 3125 7208 3181
rect 7233 3125 7289 3181
rect 7314 3125 7370 3181
rect 5191 3045 5247 3101
rect 5273 3045 5329 3101
rect 5355 3045 5411 3101
rect 5437 3045 5493 3101
rect 5519 3045 5575 3101
rect 5601 3045 5657 3101
rect 5683 3045 5739 3101
rect 5765 3045 5821 3101
rect 5847 3045 5903 3101
rect 5929 3045 5985 3101
rect 6011 3045 6067 3101
rect 6093 3045 6149 3101
rect 6175 3045 6231 3101
rect 6257 3045 6313 3101
rect 6339 3045 6395 3101
rect 6421 3045 6477 3101
rect 6503 3045 6559 3101
rect 6585 3045 6641 3101
rect 6666 3045 6722 3101
rect 6747 3045 6803 3101
rect 6828 3045 6884 3101
rect 6909 3045 6965 3101
rect 6990 3045 7046 3101
rect 7071 3045 7127 3101
rect 7152 3045 7208 3101
rect 7233 3045 7289 3101
rect 7314 3045 7370 3101
rect 5191 2965 5247 3021
rect 5273 2965 5329 3021
rect 5355 2965 5411 3021
rect 5437 2965 5493 3021
rect 5519 2965 5575 3021
rect 5601 2965 5657 3021
rect 5683 2965 5739 3021
rect 5765 2965 5821 3021
rect 5847 2965 5903 3021
rect 5929 2965 5985 3021
rect 6011 2965 6067 3021
rect 6093 2965 6149 3021
rect 6175 2965 6231 3021
rect 6257 2965 6313 3021
rect 6339 2965 6395 3021
rect 6421 2965 6477 3021
rect 6503 2965 6559 3021
rect 6585 2965 6641 3021
rect 6666 2965 6722 3021
rect 6747 2965 6803 3021
rect 6828 2965 6884 3021
rect 6909 2965 6965 3021
rect 6990 2965 7046 3021
rect 7071 2965 7127 3021
rect 7152 2965 7208 3021
rect 7233 2965 7289 3021
rect 7314 2965 7370 3021
rect 5191 2885 5247 2941
rect 5273 2885 5329 2941
rect 5355 2885 5411 2941
rect 5437 2885 5493 2941
rect 5519 2885 5575 2941
rect 5601 2885 5657 2941
rect 5683 2885 5739 2941
rect 5765 2885 5821 2941
rect 5847 2885 5903 2941
rect 5929 2885 5985 2941
rect 6011 2885 6067 2941
rect 6093 2885 6149 2941
rect 6175 2885 6231 2941
rect 6257 2885 6313 2941
rect 6339 2885 6395 2941
rect 6421 2885 6477 2941
rect 6503 2885 6559 2941
rect 6585 2885 6641 2941
rect 6666 2885 6722 2941
rect 6747 2885 6803 2941
rect 6828 2885 6884 2941
rect 6909 2885 6965 2941
rect 6990 2885 7046 2941
rect 7071 2885 7127 2941
rect 7152 2885 7208 2941
rect 7233 2885 7289 2941
rect 7314 2885 7370 2941
rect 5191 2805 5247 2861
rect 5273 2805 5329 2861
rect 5355 2805 5411 2861
rect 5437 2805 5493 2861
rect 5519 2805 5575 2861
rect 5601 2805 5657 2861
rect 5683 2805 5739 2861
rect 5765 2805 5821 2861
rect 5847 2805 5903 2861
rect 5929 2805 5985 2861
rect 6011 2805 6067 2861
rect 6093 2805 6149 2861
rect 6175 2805 6231 2861
rect 6257 2805 6313 2861
rect 6339 2805 6395 2861
rect 6421 2805 6477 2861
rect 6503 2805 6559 2861
rect 6585 2805 6641 2861
rect 6666 2805 6722 2861
rect 6747 2805 6803 2861
rect 6828 2805 6884 2861
rect 6909 2805 6965 2861
rect 6990 2805 7046 2861
rect 7071 2805 7127 2861
rect 7152 2805 7208 2861
rect 7233 2805 7289 2861
rect 7314 2805 7370 2861
rect 5191 2725 5247 2781
rect 5273 2725 5329 2781
rect 5355 2725 5411 2781
rect 5437 2725 5493 2781
rect 5519 2725 5575 2781
rect 5601 2725 5657 2781
rect 5683 2725 5739 2781
rect 5765 2725 5821 2781
rect 5847 2725 5903 2781
rect 5929 2725 5985 2781
rect 6011 2725 6067 2781
rect 6093 2725 6149 2781
rect 6175 2725 6231 2781
rect 6257 2725 6313 2781
rect 6339 2725 6395 2781
rect 6421 2725 6477 2781
rect 6503 2725 6559 2781
rect 6585 2725 6641 2781
rect 6666 2725 6722 2781
rect 6747 2725 6803 2781
rect 6828 2725 6884 2781
rect 6909 2725 6965 2781
rect 6990 2725 7046 2781
rect 7071 2725 7127 2781
rect 7152 2725 7208 2781
rect 7233 2725 7289 2781
rect 7314 2725 7370 2781
rect 5191 2645 5247 2701
rect 5273 2645 5329 2701
rect 5355 2645 5411 2701
rect 5437 2645 5493 2701
rect 5519 2645 5575 2701
rect 5601 2645 5657 2701
rect 5683 2645 5739 2701
rect 5765 2645 5821 2701
rect 5847 2645 5903 2701
rect 5929 2645 5985 2701
rect 6011 2645 6067 2701
rect 6093 2645 6149 2701
rect 6175 2645 6231 2701
rect 6257 2645 6313 2701
rect 6339 2645 6395 2701
rect 6421 2645 6477 2701
rect 6503 2645 6559 2701
rect 6585 2645 6641 2701
rect 6666 2645 6722 2701
rect 6747 2645 6803 2701
rect 6828 2645 6884 2701
rect 6909 2645 6965 2701
rect 6990 2645 7046 2701
rect 7071 2645 7127 2701
rect 7152 2645 7208 2701
rect 7233 2645 7289 2701
rect 7314 2645 7370 2701
rect 5191 2565 5247 2621
rect 5273 2565 5329 2621
rect 5355 2565 5411 2621
rect 5437 2565 5493 2621
rect 5519 2565 5575 2621
rect 5601 2565 5657 2621
rect 5683 2565 5739 2621
rect 5765 2565 5821 2621
rect 5847 2565 5903 2621
rect 5929 2565 5985 2621
rect 6011 2565 6067 2621
rect 6093 2565 6149 2621
rect 6175 2565 6231 2621
rect 6257 2565 6313 2621
rect 6339 2565 6395 2621
rect 6421 2565 6477 2621
rect 6503 2565 6559 2621
rect 6585 2565 6641 2621
rect 6666 2565 6722 2621
rect 6747 2565 6803 2621
rect 6828 2565 6884 2621
rect 6909 2565 6965 2621
rect 6990 2565 7046 2621
rect 7071 2565 7127 2621
rect 7152 2565 7208 2621
rect 7233 2565 7289 2621
rect 7314 2565 7370 2621
rect 5191 2485 5247 2541
rect 5273 2485 5329 2541
rect 5355 2485 5411 2541
rect 5437 2485 5493 2541
rect 5519 2485 5575 2541
rect 5601 2485 5657 2541
rect 5683 2485 5739 2541
rect 5765 2485 5821 2541
rect 5847 2485 5903 2541
rect 5929 2485 5985 2541
rect 6011 2485 6067 2541
rect 6093 2485 6149 2541
rect 6175 2485 6231 2541
rect 6257 2485 6313 2541
rect 6339 2485 6395 2541
rect 6421 2485 6477 2541
rect 6503 2485 6559 2541
rect 6585 2485 6641 2541
rect 6666 2485 6722 2541
rect 6747 2485 6803 2541
rect 6828 2485 6884 2541
rect 6909 2485 6965 2541
rect 6990 2485 7046 2541
rect 7071 2485 7127 2541
rect 7152 2485 7208 2541
rect 7233 2485 7289 2541
rect 7314 2485 7370 2541
rect 7587 5036 7643 5092
rect 7669 5036 7725 5092
rect 7751 5036 7807 5092
rect 7833 5036 7889 5092
rect 7915 5036 7971 5092
rect 7997 5036 8053 5092
rect 8079 5036 8135 5092
rect 8161 5036 8217 5092
rect 8243 5036 8299 5092
rect 8325 5036 8381 5092
rect 8407 5036 8463 5092
rect 8489 5036 8545 5092
rect 8571 5036 8627 5092
rect 8653 5036 8709 5092
rect 8735 5036 8791 5092
rect 8817 5036 8873 5092
rect 8899 5036 8955 5092
rect 8981 5036 9037 5092
rect 9063 5036 9119 5092
rect 9145 5036 9201 5092
rect 9227 5036 9283 5092
rect 9308 5036 9364 5092
rect 9389 5036 9445 5092
rect 9470 5036 9526 5092
rect 9551 5036 9607 5092
rect 9632 5036 9688 5092
rect 9713 5036 9769 5092
rect 7587 4956 7643 5012
rect 7669 4956 7725 5012
rect 7751 4956 7807 5012
rect 7833 4956 7889 5012
rect 7915 4956 7971 5012
rect 7997 4956 8053 5012
rect 8079 4956 8135 5012
rect 8161 4956 8217 5012
rect 8243 4956 8299 5012
rect 8325 4956 8381 5012
rect 8407 4956 8463 5012
rect 8489 4956 8545 5012
rect 8571 4956 8627 5012
rect 8653 4956 8709 5012
rect 8735 4956 8791 5012
rect 8817 4956 8873 5012
rect 8899 4956 8955 5012
rect 8981 4956 9037 5012
rect 9063 4956 9119 5012
rect 9145 4956 9201 5012
rect 9227 4956 9283 5012
rect 9308 4956 9364 5012
rect 9389 4956 9445 5012
rect 9470 4956 9526 5012
rect 9551 4956 9607 5012
rect 9632 4956 9688 5012
rect 9713 4956 9769 5012
rect 7587 4876 7643 4932
rect 7669 4876 7725 4932
rect 7751 4876 7807 4932
rect 7833 4876 7889 4932
rect 7915 4876 7971 4932
rect 7997 4876 8053 4932
rect 8079 4876 8135 4932
rect 8161 4876 8217 4932
rect 8243 4876 8299 4932
rect 8325 4876 8381 4932
rect 8407 4876 8463 4932
rect 8489 4876 8545 4932
rect 8571 4876 8627 4932
rect 8653 4876 8709 4932
rect 8735 4876 8791 4932
rect 8817 4876 8873 4932
rect 8899 4876 8955 4932
rect 8981 4876 9037 4932
rect 9063 4876 9119 4932
rect 9145 4876 9201 4932
rect 9227 4876 9283 4932
rect 9308 4876 9364 4932
rect 9389 4876 9445 4932
rect 9470 4876 9526 4932
rect 9551 4876 9607 4932
rect 9632 4876 9688 4932
rect 9713 4876 9769 4932
rect 7587 4796 7643 4852
rect 7669 4796 7725 4852
rect 7751 4796 7807 4852
rect 7833 4796 7889 4852
rect 7915 4796 7971 4852
rect 7997 4796 8053 4852
rect 8079 4796 8135 4852
rect 8161 4796 8217 4852
rect 8243 4796 8299 4852
rect 8325 4796 8381 4852
rect 8407 4796 8463 4852
rect 8489 4796 8545 4852
rect 8571 4796 8627 4852
rect 8653 4796 8709 4852
rect 8735 4796 8791 4852
rect 8817 4796 8873 4852
rect 8899 4796 8955 4852
rect 8981 4796 9037 4852
rect 9063 4796 9119 4852
rect 9145 4796 9201 4852
rect 9227 4796 9283 4852
rect 9308 4796 9364 4852
rect 9389 4796 9445 4852
rect 9470 4796 9526 4852
rect 9551 4796 9607 4852
rect 9632 4796 9688 4852
rect 9713 4796 9769 4852
rect 7587 4716 7643 4772
rect 7669 4716 7725 4772
rect 7751 4716 7807 4772
rect 7833 4716 7889 4772
rect 7915 4716 7971 4772
rect 7997 4716 8053 4772
rect 8079 4716 8135 4772
rect 8161 4716 8217 4772
rect 8243 4716 8299 4772
rect 8325 4716 8381 4772
rect 8407 4716 8463 4772
rect 8489 4716 8545 4772
rect 8571 4716 8627 4772
rect 8653 4716 8709 4772
rect 8735 4716 8791 4772
rect 8817 4716 8873 4772
rect 8899 4716 8955 4772
rect 8981 4716 9037 4772
rect 9063 4716 9119 4772
rect 9145 4716 9201 4772
rect 9227 4716 9283 4772
rect 9308 4716 9364 4772
rect 9389 4716 9445 4772
rect 9470 4716 9526 4772
rect 9551 4716 9607 4772
rect 9632 4716 9688 4772
rect 9713 4716 9769 4772
rect 7587 4636 7643 4692
rect 7669 4636 7725 4692
rect 7751 4636 7807 4692
rect 7833 4636 7889 4692
rect 7915 4636 7971 4692
rect 7997 4636 8053 4692
rect 8079 4636 8135 4692
rect 8161 4636 8217 4692
rect 8243 4636 8299 4692
rect 8325 4636 8381 4692
rect 8407 4636 8463 4692
rect 8489 4636 8545 4692
rect 8571 4636 8627 4692
rect 8653 4636 8709 4692
rect 8735 4636 8791 4692
rect 8817 4636 8873 4692
rect 8899 4636 8955 4692
rect 8981 4636 9037 4692
rect 9063 4636 9119 4692
rect 9145 4636 9201 4692
rect 9227 4636 9283 4692
rect 9308 4636 9364 4692
rect 9389 4636 9445 4692
rect 9470 4636 9526 4692
rect 9551 4636 9607 4692
rect 9632 4636 9688 4692
rect 9713 4636 9769 4692
rect 7587 4556 7643 4612
rect 7669 4556 7725 4612
rect 7751 4556 7807 4612
rect 7833 4556 7889 4612
rect 7915 4556 7971 4612
rect 7997 4556 8053 4612
rect 8079 4556 8135 4612
rect 8161 4556 8217 4612
rect 8243 4556 8299 4612
rect 8325 4556 8381 4612
rect 8407 4556 8463 4612
rect 8489 4556 8545 4612
rect 8571 4556 8627 4612
rect 8653 4556 8709 4612
rect 8735 4556 8791 4612
rect 8817 4556 8873 4612
rect 8899 4556 8955 4612
rect 8981 4556 9037 4612
rect 9063 4556 9119 4612
rect 9145 4556 9201 4612
rect 9227 4556 9283 4612
rect 9308 4556 9364 4612
rect 9389 4556 9445 4612
rect 9470 4556 9526 4612
rect 9551 4556 9607 4612
rect 9632 4556 9688 4612
rect 9713 4556 9769 4612
rect 7587 4476 7643 4532
rect 7669 4476 7725 4532
rect 7751 4476 7807 4532
rect 7833 4476 7889 4532
rect 7915 4476 7971 4532
rect 7997 4476 8053 4532
rect 8079 4476 8135 4532
rect 8161 4476 8217 4532
rect 8243 4476 8299 4532
rect 8325 4476 8381 4532
rect 8407 4476 8463 4532
rect 8489 4476 8545 4532
rect 8571 4476 8627 4532
rect 8653 4476 8709 4532
rect 8735 4476 8791 4532
rect 8817 4476 8873 4532
rect 8899 4476 8955 4532
rect 8981 4476 9037 4532
rect 9063 4476 9119 4532
rect 9145 4476 9201 4532
rect 9227 4476 9283 4532
rect 9308 4476 9364 4532
rect 9389 4476 9445 4532
rect 9470 4476 9526 4532
rect 9551 4476 9607 4532
rect 9632 4476 9688 4532
rect 9713 4476 9769 4532
rect 7587 4396 7643 4452
rect 7669 4396 7725 4452
rect 7751 4396 7807 4452
rect 7833 4396 7889 4452
rect 7915 4396 7971 4452
rect 7997 4396 8053 4452
rect 8079 4396 8135 4452
rect 8161 4396 8217 4452
rect 8243 4396 8299 4452
rect 8325 4396 8381 4452
rect 8407 4396 8463 4452
rect 8489 4396 8545 4452
rect 8571 4396 8627 4452
rect 8653 4396 8709 4452
rect 8735 4396 8791 4452
rect 8817 4396 8873 4452
rect 8899 4396 8955 4452
rect 8981 4396 9037 4452
rect 9063 4396 9119 4452
rect 9145 4396 9201 4452
rect 9227 4396 9283 4452
rect 9308 4396 9364 4452
rect 9389 4396 9445 4452
rect 9470 4396 9526 4452
rect 9551 4396 9607 4452
rect 9632 4396 9688 4452
rect 9713 4396 9769 4452
rect 7587 4316 7643 4372
rect 7669 4316 7725 4372
rect 7751 4316 7807 4372
rect 7833 4316 7889 4372
rect 7915 4316 7971 4372
rect 7997 4316 8053 4372
rect 8079 4316 8135 4372
rect 8161 4316 8217 4372
rect 8243 4316 8299 4372
rect 8325 4316 8381 4372
rect 8407 4316 8463 4372
rect 8489 4316 8545 4372
rect 8571 4316 8627 4372
rect 8653 4316 8709 4372
rect 8735 4316 8791 4372
rect 8817 4316 8873 4372
rect 8899 4316 8955 4372
rect 8981 4316 9037 4372
rect 9063 4316 9119 4372
rect 9145 4316 9201 4372
rect 9227 4316 9283 4372
rect 9308 4316 9364 4372
rect 9389 4316 9445 4372
rect 9470 4316 9526 4372
rect 9551 4316 9607 4372
rect 9632 4316 9688 4372
rect 9713 4316 9769 4372
rect 7587 4236 7643 4292
rect 7669 4236 7725 4292
rect 7751 4236 7807 4292
rect 7833 4236 7889 4292
rect 7915 4236 7971 4292
rect 7997 4236 8053 4292
rect 8079 4236 8135 4292
rect 8161 4236 8217 4292
rect 8243 4236 8299 4292
rect 8325 4236 8381 4292
rect 8407 4236 8463 4292
rect 8489 4236 8545 4292
rect 8571 4236 8627 4292
rect 8653 4236 8709 4292
rect 8735 4236 8791 4292
rect 8817 4236 8873 4292
rect 8899 4236 8955 4292
rect 8981 4236 9037 4292
rect 9063 4236 9119 4292
rect 9145 4236 9201 4292
rect 9227 4236 9283 4292
rect 9308 4236 9364 4292
rect 9389 4236 9445 4292
rect 9470 4236 9526 4292
rect 9551 4236 9607 4292
rect 9632 4236 9688 4292
rect 9713 4236 9769 4292
rect 7587 4156 7643 4212
rect 7669 4156 7725 4212
rect 7751 4156 7807 4212
rect 7833 4156 7889 4212
rect 7915 4156 7971 4212
rect 7997 4156 8053 4212
rect 8079 4156 8135 4212
rect 8161 4156 8217 4212
rect 8243 4156 8299 4212
rect 8325 4156 8381 4212
rect 8407 4156 8463 4212
rect 8489 4156 8545 4212
rect 8571 4156 8627 4212
rect 8653 4156 8709 4212
rect 8735 4156 8791 4212
rect 8817 4156 8873 4212
rect 8899 4156 8955 4212
rect 8981 4156 9037 4212
rect 9063 4156 9119 4212
rect 9145 4156 9201 4212
rect 9227 4156 9283 4212
rect 9308 4156 9364 4212
rect 9389 4156 9445 4212
rect 9470 4156 9526 4212
rect 9551 4156 9607 4212
rect 9632 4156 9688 4212
rect 9713 4156 9769 4212
rect 7587 4076 7643 4132
rect 7669 4076 7725 4132
rect 7751 4076 7807 4132
rect 7833 4076 7889 4132
rect 7915 4076 7971 4132
rect 7997 4076 8053 4132
rect 8079 4076 8135 4132
rect 8161 4076 8217 4132
rect 8243 4076 8299 4132
rect 8325 4076 8381 4132
rect 8407 4076 8463 4132
rect 8489 4076 8545 4132
rect 8571 4076 8627 4132
rect 8653 4076 8709 4132
rect 8735 4076 8791 4132
rect 8817 4076 8873 4132
rect 8899 4076 8955 4132
rect 8981 4076 9037 4132
rect 9063 4076 9119 4132
rect 9145 4076 9201 4132
rect 9227 4076 9283 4132
rect 9308 4076 9364 4132
rect 9389 4076 9445 4132
rect 9470 4076 9526 4132
rect 9551 4076 9607 4132
rect 9632 4076 9688 4132
rect 9713 4076 9769 4132
rect 7587 3996 7643 4052
rect 7669 3996 7725 4052
rect 7751 3996 7807 4052
rect 7833 3996 7889 4052
rect 7915 3996 7971 4052
rect 7997 3996 8053 4052
rect 8079 3996 8135 4052
rect 8161 3996 8217 4052
rect 8243 3996 8299 4052
rect 8325 3996 8381 4052
rect 8407 3996 8463 4052
rect 8489 3996 8545 4052
rect 8571 3996 8627 4052
rect 8653 3996 8709 4052
rect 8735 3996 8791 4052
rect 8817 3996 8873 4052
rect 8899 3996 8955 4052
rect 8981 3996 9037 4052
rect 9063 3996 9119 4052
rect 9145 3996 9201 4052
rect 9227 3996 9283 4052
rect 9308 3996 9364 4052
rect 9389 3996 9445 4052
rect 9470 3996 9526 4052
rect 9551 3996 9607 4052
rect 9632 3996 9688 4052
rect 9713 3996 9769 4052
rect 7587 3916 7643 3972
rect 7669 3916 7725 3972
rect 7751 3916 7807 3972
rect 7833 3916 7889 3972
rect 7915 3916 7971 3972
rect 7997 3916 8053 3972
rect 8079 3916 8135 3972
rect 8161 3916 8217 3972
rect 8243 3916 8299 3972
rect 8325 3916 8381 3972
rect 8407 3916 8463 3972
rect 8489 3916 8545 3972
rect 8571 3916 8627 3972
rect 8653 3916 8709 3972
rect 8735 3916 8791 3972
rect 8817 3916 8873 3972
rect 8899 3916 8955 3972
rect 8981 3916 9037 3972
rect 9063 3916 9119 3972
rect 9145 3916 9201 3972
rect 9227 3916 9283 3972
rect 9308 3916 9364 3972
rect 9389 3916 9445 3972
rect 9470 3916 9526 3972
rect 9551 3916 9607 3972
rect 9632 3916 9688 3972
rect 9713 3916 9769 3972
rect 7587 3836 7643 3892
rect 7669 3836 7725 3892
rect 7751 3836 7807 3892
rect 7833 3836 7889 3892
rect 7915 3836 7971 3892
rect 7997 3836 8053 3892
rect 8079 3836 8135 3892
rect 8161 3836 8217 3892
rect 8243 3836 8299 3892
rect 8325 3836 8381 3892
rect 8407 3836 8463 3892
rect 8489 3836 8545 3892
rect 8571 3836 8627 3892
rect 8653 3836 8709 3892
rect 8735 3836 8791 3892
rect 8817 3836 8873 3892
rect 8899 3836 8955 3892
rect 8981 3836 9037 3892
rect 9063 3836 9119 3892
rect 9145 3836 9201 3892
rect 9227 3836 9283 3892
rect 9308 3836 9364 3892
rect 9389 3836 9445 3892
rect 9470 3836 9526 3892
rect 9551 3836 9607 3892
rect 9632 3836 9688 3892
rect 9713 3836 9769 3892
rect 7587 3756 7643 3812
rect 7669 3756 7725 3812
rect 7751 3756 7807 3812
rect 7833 3756 7889 3812
rect 7915 3756 7971 3812
rect 7997 3756 8053 3812
rect 8079 3756 8135 3812
rect 8161 3756 8217 3812
rect 8243 3756 8299 3812
rect 8325 3756 8381 3812
rect 8407 3756 8463 3812
rect 8489 3756 8545 3812
rect 8571 3756 8627 3812
rect 8653 3756 8709 3812
rect 8735 3756 8791 3812
rect 8817 3756 8873 3812
rect 8899 3756 8955 3812
rect 8981 3756 9037 3812
rect 9063 3756 9119 3812
rect 9145 3756 9201 3812
rect 9227 3756 9283 3812
rect 9308 3756 9364 3812
rect 9389 3756 9445 3812
rect 9470 3756 9526 3812
rect 9551 3756 9607 3812
rect 9632 3756 9688 3812
rect 9713 3756 9769 3812
rect 7587 3676 7643 3732
rect 7669 3676 7725 3732
rect 7751 3676 7807 3732
rect 7833 3676 7889 3732
rect 7915 3676 7971 3732
rect 7997 3676 8053 3732
rect 8079 3676 8135 3732
rect 8161 3676 8217 3732
rect 8243 3676 8299 3732
rect 8325 3676 8381 3732
rect 8407 3676 8463 3732
rect 8489 3676 8545 3732
rect 8571 3676 8627 3732
rect 8653 3676 8709 3732
rect 8735 3676 8791 3732
rect 8817 3676 8873 3732
rect 8899 3676 8955 3732
rect 8981 3676 9037 3732
rect 9063 3676 9119 3732
rect 9145 3676 9201 3732
rect 9227 3676 9283 3732
rect 9308 3676 9364 3732
rect 9389 3676 9445 3732
rect 9470 3676 9526 3732
rect 9551 3676 9607 3732
rect 9632 3676 9688 3732
rect 9713 3676 9769 3732
rect 7587 3596 7643 3652
rect 7669 3596 7725 3652
rect 7751 3596 7807 3652
rect 7833 3596 7889 3652
rect 7915 3596 7971 3652
rect 7997 3596 8053 3652
rect 8079 3596 8135 3652
rect 8161 3596 8217 3652
rect 8243 3596 8299 3652
rect 8325 3596 8381 3652
rect 8407 3596 8463 3652
rect 8489 3596 8545 3652
rect 8571 3596 8627 3652
rect 8653 3596 8709 3652
rect 8735 3596 8791 3652
rect 8817 3596 8873 3652
rect 8899 3596 8955 3652
rect 8981 3596 9037 3652
rect 9063 3596 9119 3652
rect 9145 3596 9201 3652
rect 9227 3596 9283 3652
rect 9308 3596 9364 3652
rect 9389 3596 9445 3652
rect 9470 3596 9526 3652
rect 9551 3596 9607 3652
rect 9632 3596 9688 3652
rect 9713 3596 9769 3652
rect 7587 3516 7643 3572
rect 7669 3516 7725 3572
rect 7751 3516 7807 3572
rect 7833 3516 7889 3572
rect 7915 3516 7971 3572
rect 7997 3516 8053 3572
rect 8079 3516 8135 3572
rect 8161 3516 8217 3572
rect 8243 3516 8299 3572
rect 8325 3516 8381 3572
rect 8407 3516 8463 3572
rect 8489 3516 8545 3572
rect 8571 3516 8627 3572
rect 8653 3516 8709 3572
rect 8735 3516 8791 3572
rect 8817 3516 8873 3572
rect 8899 3516 8955 3572
rect 8981 3516 9037 3572
rect 9063 3516 9119 3572
rect 9145 3516 9201 3572
rect 9227 3516 9283 3572
rect 9308 3516 9364 3572
rect 9389 3516 9445 3572
rect 9470 3516 9526 3572
rect 9551 3516 9607 3572
rect 9632 3516 9688 3572
rect 9713 3516 9769 3572
rect 7587 3436 7643 3492
rect 7669 3436 7725 3492
rect 7751 3436 7807 3492
rect 7833 3436 7889 3492
rect 7915 3436 7971 3492
rect 7997 3436 8053 3492
rect 8079 3436 8135 3492
rect 8161 3436 8217 3492
rect 8243 3436 8299 3492
rect 8325 3436 8381 3492
rect 8407 3436 8463 3492
rect 8489 3436 8545 3492
rect 8571 3436 8627 3492
rect 8653 3436 8709 3492
rect 8735 3436 8791 3492
rect 8817 3436 8873 3492
rect 8899 3436 8955 3492
rect 8981 3436 9037 3492
rect 9063 3436 9119 3492
rect 9145 3436 9201 3492
rect 9227 3436 9283 3492
rect 9308 3436 9364 3492
rect 9389 3436 9445 3492
rect 9470 3436 9526 3492
rect 9551 3436 9607 3492
rect 9632 3436 9688 3492
rect 9713 3436 9769 3492
rect 7587 3356 7643 3412
rect 7669 3356 7725 3412
rect 7751 3356 7807 3412
rect 7833 3356 7889 3412
rect 7915 3356 7971 3412
rect 7997 3356 8053 3412
rect 8079 3356 8135 3412
rect 8161 3356 8217 3412
rect 8243 3356 8299 3412
rect 8325 3356 8381 3412
rect 8407 3356 8463 3412
rect 8489 3356 8545 3412
rect 8571 3356 8627 3412
rect 8653 3356 8709 3412
rect 8735 3356 8791 3412
rect 8817 3356 8873 3412
rect 8899 3356 8955 3412
rect 8981 3356 9037 3412
rect 9063 3356 9119 3412
rect 9145 3356 9201 3412
rect 9227 3356 9283 3412
rect 9308 3356 9364 3412
rect 9389 3356 9445 3412
rect 9470 3356 9526 3412
rect 9551 3356 9607 3412
rect 9632 3356 9688 3412
rect 9713 3356 9769 3412
rect 7587 3276 7643 3332
rect 7669 3276 7725 3332
rect 7751 3276 7807 3332
rect 7833 3276 7889 3332
rect 7915 3276 7971 3332
rect 7997 3276 8053 3332
rect 8079 3276 8135 3332
rect 8161 3276 8217 3332
rect 8243 3276 8299 3332
rect 8325 3276 8381 3332
rect 8407 3276 8463 3332
rect 8489 3276 8545 3332
rect 8571 3276 8627 3332
rect 8653 3276 8709 3332
rect 8735 3276 8791 3332
rect 8817 3276 8873 3332
rect 8899 3276 8955 3332
rect 8981 3276 9037 3332
rect 9063 3276 9119 3332
rect 9145 3276 9201 3332
rect 9227 3276 9283 3332
rect 9308 3276 9364 3332
rect 9389 3276 9445 3332
rect 9470 3276 9526 3332
rect 9551 3276 9607 3332
rect 9632 3276 9688 3332
rect 9713 3276 9769 3332
rect 7587 3196 7643 3252
rect 7669 3196 7725 3252
rect 7751 3196 7807 3252
rect 7833 3196 7889 3252
rect 7915 3196 7971 3252
rect 7997 3196 8053 3252
rect 8079 3196 8135 3252
rect 8161 3196 8217 3252
rect 8243 3196 8299 3252
rect 8325 3196 8381 3252
rect 8407 3196 8463 3252
rect 8489 3196 8545 3252
rect 8571 3196 8627 3252
rect 8653 3196 8709 3252
rect 8735 3196 8791 3252
rect 8817 3196 8873 3252
rect 8899 3196 8955 3252
rect 8981 3196 9037 3252
rect 9063 3196 9119 3252
rect 9145 3196 9201 3252
rect 9227 3196 9283 3252
rect 9308 3196 9364 3252
rect 9389 3196 9445 3252
rect 9470 3196 9526 3252
rect 9551 3196 9607 3252
rect 9632 3196 9688 3252
rect 9713 3196 9769 3252
rect 7587 3116 7643 3172
rect 7669 3116 7725 3172
rect 7751 3116 7807 3172
rect 7833 3116 7889 3172
rect 7915 3116 7971 3172
rect 7997 3116 8053 3172
rect 8079 3116 8135 3172
rect 8161 3116 8217 3172
rect 8243 3116 8299 3172
rect 8325 3116 8381 3172
rect 8407 3116 8463 3172
rect 8489 3116 8545 3172
rect 8571 3116 8627 3172
rect 8653 3116 8709 3172
rect 8735 3116 8791 3172
rect 8817 3116 8873 3172
rect 8899 3116 8955 3172
rect 8981 3116 9037 3172
rect 9063 3116 9119 3172
rect 9145 3116 9201 3172
rect 9227 3116 9283 3172
rect 9308 3116 9364 3172
rect 9389 3116 9445 3172
rect 9470 3116 9526 3172
rect 9551 3116 9607 3172
rect 9632 3116 9688 3172
rect 9713 3116 9769 3172
rect 7587 3036 7643 3092
rect 7669 3036 7725 3092
rect 7751 3036 7807 3092
rect 7833 3036 7889 3092
rect 7915 3036 7971 3092
rect 7997 3036 8053 3092
rect 8079 3036 8135 3092
rect 8161 3036 8217 3092
rect 8243 3036 8299 3092
rect 8325 3036 8381 3092
rect 8407 3036 8463 3092
rect 8489 3036 8545 3092
rect 8571 3036 8627 3092
rect 8653 3036 8709 3092
rect 8735 3036 8791 3092
rect 8817 3036 8873 3092
rect 8899 3036 8955 3092
rect 8981 3036 9037 3092
rect 9063 3036 9119 3092
rect 9145 3036 9201 3092
rect 9227 3036 9283 3092
rect 9308 3036 9364 3092
rect 9389 3036 9445 3092
rect 9470 3036 9526 3092
rect 9551 3036 9607 3092
rect 9632 3036 9688 3092
rect 9713 3036 9769 3092
rect 7587 2956 7643 3012
rect 7669 2956 7725 3012
rect 7751 2956 7807 3012
rect 7833 2956 7889 3012
rect 7915 2956 7971 3012
rect 7997 2956 8053 3012
rect 8079 2956 8135 3012
rect 8161 2956 8217 3012
rect 8243 2956 8299 3012
rect 8325 2956 8381 3012
rect 8407 2956 8463 3012
rect 8489 2956 8545 3012
rect 8571 2956 8627 3012
rect 8653 2956 8709 3012
rect 8735 2956 8791 3012
rect 8817 2956 8873 3012
rect 8899 2956 8955 3012
rect 8981 2956 9037 3012
rect 9063 2956 9119 3012
rect 9145 2956 9201 3012
rect 9227 2956 9283 3012
rect 9308 2956 9364 3012
rect 9389 2956 9445 3012
rect 9470 2956 9526 3012
rect 9551 2956 9607 3012
rect 9632 2956 9688 3012
rect 9713 2956 9769 3012
rect 7587 2876 7643 2932
rect 7669 2876 7725 2932
rect 7751 2876 7807 2932
rect 7833 2876 7889 2932
rect 7915 2876 7971 2932
rect 7997 2876 8053 2932
rect 8079 2876 8135 2932
rect 8161 2876 8217 2932
rect 8243 2876 8299 2932
rect 8325 2876 8381 2932
rect 8407 2876 8463 2932
rect 8489 2876 8545 2932
rect 8571 2876 8627 2932
rect 8653 2876 8709 2932
rect 8735 2876 8791 2932
rect 8817 2876 8873 2932
rect 8899 2876 8955 2932
rect 8981 2876 9037 2932
rect 9063 2876 9119 2932
rect 9145 2876 9201 2932
rect 9227 2876 9283 2932
rect 9308 2876 9364 2932
rect 9389 2876 9445 2932
rect 9470 2876 9526 2932
rect 9551 2876 9607 2932
rect 9632 2876 9688 2932
rect 9713 2876 9769 2932
rect 7587 2796 7643 2852
rect 7669 2796 7725 2852
rect 7751 2796 7807 2852
rect 7833 2796 7889 2852
rect 7915 2796 7971 2852
rect 7997 2796 8053 2852
rect 8079 2796 8135 2852
rect 8161 2796 8217 2852
rect 8243 2796 8299 2852
rect 8325 2796 8381 2852
rect 8407 2796 8463 2852
rect 8489 2796 8545 2852
rect 8571 2796 8627 2852
rect 8653 2796 8709 2852
rect 8735 2796 8791 2852
rect 8817 2796 8873 2852
rect 8899 2796 8955 2852
rect 8981 2796 9037 2852
rect 9063 2796 9119 2852
rect 9145 2796 9201 2852
rect 9227 2796 9283 2852
rect 9308 2796 9364 2852
rect 9389 2796 9445 2852
rect 9470 2796 9526 2852
rect 9551 2796 9607 2852
rect 9632 2796 9688 2852
rect 9713 2796 9769 2852
rect 7587 2716 7643 2772
rect 7669 2716 7725 2772
rect 7751 2716 7807 2772
rect 7833 2716 7889 2772
rect 7915 2716 7971 2772
rect 7997 2716 8053 2772
rect 8079 2716 8135 2772
rect 8161 2716 8217 2772
rect 8243 2716 8299 2772
rect 8325 2716 8381 2772
rect 8407 2716 8463 2772
rect 8489 2716 8545 2772
rect 8571 2716 8627 2772
rect 8653 2716 8709 2772
rect 8735 2716 8791 2772
rect 8817 2716 8873 2772
rect 8899 2716 8955 2772
rect 8981 2716 9037 2772
rect 9063 2716 9119 2772
rect 9145 2716 9201 2772
rect 9227 2716 9283 2772
rect 9308 2716 9364 2772
rect 9389 2716 9445 2772
rect 9470 2716 9526 2772
rect 9551 2716 9607 2772
rect 9632 2716 9688 2772
rect 9713 2716 9769 2772
rect 7587 2636 7643 2692
rect 7669 2636 7725 2692
rect 7751 2636 7807 2692
rect 7833 2636 7889 2692
rect 7915 2636 7971 2692
rect 7997 2636 8053 2692
rect 8079 2636 8135 2692
rect 8161 2636 8217 2692
rect 8243 2636 8299 2692
rect 8325 2636 8381 2692
rect 8407 2636 8463 2692
rect 8489 2636 8545 2692
rect 8571 2636 8627 2692
rect 8653 2636 8709 2692
rect 8735 2636 8791 2692
rect 8817 2636 8873 2692
rect 8899 2636 8955 2692
rect 8981 2636 9037 2692
rect 9063 2636 9119 2692
rect 9145 2636 9201 2692
rect 9227 2636 9283 2692
rect 9308 2636 9364 2692
rect 9389 2636 9445 2692
rect 9470 2636 9526 2692
rect 9551 2636 9607 2692
rect 9632 2636 9688 2692
rect 9713 2636 9769 2692
rect 7587 2556 7643 2612
rect 7669 2556 7725 2612
rect 7751 2556 7807 2612
rect 7833 2556 7889 2612
rect 7915 2556 7971 2612
rect 7997 2556 8053 2612
rect 8079 2556 8135 2612
rect 8161 2556 8217 2612
rect 8243 2556 8299 2612
rect 8325 2556 8381 2612
rect 8407 2556 8463 2612
rect 8489 2556 8545 2612
rect 8571 2556 8627 2612
rect 8653 2556 8709 2612
rect 8735 2556 8791 2612
rect 8817 2556 8873 2612
rect 8899 2556 8955 2612
rect 8981 2556 9037 2612
rect 9063 2556 9119 2612
rect 9145 2556 9201 2612
rect 9227 2556 9283 2612
rect 9308 2556 9364 2612
rect 9389 2556 9445 2612
rect 9470 2556 9526 2612
rect 9551 2556 9607 2612
rect 9632 2556 9688 2612
rect 9713 2556 9769 2612
rect 7587 2476 7643 2532
rect 7669 2476 7725 2532
rect 7751 2476 7807 2532
rect 7833 2476 7889 2532
rect 7915 2476 7971 2532
rect 7997 2476 8053 2532
rect 8079 2476 8135 2532
rect 8161 2476 8217 2532
rect 8243 2476 8299 2532
rect 8325 2476 8381 2532
rect 8407 2476 8463 2532
rect 8489 2476 8545 2532
rect 8571 2476 8627 2532
rect 8653 2476 8709 2532
rect 8735 2476 8791 2532
rect 8817 2476 8873 2532
rect 8899 2476 8955 2532
rect 8981 2476 9037 2532
rect 9063 2476 9119 2532
rect 9145 2476 9201 2532
rect 9227 2476 9283 2532
rect 9308 2476 9364 2532
rect 9389 2476 9445 2532
rect 9470 2476 9526 2532
rect 9551 2476 9607 2532
rect 9632 2476 9688 2532
rect 9713 2476 9769 2532
<< metal3 >>
rect 2525 39009 5002 39015
rect 2525 38953 2534 39009
rect 2590 38953 2617 39009
rect 2673 38953 2700 39009
rect 2756 38953 2783 39009
rect 2839 38953 2866 39009
rect 2922 38953 2949 39009
rect 3005 38953 3032 39009
rect 3088 38953 3115 39009
rect 3171 38953 3198 39009
rect 3254 38953 3281 39009
rect 3337 38953 3364 39009
rect 3420 38953 3447 39009
rect 3503 38953 3530 39009
rect 3586 38953 3613 39009
rect 3669 38953 3696 39009
rect 3752 38953 3779 39009
rect 3835 38953 3862 39009
rect 3918 38953 3945 39009
rect 4001 38953 4028 39009
rect 4084 38953 4111 39009
rect 4167 38953 4194 39009
rect 4250 38953 4276 39009
rect 4332 38953 4358 39009
rect 4414 38953 4440 39009
rect 4496 38953 4522 39009
rect 4578 38953 4604 39009
rect 4660 38953 4686 39009
rect 4742 38953 4768 39009
rect 4824 38953 4850 39009
rect 4906 38953 4932 39009
rect 4988 38953 5002 39009
rect 2525 38925 5002 38953
rect 2525 38869 2534 38925
rect 2590 38869 2617 38925
rect 2673 38869 2700 38925
rect 2756 38869 2783 38925
rect 2839 38869 2866 38925
rect 2922 38869 2949 38925
rect 3005 38869 3032 38925
rect 3088 38869 3115 38925
rect 3171 38869 3198 38925
rect 3254 38869 3281 38925
rect 3337 38869 3364 38925
rect 3420 38869 3447 38925
rect 3503 38869 3530 38925
rect 3586 38869 3613 38925
rect 3669 38869 3696 38925
rect 3752 38869 3779 38925
rect 3835 38869 3862 38925
rect 3918 38869 3945 38925
rect 4001 38869 4028 38925
rect 4084 38869 4111 38925
rect 4167 38869 4194 38925
rect 4250 38869 4276 38925
rect 4332 38869 4358 38925
rect 4414 38869 4440 38925
rect 4496 38869 4522 38925
rect 4578 38869 4604 38925
rect 4660 38869 4686 38925
rect 4742 38869 4768 38925
rect 4824 38869 4850 38925
rect 4906 38869 4932 38925
rect 4988 38869 5002 38925
rect 2525 38841 5002 38869
rect 2525 38785 2534 38841
rect 2590 38785 2617 38841
rect 2673 38785 2700 38841
rect 2756 38785 2783 38841
rect 2839 38785 2866 38841
rect 2922 38785 2949 38841
rect 3005 38785 3032 38841
rect 3088 38785 3115 38841
rect 3171 38785 3198 38841
rect 3254 38785 3281 38841
rect 3337 38785 3364 38841
rect 3420 38785 3447 38841
rect 3503 38785 3530 38841
rect 3586 38785 3613 38841
rect 3669 38785 3696 38841
rect 3752 38785 3779 38841
rect 3835 38785 3862 38841
rect 3918 38785 3945 38841
rect 4001 38785 4028 38841
rect 4084 38785 4111 38841
rect 4167 38785 4194 38841
rect 4250 38785 4276 38841
rect 4332 38785 4358 38841
rect 4414 38785 4440 38841
rect 4496 38785 4522 38841
rect 4578 38785 4604 38841
rect 4660 38785 4686 38841
rect 4742 38785 4768 38841
rect 4824 38785 4850 38841
rect 4906 38785 4932 38841
rect 4988 38785 5002 38841
rect 2525 38757 5002 38785
rect 2525 38701 2534 38757
rect 2590 38701 2617 38757
rect 2673 38701 2700 38757
rect 2756 38701 2783 38757
rect 2839 38701 2866 38757
rect 2922 38701 2949 38757
rect 3005 38701 3032 38757
rect 3088 38701 3115 38757
rect 3171 38701 3198 38757
rect 3254 38701 3281 38757
rect 3337 38701 3364 38757
rect 3420 38701 3447 38757
rect 3503 38701 3530 38757
rect 3586 38701 3613 38757
rect 3669 38701 3696 38757
rect 3752 38701 3779 38757
rect 3835 38701 3862 38757
rect 3918 38701 3945 38757
rect 4001 38701 4028 38757
rect 4084 38701 4111 38757
rect 4167 38701 4194 38757
rect 4250 38701 4276 38757
rect 4332 38701 4358 38757
rect 4414 38701 4440 38757
rect 4496 38701 4522 38757
rect 4578 38701 4604 38757
rect 4660 38701 4686 38757
rect 4742 38701 4768 38757
rect 4824 38701 4850 38757
rect 4906 38701 4932 38757
rect 4988 38701 5002 38757
rect 2525 38673 5002 38701
rect 2525 38617 2534 38673
rect 2590 38617 2617 38673
rect 2673 38617 2700 38673
rect 2756 38617 2783 38673
rect 2839 38617 2866 38673
rect 2922 38617 2949 38673
rect 3005 38617 3032 38673
rect 3088 38617 3115 38673
rect 3171 38617 3198 38673
rect 3254 38617 3281 38673
rect 3337 38617 3364 38673
rect 3420 38617 3447 38673
rect 3503 38617 3530 38673
rect 3586 38617 3613 38673
rect 3669 38617 3696 38673
rect 3752 38617 3779 38673
rect 3835 38617 3862 38673
rect 3918 38617 3945 38673
rect 4001 38617 4028 38673
rect 4084 38617 4111 38673
rect 4167 38617 4194 38673
rect 4250 38617 4276 38673
rect 4332 38617 4358 38673
rect 4414 38617 4440 38673
rect 4496 38617 4522 38673
rect 4578 38617 4604 38673
rect 4660 38617 4686 38673
rect 4742 38617 4768 38673
rect 4824 38617 4850 38673
rect 4906 38617 4932 38673
rect 4988 38617 5002 38673
rect 2525 38589 5002 38617
rect 2525 38533 2534 38589
rect 2590 38533 2617 38589
rect 2673 38533 2700 38589
rect 2756 38533 2783 38589
rect 2839 38533 2866 38589
rect 2922 38533 2949 38589
rect 3005 38533 3032 38589
rect 3088 38533 3115 38589
rect 3171 38533 3198 38589
rect 3254 38533 3281 38589
rect 3337 38533 3364 38589
rect 3420 38533 3447 38589
rect 3503 38533 3530 38589
rect 3586 38533 3613 38589
rect 3669 38533 3696 38589
rect 3752 38533 3779 38589
rect 3835 38533 3862 38589
rect 3918 38533 3945 38589
rect 4001 38533 4028 38589
rect 4084 38533 4111 38589
rect 4167 38533 4194 38589
rect 4250 38533 4276 38589
rect 4332 38533 4358 38589
rect 4414 38533 4440 38589
rect 4496 38533 4522 38589
rect 4578 38533 4604 38589
rect 4660 38533 4686 38589
rect 4742 38533 4768 38589
rect 4824 38533 4850 38589
rect 4906 38533 4932 38589
rect 4988 38533 5002 38589
rect 2525 38505 5002 38533
rect 2525 38449 2534 38505
rect 2590 38449 2617 38505
rect 2673 38449 2700 38505
rect 2756 38449 2783 38505
rect 2839 38449 2866 38505
rect 2922 38449 2949 38505
rect 3005 38449 3032 38505
rect 3088 38449 3115 38505
rect 3171 38449 3198 38505
rect 3254 38449 3281 38505
rect 3337 38449 3364 38505
rect 3420 38449 3447 38505
rect 3503 38449 3530 38505
rect 3586 38449 3613 38505
rect 3669 38449 3696 38505
rect 3752 38449 3779 38505
rect 3835 38449 3862 38505
rect 3918 38449 3945 38505
rect 4001 38449 4028 38505
rect 4084 38449 4111 38505
rect 4167 38449 4194 38505
rect 4250 38449 4276 38505
rect 4332 38449 4358 38505
rect 4414 38449 4440 38505
rect 4496 38449 4522 38505
rect 4578 38449 4604 38505
rect 4660 38449 4686 38505
rect 4742 38449 4768 38505
rect 4824 38449 4850 38505
rect 4906 38449 4932 38505
rect 4988 38449 5002 38505
rect 2525 38421 5002 38449
rect 2525 38365 2534 38421
rect 2590 38365 2617 38421
rect 2673 38365 2700 38421
rect 2756 38365 2783 38421
rect 2839 38365 2866 38421
rect 2922 38365 2949 38421
rect 3005 38365 3032 38421
rect 3088 38365 3115 38421
rect 3171 38365 3198 38421
rect 3254 38365 3281 38421
rect 3337 38365 3364 38421
rect 3420 38365 3447 38421
rect 3503 38365 3530 38421
rect 3586 38365 3613 38421
rect 3669 38365 3696 38421
rect 3752 38365 3779 38421
rect 3835 38365 3862 38421
rect 3918 38365 3945 38421
rect 4001 38365 4028 38421
rect 4084 38365 4111 38421
rect 4167 38365 4194 38421
rect 4250 38365 4276 38421
rect 4332 38365 4358 38421
rect 4414 38365 4440 38421
rect 4496 38365 4522 38421
rect 4578 38365 4604 38421
rect 4660 38365 4686 38421
rect 4742 38365 4768 38421
rect 4824 38365 4850 38421
rect 4906 38365 4932 38421
rect 4988 38365 5002 38421
rect 2525 38337 5002 38365
rect 2525 38281 2534 38337
rect 2590 38281 2617 38337
rect 2673 38281 2700 38337
rect 2756 38281 2783 38337
rect 2839 38281 2866 38337
rect 2922 38281 2949 38337
rect 3005 38281 3032 38337
rect 3088 38281 3115 38337
rect 3171 38281 3198 38337
rect 3254 38281 3281 38337
rect 3337 38281 3364 38337
rect 3420 38281 3447 38337
rect 3503 38281 3530 38337
rect 3586 38281 3613 38337
rect 3669 38281 3696 38337
rect 3752 38281 3779 38337
rect 3835 38281 3862 38337
rect 3918 38281 3945 38337
rect 4001 38281 4028 38337
rect 4084 38281 4111 38337
rect 4167 38281 4194 38337
rect 4250 38281 4276 38337
rect 4332 38281 4358 38337
rect 4414 38281 4440 38337
rect 4496 38281 4522 38337
rect 4578 38281 4604 38337
rect 4660 38281 4686 38337
rect 4742 38281 4768 38337
rect 4824 38281 4850 38337
rect 4906 38281 4932 38337
rect 4988 38281 5002 38337
rect 2525 38253 5002 38281
rect 2525 38197 2534 38253
rect 2590 38197 2617 38253
rect 2673 38197 2700 38253
rect 2756 38197 2783 38253
rect 2839 38197 2866 38253
rect 2922 38197 2949 38253
rect 3005 38197 3032 38253
rect 3088 38197 3115 38253
rect 3171 38197 3198 38253
rect 3254 38197 3281 38253
rect 3337 38197 3364 38253
rect 3420 38197 3447 38253
rect 3503 38197 3530 38253
rect 3586 38197 3613 38253
rect 3669 38197 3696 38253
rect 3752 38197 3779 38253
rect 3835 38197 3862 38253
rect 3918 38197 3945 38253
rect 4001 38197 4028 38253
rect 4084 38197 4111 38253
rect 4167 38197 4194 38253
rect 4250 38197 4276 38253
rect 4332 38197 4358 38253
rect 4414 38197 4440 38253
rect 4496 38197 4522 38253
rect 4578 38197 4604 38253
rect 4660 38197 4686 38253
rect 4742 38197 4768 38253
rect 4824 38197 4850 38253
rect 4906 38197 4932 38253
rect 4988 38197 5002 38253
rect 2525 38169 5002 38197
rect 2525 38113 2534 38169
rect 2590 38113 2617 38169
rect 2673 38113 2700 38169
rect 2756 38113 2783 38169
rect 2839 38113 2866 38169
rect 2922 38113 2949 38169
rect 3005 38113 3032 38169
rect 3088 38113 3115 38169
rect 3171 38113 3198 38169
rect 3254 38113 3281 38169
rect 3337 38113 3364 38169
rect 3420 38113 3447 38169
rect 3503 38113 3530 38169
rect 3586 38113 3613 38169
rect 3669 38113 3696 38169
rect 3752 38113 3779 38169
rect 3835 38113 3862 38169
rect 3918 38113 3945 38169
rect 4001 38113 4028 38169
rect 4084 38113 4111 38169
rect 4167 38113 4194 38169
rect 4250 38113 4276 38169
rect 4332 38113 4358 38169
rect 4414 38113 4440 38169
rect 4496 38113 4522 38169
rect 4578 38113 4604 38169
rect 4660 38113 4686 38169
rect 4742 38113 4768 38169
rect 4824 38113 4850 38169
rect 4906 38113 4932 38169
rect 4988 38113 5002 38169
rect 2525 38073 5002 38113
rect 2525 38017 2531 38073
rect 2587 38017 2649 38073
rect 2705 38017 2767 38073
rect 2823 38017 5002 38073
rect 2525 37988 5002 38017
rect 2525 37932 2531 37988
rect 2587 37932 2649 37988
rect 2705 37932 2767 37988
rect 2823 37932 5002 37988
rect 2525 37903 5002 37932
rect 2525 37847 2531 37903
rect 2587 37847 2649 37903
rect 2705 37847 2767 37903
rect 2823 37847 5002 37903
rect 2525 37818 5002 37847
rect 2525 37762 2531 37818
rect 2587 37762 2649 37818
rect 2705 37762 2767 37818
rect 2823 37762 5002 37818
rect 2525 37733 5002 37762
rect 2525 37677 2531 37733
rect 2587 37677 2649 37733
rect 2705 37677 2767 37733
rect 2823 37677 5002 37733
rect 2525 37648 5002 37677
rect 2525 37592 2531 37648
rect 2587 37592 2649 37648
rect 2705 37592 2767 37648
rect 2823 37592 5002 37648
rect 2525 37563 5002 37592
rect 2525 37507 2531 37563
rect 2587 37507 2649 37563
rect 2705 37507 2767 37563
rect 2823 37507 5002 37563
rect 2525 37478 5002 37507
rect 2525 37422 2531 37478
rect 2587 37422 2649 37478
rect 2705 37422 2767 37478
rect 2823 37422 5002 37478
rect 2525 37393 5002 37422
rect 2525 37337 2531 37393
rect 2587 37337 2649 37393
rect 2705 37337 2767 37393
rect 2823 37337 5002 37393
rect 2525 37308 5002 37337
rect 2525 37252 2531 37308
rect 2587 37252 2649 37308
rect 2705 37252 2767 37308
rect 2823 37252 5002 37308
rect 2525 37222 5002 37252
rect 2525 37166 2531 37222
rect 2587 37166 2649 37222
rect 2705 37166 2767 37222
rect 2823 37166 5002 37222
rect 2525 37136 5002 37166
rect 2525 37080 2531 37136
rect 2587 37080 2649 37136
rect 2705 37080 2767 37136
rect 2823 37080 5002 37136
rect 2525 37050 5002 37080
rect 2525 36994 2531 37050
rect 2587 36994 2649 37050
rect 2705 36994 2767 37050
rect 2823 36994 5002 37050
rect 2525 36964 5002 36994
rect 2525 36908 2531 36964
rect 2587 36908 2649 36964
rect 2705 36908 2767 36964
rect 2823 36908 5002 36964
rect 2525 36878 5002 36908
rect 2525 36822 2531 36878
rect 2587 36822 2649 36878
rect 2705 36822 2767 36878
rect 2823 36822 5002 36878
rect 2525 36772 5002 36822
rect 2525 36716 2538 36772
rect 2594 36716 2632 36772
rect 2688 36716 2726 36772
rect 2782 36716 2820 36772
rect 2876 36716 2914 36772
rect 2970 36716 3008 36772
rect 3064 36716 5002 36772
rect 2525 36692 5002 36716
rect 2525 36636 2538 36692
rect 2594 36636 2632 36692
rect 2688 36636 2726 36692
rect 2782 36636 2820 36692
rect 2876 36636 2914 36692
rect 2970 36636 3008 36692
rect 3064 36650 5002 36692
rect 3064 36636 3099 36650
rect 2525 36612 3099 36636
rect 2525 36556 2538 36612
rect 2594 36556 2632 36612
rect 2688 36556 2726 36612
rect 2782 36556 2820 36612
rect 2876 36556 2914 36612
rect 2970 36556 3008 36612
rect 3064 36594 3099 36612
rect 3155 36594 5002 36650
rect 3064 36562 5002 36594
rect 3064 36556 3112 36562
rect 2525 36532 3112 36556
rect 2525 36476 2538 36532
rect 2594 36476 2632 36532
rect 2688 36476 2726 36532
rect 2782 36476 2820 36532
rect 2876 36476 2914 36532
rect 2970 36476 3008 36532
rect 3064 36506 3112 36532
rect 3168 36506 3206 36562
rect 3262 36506 5002 36562
rect 3064 36476 5002 36506
rect 2525 36452 3112 36476
rect 2525 36396 2538 36452
rect 2594 36396 2632 36452
rect 2688 36396 2726 36452
rect 2782 36396 2820 36452
rect 2876 36396 2914 36452
rect 2970 36396 3008 36452
rect 3064 36420 3112 36452
rect 3168 36420 3206 36476
rect 3262 36420 5002 36476
rect 3064 36415 5002 36420
rect 3064 36396 3321 36415
rect 2525 36390 3321 36396
rect 2525 36372 3112 36390
rect 2525 36316 2538 36372
rect 2594 36316 2632 36372
rect 2688 36316 2726 36372
rect 2782 36316 2820 36372
rect 2876 36316 2914 36372
rect 2970 36316 3008 36372
rect 3064 36334 3112 36372
rect 3168 36334 3206 36390
rect 3262 36359 3321 36390
rect 3377 36359 5002 36415
rect 3262 36334 5002 36359
rect 3064 36316 5002 36334
rect 2525 36294 5002 36316
rect 2525 36292 3109 36294
rect 2525 36236 2538 36292
rect 2594 36236 2632 36292
rect 2688 36236 2726 36292
rect 2782 36236 2820 36292
rect 2876 36236 2914 36292
rect 2970 36236 3008 36292
rect 3064 36238 3109 36292
rect 3165 36238 3193 36294
rect 3249 36238 3277 36294
rect 3333 36238 3360 36294
rect 3416 36238 3443 36294
rect 3499 36238 3526 36294
rect 3582 36238 3609 36294
rect 3665 36238 3692 36294
rect 3748 36238 3775 36294
rect 3831 36238 3858 36294
rect 3914 36238 3941 36294
rect 3997 36238 4024 36294
rect 4080 36238 4107 36294
rect 4163 36238 4190 36294
rect 4246 36238 4273 36294
rect 4329 36238 4356 36294
rect 4412 36238 4439 36294
rect 4495 36238 4522 36294
rect 4578 36238 4605 36294
rect 4661 36238 4688 36294
rect 4744 36238 4771 36294
rect 4827 36238 4854 36294
rect 4910 36238 4937 36294
rect 4993 36238 5002 36294
rect 3064 36236 5002 36238
rect 2525 36214 5002 36236
rect 2525 36212 3109 36214
rect 2525 36156 2538 36212
rect 2594 36156 2632 36212
rect 2688 36156 2726 36212
rect 2782 36156 2820 36212
rect 2876 36156 2914 36212
rect 2970 36156 3008 36212
rect 3064 36158 3109 36212
rect 3165 36158 3193 36214
rect 3249 36158 3277 36214
rect 3333 36158 3360 36214
rect 3416 36158 3443 36214
rect 3499 36158 3526 36214
rect 3582 36158 3609 36214
rect 3665 36158 3692 36214
rect 3748 36158 3775 36214
rect 3831 36158 3858 36214
rect 3914 36158 3941 36214
rect 3997 36158 4024 36214
rect 4080 36158 4107 36214
rect 4163 36158 4190 36214
rect 4246 36158 4273 36214
rect 4329 36158 4356 36214
rect 4412 36158 4439 36214
rect 4495 36158 4522 36214
rect 4578 36158 4605 36214
rect 4661 36158 4688 36214
rect 4744 36158 4771 36214
rect 4827 36158 4854 36214
rect 4910 36158 4937 36214
rect 4993 36158 5002 36214
rect 3064 36156 5002 36158
rect 2525 36134 5002 36156
rect 2525 36132 3109 36134
rect 2525 36076 2538 36132
rect 2594 36076 2632 36132
rect 2688 36076 2726 36132
rect 2782 36076 2820 36132
rect 2876 36076 2914 36132
rect 2970 36076 3008 36132
rect 3064 36078 3109 36132
rect 3165 36078 3193 36134
rect 3249 36078 3277 36134
rect 3333 36078 3360 36134
rect 3416 36078 3443 36134
rect 3499 36078 3526 36134
rect 3582 36078 3609 36134
rect 3665 36078 3692 36134
rect 3748 36078 3775 36134
rect 3831 36078 3858 36134
rect 3914 36078 3941 36134
rect 3997 36078 4024 36134
rect 4080 36078 4107 36134
rect 4163 36078 4190 36134
rect 4246 36078 4273 36134
rect 4329 36078 4356 36134
rect 4412 36078 4439 36134
rect 4495 36078 4522 36134
rect 4578 36078 4605 36134
rect 4661 36078 4688 36134
rect 4744 36078 4771 36134
rect 4827 36078 4854 36134
rect 4910 36078 4937 36134
rect 4993 36078 5002 36134
rect 3064 36076 5002 36078
rect 2525 36054 5002 36076
rect 2525 36052 3109 36054
rect 2525 35996 2538 36052
rect 2594 35996 2632 36052
rect 2688 35996 2726 36052
rect 2782 35996 2820 36052
rect 2876 35996 2914 36052
rect 2970 35996 3008 36052
rect 3064 35998 3109 36052
rect 3165 35998 3193 36054
rect 3249 35998 3277 36054
rect 3333 35998 3360 36054
rect 3416 35998 3443 36054
rect 3499 35998 3526 36054
rect 3582 35998 3609 36054
rect 3665 35998 3692 36054
rect 3748 35998 3775 36054
rect 3831 35998 3858 36054
rect 3914 35998 3941 36054
rect 3997 35998 4024 36054
rect 4080 35998 4107 36054
rect 4163 35998 4190 36054
rect 4246 35998 4273 36054
rect 4329 35998 4356 36054
rect 4412 35998 4439 36054
rect 4495 35998 4522 36054
rect 4578 35998 4605 36054
rect 4661 35998 4688 36054
rect 4744 35998 4771 36054
rect 4827 35998 4854 36054
rect 4910 35998 4937 36054
rect 4993 35998 5002 36054
rect 3064 35996 5002 35998
rect 2525 35974 5002 35996
rect 2525 35972 3109 35974
rect 2525 35916 2538 35972
rect 2594 35916 2632 35972
rect 2688 35916 2726 35972
rect 2782 35916 2820 35972
rect 2876 35916 2914 35972
rect 2970 35916 3008 35972
rect 3064 35918 3109 35972
rect 3165 35918 3193 35974
rect 3249 35918 3277 35974
rect 3333 35918 3360 35974
rect 3416 35918 3443 35974
rect 3499 35918 3526 35974
rect 3582 35918 3609 35974
rect 3665 35918 3692 35974
rect 3748 35918 3775 35974
rect 3831 35918 3858 35974
rect 3914 35918 3941 35974
rect 3997 35918 4024 35974
rect 4080 35918 4107 35974
rect 4163 35918 4190 35974
rect 4246 35918 4273 35974
rect 4329 35918 4356 35974
rect 4412 35918 4439 35974
rect 4495 35918 4522 35974
rect 4578 35918 4605 35974
rect 4661 35918 4688 35974
rect 4744 35918 4771 35974
rect 4827 35918 4854 35974
rect 4910 35918 4937 35974
rect 4993 35918 5002 35974
rect 3064 35916 5002 35918
rect 2525 35894 5002 35916
rect 2525 35892 3109 35894
rect 2525 35836 2538 35892
rect 2594 35836 2632 35892
rect 2688 35836 2726 35892
rect 2782 35836 2820 35892
rect 2876 35836 2914 35892
rect 2970 35836 3008 35892
rect 3064 35838 3109 35892
rect 3165 35838 3193 35894
rect 3249 35838 3277 35894
rect 3333 35838 3360 35894
rect 3416 35838 3443 35894
rect 3499 35838 3526 35894
rect 3582 35838 3609 35894
rect 3665 35838 3692 35894
rect 3748 35838 3775 35894
rect 3831 35838 3858 35894
rect 3914 35838 3941 35894
rect 3997 35838 4024 35894
rect 4080 35838 4107 35894
rect 4163 35838 4190 35894
rect 4246 35838 4273 35894
rect 4329 35838 4356 35894
rect 4412 35838 4439 35894
rect 4495 35838 4522 35894
rect 4578 35838 4605 35894
rect 4661 35838 4688 35894
rect 4744 35838 4771 35894
rect 4827 35838 4854 35894
rect 4910 35838 4937 35894
rect 4993 35838 5002 35894
rect 3064 35836 5002 35838
rect 2525 35814 5002 35836
rect 2525 35812 3109 35814
rect 2525 35756 2538 35812
rect 2594 35756 2632 35812
rect 2688 35756 2726 35812
rect 2782 35756 2820 35812
rect 2876 35756 2914 35812
rect 2970 35756 3008 35812
rect 3064 35758 3109 35812
rect 3165 35758 3193 35814
rect 3249 35758 3277 35814
rect 3333 35758 3360 35814
rect 3416 35758 3443 35814
rect 3499 35758 3526 35814
rect 3582 35758 3609 35814
rect 3665 35758 3692 35814
rect 3748 35758 3775 35814
rect 3831 35758 3858 35814
rect 3914 35758 3941 35814
rect 3997 35758 4024 35814
rect 4080 35758 4107 35814
rect 4163 35758 4190 35814
rect 4246 35758 4273 35814
rect 4329 35758 4356 35814
rect 4412 35758 4439 35814
rect 4495 35758 4522 35814
rect 4578 35758 4605 35814
rect 4661 35758 4688 35814
rect 4744 35758 4771 35814
rect 4827 35758 4854 35814
rect 4910 35758 4937 35814
rect 4993 35758 5002 35814
rect 3064 35756 5002 35758
rect 2525 35734 5002 35756
rect 2525 35732 3109 35734
rect 2525 35676 2538 35732
rect 2594 35676 2632 35732
rect 2688 35676 2726 35732
rect 2782 35676 2820 35732
rect 2876 35676 2914 35732
rect 2970 35676 3008 35732
rect 3064 35678 3109 35732
rect 3165 35678 3193 35734
rect 3249 35678 3277 35734
rect 3333 35678 3360 35734
rect 3416 35678 3443 35734
rect 3499 35678 3526 35734
rect 3582 35678 3609 35734
rect 3665 35678 3692 35734
rect 3748 35678 3775 35734
rect 3831 35678 3858 35734
rect 3914 35678 3941 35734
rect 3997 35678 4024 35734
rect 4080 35678 4107 35734
rect 4163 35678 4190 35734
rect 4246 35678 4273 35734
rect 4329 35678 4356 35734
rect 4412 35678 4439 35734
rect 4495 35678 4522 35734
rect 4578 35678 4605 35734
rect 4661 35678 4688 35734
rect 4744 35678 4771 35734
rect 4827 35678 4854 35734
rect 4910 35678 4937 35734
rect 4993 35678 5002 35734
rect 3064 35676 5002 35678
rect 2525 35654 5002 35676
rect 2525 35652 3109 35654
rect 2525 35596 2538 35652
rect 2594 35596 2632 35652
rect 2688 35596 2726 35652
rect 2782 35596 2820 35652
rect 2876 35596 2914 35652
rect 2970 35596 3008 35652
rect 3064 35598 3109 35652
rect 3165 35598 3193 35654
rect 3249 35598 3277 35654
rect 3333 35598 3360 35654
rect 3416 35598 3443 35654
rect 3499 35598 3526 35654
rect 3582 35598 3609 35654
rect 3665 35598 3692 35654
rect 3748 35598 3775 35654
rect 3831 35598 3858 35654
rect 3914 35598 3941 35654
rect 3997 35598 4024 35654
rect 4080 35598 4107 35654
rect 4163 35598 4190 35654
rect 4246 35598 4273 35654
rect 4329 35598 4356 35654
rect 4412 35598 4439 35654
rect 4495 35598 4522 35654
rect 4578 35598 4605 35654
rect 4661 35598 4688 35654
rect 4744 35598 4771 35654
rect 4827 35598 4854 35654
rect 4910 35598 4937 35654
rect 4993 35598 5002 35654
rect 3064 35596 5002 35598
rect 2525 35574 5002 35596
rect 2525 35572 3109 35574
rect 2525 35516 2538 35572
rect 2594 35516 2632 35572
rect 2688 35516 2726 35572
rect 2782 35516 2820 35572
rect 2876 35516 2914 35572
rect 2970 35516 3008 35572
rect 3064 35518 3109 35572
rect 3165 35518 3193 35574
rect 3249 35518 3277 35574
rect 3333 35518 3360 35574
rect 3416 35518 3443 35574
rect 3499 35518 3526 35574
rect 3582 35518 3609 35574
rect 3665 35518 3692 35574
rect 3748 35518 3775 35574
rect 3831 35518 3858 35574
rect 3914 35518 3941 35574
rect 3997 35518 4024 35574
rect 4080 35518 4107 35574
rect 4163 35518 4190 35574
rect 4246 35518 4273 35574
rect 4329 35518 4356 35574
rect 4412 35518 4439 35574
rect 4495 35518 4522 35574
rect 4578 35518 4605 35574
rect 4661 35518 4688 35574
rect 4744 35518 4771 35574
rect 4827 35518 4854 35574
rect 4910 35518 4937 35574
rect 4993 35518 5002 35574
rect 3064 35516 5002 35518
rect 2525 35494 5002 35516
rect 2525 35491 3109 35494
rect 2525 35435 2538 35491
rect 2594 35435 2632 35491
rect 2688 35435 2726 35491
rect 2782 35435 2820 35491
rect 2876 35435 2914 35491
rect 2970 35435 3008 35491
rect 3064 35438 3109 35491
rect 3165 35438 3193 35494
rect 3249 35438 3277 35494
rect 3333 35438 3360 35494
rect 3416 35438 3443 35494
rect 3499 35438 3526 35494
rect 3582 35438 3609 35494
rect 3665 35438 3692 35494
rect 3748 35438 3775 35494
rect 3831 35438 3858 35494
rect 3914 35438 3941 35494
rect 3997 35438 4024 35494
rect 4080 35438 4107 35494
rect 4163 35438 4190 35494
rect 4246 35438 4273 35494
rect 4329 35438 4356 35494
rect 4412 35438 4439 35494
rect 4495 35438 4522 35494
rect 4578 35438 4605 35494
rect 4661 35438 4688 35494
rect 4744 35438 4771 35494
rect 4827 35438 4854 35494
rect 4910 35438 4937 35494
rect 4993 35438 5002 35494
rect 3064 35435 5002 35438
rect 2525 35414 5002 35435
rect 2525 35410 3109 35414
rect 2525 35354 2538 35410
rect 2594 35354 2632 35410
rect 2688 35354 2726 35410
rect 2782 35354 2820 35410
rect 2876 35354 2914 35410
rect 2970 35354 3008 35410
rect 3064 35358 3109 35410
rect 3165 35358 3193 35414
rect 3249 35358 3277 35414
rect 3333 35358 3360 35414
rect 3416 35358 3443 35414
rect 3499 35358 3526 35414
rect 3582 35358 3609 35414
rect 3665 35358 3692 35414
rect 3748 35358 3775 35414
rect 3831 35358 3858 35414
rect 3914 35358 3941 35414
rect 3997 35358 4024 35414
rect 4080 35358 4107 35414
rect 4163 35358 4190 35414
rect 4246 35358 4273 35414
rect 4329 35358 4356 35414
rect 4412 35358 4439 35414
rect 4495 35358 4522 35414
rect 4578 35358 4605 35414
rect 4661 35358 4688 35414
rect 4744 35358 4771 35414
rect 4827 35358 4854 35414
rect 4910 35358 4937 35414
rect 4993 35358 5002 35414
rect 3064 35354 5002 35358
rect 2525 35334 5002 35354
rect 2525 35329 3109 35334
rect 2525 35273 2538 35329
rect 2594 35273 2632 35329
rect 2688 35273 2726 35329
rect 2782 35273 2820 35329
rect 2876 35273 2914 35329
rect 2970 35273 3008 35329
rect 3064 35278 3109 35329
rect 3165 35278 3193 35334
rect 3249 35278 3277 35334
rect 3333 35278 3360 35334
rect 3416 35278 3443 35334
rect 3499 35278 3526 35334
rect 3582 35278 3609 35334
rect 3665 35278 3692 35334
rect 3748 35278 3775 35334
rect 3831 35278 3858 35334
rect 3914 35278 3941 35334
rect 3997 35278 4024 35334
rect 4080 35278 4107 35334
rect 4163 35278 4190 35334
rect 4246 35278 4273 35334
rect 4329 35278 4356 35334
rect 4412 35278 4439 35334
rect 4495 35278 4522 35334
rect 4578 35278 4605 35334
rect 4661 35278 4688 35334
rect 4744 35278 4771 35334
rect 4827 35278 4854 35334
rect 4910 35278 4937 35334
rect 4993 35278 5002 35334
rect 3064 35273 5002 35278
rect 2525 35254 5002 35273
rect 2525 35248 3109 35254
rect 2525 35192 2538 35248
rect 2594 35192 2632 35248
rect 2688 35192 2726 35248
rect 2782 35192 2820 35248
rect 2876 35192 2914 35248
rect 2970 35192 3008 35248
rect 3064 35198 3109 35248
rect 3165 35198 3193 35254
rect 3249 35198 3277 35254
rect 3333 35198 3360 35254
rect 3416 35198 3443 35254
rect 3499 35198 3526 35254
rect 3582 35198 3609 35254
rect 3665 35198 3692 35254
rect 3748 35198 3775 35254
rect 3831 35198 3858 35254
rect 3914 35198 3941 35254
rect 3997 35198 4024 35254
rect 4080 35198 4107 35254
rect 4163 35198 4190 35254
rect 4246 35198 4273 35254
rect 4329 35198 4356 35254
rect 4412 35198 4439 35254
rect 4495 35198 4522 35254
rect 4578 35198 4605 35254
rect 4661 35198 4688 35254
rect 4744 35198 4771 35254
rect 4827 35198 4854 35254
rect 4910 35198 4937 35254
rect 4993 35198 5002 35254
rect 3064 35192 5002 35198
rect 2525 35179 5002 35192
tri 2525 35174 2530 35179 ne
rect 2530 35174 5002 35179
tri 2530 35150 2554 35174 ne
rect 2554 35150 3109 35174
tri 2554 35139 2565 35150 ne
rect 2565 35139 2821 35150
tri 2565 35083 2621 35139 ne
rect 2621 35083 2675 35139
rect 2731 35094 2821 35139
rect 2877 35094 2914 35150
rect 2970 35094 3006 35150
rect 3062 35118 3109 35150
rect 3165 35118 3193 35174
rect 3249 35118 3277 35174
rect 3333 35118 3360 35174
rect 3416 35118 3443 35174
rect 3499 35118 3526 35174
rect 3582 35118 3609 35174
rect 3665 35118 3692 35174
rect 3748 35118 3775 35174
rect 3831 35118 3858 35174
rect 3914 35118 3941 35174
rect 3997 35118 4024 35174
rect 4080 35118 4107 35174
rect 4163 35118 4190 35174
rect 4246 35118 4273 35174
rect 4329 35118 4356 35174
rect 4412 35118 4439 35174
rect 4495 35118 4522 35174
rect 4578 35118 4605 35174
rect 4661 35118 4688 35174
rect 4744 35118 4771 35174
rect 4827 35118 4854 35174
rect 4910 35118 4937 35174
rect 4993 35118 5002 35174
rect 3062 35094 5002 35118
rect 2731 35083 3109 35094
tri 2621 35070 2634 35083 ne
rect 2634 35070 3109 35083
tri 2634 35058 2646 35070 ne
rect 2646 35058 3109 35070
tri 2646 35052 2652 35058 ne
rect 2652 35052 2821 35058
tri 2652 35002 2702 35052 ne
rect 2702 35002 2821 35052
rect 2877 35002 2914 35058
rect 2970 35002 3006 35058
rect 3062 35038 3109 35058
rect 3165 35038 3193 35094
rect 3249 35038 3277 35094
rect 3333 35038 3360 35094
rect 3416 35038 3443 35094
rect 3499 35038 3526 35094
rect 3582 35038 3609 35094
rect 3665 35038 3692 35094
rect 3748 35038 3775 35094
rect 3831 35038 3858 35094
rect 3914 35038 3941 35094
rect 3997 35038 4024 35094
rect 4080 35038 4107 35094
rect 4163 35038 4190 35094
rect 4246 35038 4273 35094
rect 4329 35038 4356 35094
rect 4412 35038 4439 35094
rect 4495 35038 4522 35094
rect 4578 35038 4605 35094
rect 4661 35038 4688 35094
rect 4744 35038 4771 35094
rect 4827 35038 4854 35094
rect 4910 35038 4937 35094
rect 4993 35038 5002 35094
rect 3062 35014 5002 35038
rect 3062 35002 3109 35014
tri 2702 34966 2738 35002 ne
rect 2738 34966 3109 35002
tri 2738 34910 2794 34966 ne
rect 2794 34910 2821 34966
rect 2877 34910 2914 34966
rect 2970 34910 3006 34966
rect 3062 34958 3109 34966
rect 3165 34958 3193 35014
rect 3249 34958 3277 35014
rect 3333 34958 3360 35014
rect 3416 34958 3443 35014
rect 3499 34958 3526 35014
rect 3582 34958 3609 35014
rect 3665 34958 3692 35014
rect 3748 34958 3775 35014
rect 3831 34958 3858 35014
rect 3914 34958 3941 35014
rect 3997 34958 4024 35014
rect 4080 34958 4107 35014
rect 4163 34958 4190 35014
rect 4246 34958 4273 35014
rect 4329 34958 4356 35014
rect 4412 34958 4439 35014
rect 4495 34958 4522 35014
rect 4578 34958 4605 35014
rect 4661 34958 4688 35014
rect 4744 34958 4771 35014
rect 4827 34958 4854 35014
rect 4910 34958 4937 35014
rect 4993 34958 5002 35014
rect 3062 34934 5002 34958
rect 3062 34910 3109 34934
tri 2794 34904 2800 34910 ne
rect 2800 34904 3109 34910
tri 2800 34882 2822 34904 ne
rect 2822 34882 3109 34904
tri 2822 34878 2826 34882 ne
rect 2826 34878 3109 34882
rect 3165 34878 3193 34934
rect 3249 34878 3277 34934
rect 3333 34878 3360 34934
rect 3416 34878 3443 34934
rect 3499 34878 3526 34934
rect 3582 34878 3609 34934
rect 3665 34878 3692 34934
rect 3748 34878 3775 34934
rect 3831 34878 3858 34934
rect 3914 34878 3941 34934
rect 3997 34878 4024 34934
rect 4080 34878 4107 34934
rect 4163 34878 4190 34934
rect 4246 34878 4273 34934
rect 4329 34878 4356 34934
rect 4412 34878 4439 34934
rect 4495 34878 4522 34934
rect 4578 34878 4605 34934
rect 4661 34878 4688 34934
rect 4744 34878 4771 34934
rect 4827 34878 4854 34934
rect 4910 34878 4937 34934
rect 4993 34878 5002 34934
tri 2826 34867 2837 34878 ne
rect 2837 34867 5002 34878
tri 2837 34854 2850 34867 ne
rect 2850 34854 5002 34867
tri 2850 34851 2853 34854 ne
rect 2853 34851 3109 34854
tri 2853 34795 2909 34851 ne
rect 2909 34795 2963 34851
rect 3019 34798 3109 34851
rect 3165 34798 3193 34854
rect 3249 34798 3277 34854
rect 3333 34798 3360 34854
rect 3416 34798 3443 34854
rect 3499 34798 3526 34854
rect 3582 34798 3609 34854
rect 3665 34798 3692 34854
rect 3748 34798 3775 34854
rect 3831 34798 3858 34854
rect 3914 34798 3941 34854
rect 3997 34798 4024 34854
rect 4080 34798 4107 34854
rect 4163 34798 4190 34854
rect 4246 34798 4273 34854
rect 4329 34798 4356 34854
rect 4412 34798 4439 34854
rect 4495 34798 4522 34854
rect 4578 34798 4605 34854
rect 4661 34798 4688 34854
rect 4744 34798 4771 34854
rect 4827 34798 4854 34854
rect 4910 34798 4937 34854
rect 4993 34798 5002 34854
rect 3019 34795 5002 34798
tri 2909 34779 2925 34795 ne
rect 2925 34779 5002 34795
tri 2925 34774 2930 34779 ne
rect 2930 34774 5002 34779
tri 2930 34764 2940 34774 ne
rect 2940 34764 3109 34774
tri 2940 34718 2986 34764 ne
rect 2986 34718 3109 34764
rect 3165 34718 3193 34774
rect 3249 34718 3277 34774
rect 3333 34718 3360 34774
rect 3416 34718 3443 34774
rect 3499 34718 3526 34774
rect 3582 34718 3609 34774
rect 3665 34718 3692 34774
rect 3748 34718 3775 34774
rect 3831 34718 3858 34774
rect 3914 34718 3941 34774
rect 3997 34718 4024 34774
rect 4080 34718 4107 34774
rect 4163 34718 4190 34774
rect 4246 34718 4273 34774
rect 4329 34718 4356 34774
rect 4412 34718 4439 34774
rect 4495 34718 4522 34774
rect 4578 34718 4605 34774
rect 4661 34718 4688 34774
rect 4744 34718 4771 34774
rect 4827 34718 4854 34774
rect 4910 34718 4937 34774
rect 4993 34718 5002 34774
tri 2986 34695 3009 34718 ne
rect 3009 34695 5002 34718
tri 3009 34694 3010 34695 ne
rect 3010 34694 5002 34695
tri 3010 34638 3066 34694 ne
rect 3066 34638 3109 34694
rect 3165 34638 3193 34694
rect 3249 34638 3277 34694
rect 3333 34638 3360 34694
rect 3416 34638 3443 34694
rect 3499 34638 3526 34694
rect 3582 34638 3609 34694
rect 3665 34638 3692 34694
rect 3748 34638 3775 34694
rect 3831 34638 3858 34694
rect 3914 34638 3941 34694
rect 3997 34638 4024 34694
rect 4080 34638 4107 34694
rect 4163 34638 4190 34694
rect 4246 34638 4273 34694
rect 4329 34638 4356 34694
rect 4412 34638 4439 34694
rect 4495 34638 4522 34694
rect 4578 34638 4605 34694
rect 4661 34638 4688 34694
rect 4744 34638 4771 34694
rect 4827 34638 4854 34694
rect 4910 34638 4937 34694
rect 4993 34638 5002 34694
tri 3066 34614 3090 34638 ne
rect 3090 34614 5002 34638
tri 3090 34604 3100 34614 ne
rect 3100 34558 3109 34614
rect 3165 34558 3193 34614
rect 3249 34558 3277 34614
rect 3333 34558 3360 34614
rect 3416 34558 3443 34614
rect 3499 34558 3526 34614
rect 3582 34558 3609 34614
rect 3665 34558 3692 34614
rect 3748 34558 3775 34614
rect 3831 34558 3858 34614
rect 3914 34558 3941 34614
rect 3997 34558 4024 34614
rect 4080 34558 4107 34614
rect 4163 34558 4190 34614
rect 4246 34558 4273 34614
rect 4329 34558 4356 34614
rect 4412 34558 4439 34614
rect 4495 34558 4522 34614
rect 4578 34558 4605 34614
rect 4661 34558 4688 34614
rect 4744 34558 4771 34614
rect 4827 34558 4854 34614
rect 4910 34558 4937 34614
rect 4993 34558 5002 34614
rect 3100 34528 5002 34558
rect 3100 34229 4703 34528
tri 4703 34229 5002 34528 nw
rect 5186 39009 7364 39015
rect 5186 38953 5195 39009
rect 5251 38953 5276 39009
rect 5332 38953 5357 39009
rect 5413 38953 5438 39009
rect 5494 38953 5519 39009
rect 5575 38953 5600 39009
rect 5656 38953 5681 39009
rect 5737 38953 5762 39009
rect 5818 38953 5843 39009
rect 5899 38953 5924 39009
rect 5980 38953 6005 39009
rect 6061 38953 6086 39009
rect 6142 38953 6167 39009
rect 6223 38953 6248 39009
rect 6304 38953 6329 39009
rect 6385 38953 6410 39009
rect 6466 38953 6491 39009
rect 6547 38953 6572 39009
rect 6628 38953 6653 39009
rect 6709 38953 6734 39009
rect 6790 38953 6815 39009
rect 6871 38953 6896 39009
rect 6952 38953 6977 39009
rect 7033 38953 7058 39009
rect 7114 38953 7139 39009
rect 7195 38953 7221 39009
rect 7277 38953 7303 39009
rect 7359 38953 7364 39009
rect 5186 38925 7364 38953
rect 5186 38869 5195 38925
rect 5251 38869 5276 38925
rect 5332 38869 5357 38925
rect 5413 38869 5438 38925
rect 5494 38869 5519 38925
rect 5575 38869 5600 38925
rect 5656 38869 5681 38925
rect 5737 38869 5762 38925
rect 5818 38869 5843 38925
rect 5899 38869 5924 38925
rect 5980 38869 6005 38925
rect 6061 38869 6086 38925
rect 6142 38869 6167 38925
rect 6223 38869 6248 38925
rect 6304 38869 6329 38925
rect 6385 38869 6410 38925
rect 6466 38869 6491 38925
rect 6547 38869 6572 38925
rect 6628 38869 6653 38925
rect 6709 38869 6734 38925
rect 6790 38869 6815 38925
rect 6871 38869 6896 38925
rect 6952 38869 6977 38925
rect 7033 38869 7058 38925
rect 7114 38869 7139 38925
rect 7195 38869 7221 38925
rect 7277 38869 7303 38925
rect 7359 38869 7364 38925
rect 5186 38841 7364 38869
rect 5186 38785 5195 38841
rect 5251 38785 5276 38841
rect 5332 38785 5357 38841
rect 5413 38785 5438 38841
rect 5494 38785 5519 38841
rect 5575 38785 5600 38841
rect 5656 38785 5681 38841
rect 5737 38785 5762 38841
rect 5818 38785 5843 38841
rect 5899 38785 5924 38841
rect 5980 38785 6005 38841
rect 6061 38785 6086 38841
rect 6142 38785 6167 38841
rect 6223 38785 6248 38841
rect 6304 38785 6329 38841
rect 6385 38785 6410 38841
rect 6466 38785 6491 38841
rect 6547 38785 6572 38841
rect 6628 38785 6653 38841
rect 6709 38785 6734 38841
rect 6790 38785 6815 38841
rect 6871 38785 6896 38841
rect 6952 38785 6977 38841
rect 7033 38785 7058 38841
rect 7114 38785 7139 38841
rect 7195 38785 7221 38841
rect 7277 38785 7303 38841
rect 7359 38785 7364 38841
rect 5186 38757 7364 38785
rect 5186 38701 5195 38757
rect 5251 38701 5276 38757
rect 5332 38701 5357 38757
rect 5413 38701 5438 38757
rect 5494 38701 5519 38757
rect 5575 38701 5600 38757
rect 5656 38701 5681 38757
rect 5737 38701 5762 38757
rect 5818 38701 5843 38757
rect 5899 38701 5924 38757
rect 5980 38701 6005 38757
rect 6061 38701 6086 38757
rect 6142 38701 6167 38757
rect 6223 38701 6248 38757
rect 6304 38701 6329 38757
rect 6385 38701 6410 38757
rect 6466 38701 6491 38757
rect 6547 38701 6572 38757
rect 6628 38701 6653 38757
rect 6709 38701 6734 38757
rect 6790 38701 6815 38757
rect 6871 38701 6896 38757
rect 6952 38701 6977 38757
rect 7033 38701 7058 38757
rect 7114 38701 7139 38757
rect 7195 38701 7221 38757
rect 7277 38701 7303 38757
rect 7359 38701 7364 38757
rect 5186 38673 7364 38701
rect 5186 38617 5195 38673
rect 5251 38617 5276 38673
rect 5332 38617 5357 38673
rect 5413 38617 5438 38673
rect 5494 38617 5519 38673
rect 5575 38617 5600 38673
rect 5656 38617 5681 38673
rect 5737 38617 5762 38673
rect 5818 38617 5843 38673
rect 5899 38617 5924 38673
rect 5980 38617 6005 38673
rect 6061 38617 6086 38673
rect 6142 38617 6167 38673
rect 6223 38617 6248 38673
rect 6304 38617 6329 38673
rect 6385 38617 6410 38673
rect 6466 38617 6491 38673
rect 6547 38617 6572 38673
rect 6628 38617 6653 38673
rect 6709 38617 6734 38673
rect 6790 38617 6815 38673
rect 6871 38617 6896 38673
rect 6952 38617 6977 38673
rect 7033 38617 7058 38673
rect 7114 38617 7139 38673
rect 7195 38617 7221 38673
rect 7277 38617 7303 38673
rect 7359 38617 7364 38673
rect 5186 38589 7364 38617
rect 5186 38533 5195 38589
rect 5251 38533 5276 38589
rect 5332 38533 5357 38589
rect 5413 38533 5438 38589
rect 5494 38533 5519 38589
rect 5575 38533 5600 38589
rect 5656 38533 5681 38589
rect 5737 38533 5762 38589
rect 5818 38533 5843 38589
rect 5899 38533 5924 38589
rect 5980 38533 6005 38589
rect 6061 38533 6086 38589
rect 6142 38533 6167 38589
rect 6223 38533 6248 38589
rect 6304 38533 6329 38589
rect 6385 38533 6410 38589
rect 6466 38533 6491 38589
rect 6547 38533 6572 38589
rect 6628 38533 6653 38589
rect 6709 38533 6734 38589
rect 6790 38533 6815 38589
rect 6871 38533 6896 38589
rect 6952 38533 6977 38589
rect 7033 38533 7058 38589
rect 7114 38533 7139 38589
rect 7195 38533 7221 38589
rect 7277 38533 7303 38589
rect 7359 38533 7364 38589
rect 5186 38505 7364 38533
rect 5186 38449 5195 38505
rect 5251 38449 5276 38505
rect 5332 38449 5357 38505
rect 5413 38449 5438 38505
rect 5494 38449 5519 38505
rect 5575 38449 5600 38505
rect 5656 38449 5681 38505
rect 5737 38449 5762 38505
rect 5818 38449 5843 38505
rect 5899 38449 5924 38505
rect 5980 38449 6005 38505
rect 6061 38449 6086 38505
rect 6142 38449 6167 38505
rect 6223 38449 6248 38505
rect 6304 38449 6329 38505
rect 6385 38449 6410 38505
rect 6466 38449 6491 38505
rect 6547 38449 6572 38505
rect 6628 38449 6653 38505
rect 6709 38449 6734 38505
rect 6790 38449 6815 38505
rect 6871 38449 6896 38505
rect 6952 38449 6977 38505
rect 7033 38449 7058 38505
rect 7114 38449 7139 38505
rect 7195 38449 7221 38505
rect 7277 38449 7303 38505
rect 7359 38449 7364 38505
rect 5186 38421 7364 38449
rect 5186 38365 5195 38421
rect 5251 38365 5276 38421
rect 5332 38365 5357 38421
rect 5413 38365 5438 38421
rect 5494 38365 5519 38421
rect 5575 38365 5600 38421
rect 5656 38365 5681 38421
rect 5737 38365 5762 38421
rect 5818 38365 5843 38421
rect 5899 38365 5924 38421
rect 5980 38365 6005 38421
rect 6061 38365 6086 38421
rect 6142 38365 6167 38421
rect 6223 38365 6248 38421
rect 6304 38365 6329 38421
rect 6385 38365 6410 38421
rect 6466 38365 6491 38421
rect 6547 38365 6572 38421
rect 6628 38365 6653 38421
rect 6709 38365 6734 38421
rect 6790 38365 6815 38421
rect 6871 38365 6896 38421
rect 6952 38365 6977 38421
rect 7033 38365 7058 38421
rect 7114 38365 7139 38421
rect 7195 38365 7221 38421
rect 7277 38365 7303 38421
rect 7359 38365 7364 38421
rect 5186 38337 7364 38365
rect 5186 38281 5195 38337
rect 5251 38281 5276 38337
rect 5332 38281 5357 38337
rect 5413 38281 5438 38337
rect 5494 38281 5519 38337
rect 5575 38281 5600 38337
rect 5656 38281 5681 38337
rect 5737 38281 5762 38337
rect 5818 38281 5843 38337
rect 5899 38281 5924 38337
rect 5980 38281 6005 38337
rect 6061 38281 6086 38337
rect 6142 38281 6167 38337
rect 6223 38281 6248 38337
rect 6304 38281 6329 38337
rect 6385 38281 6410 38337
rect 6466 38281 6491 38337
rect 6547 38281 6572 38337
rect 6628 38281 6653 38337
rect 6709 38281 6734 38337
rect 6790 38281 6815 38337
rect 6871 38281 6896 38337
rect 6952 38281 6977 38337
rect 7033 38281 7058 38337
rect 7114 38281 7139 38337
rect 7195 38281 7221 38337
rect 7277 38281 7303 38337
rect 7359 38281 7364 38337
rect 5186 38253 7364 38281
rect 5186 38197 5195 38253
rect 5251 38197 5276 38253
rect 5332 38197 5357 38253
rect 5413 38197 5438 38253
rect 5494 38197 5519 38253
rect 5575 38197 5600 38253
rect 5656 38197 5681 38253
rect 5737 38197 5762 38253
rect 5818 38197 5843 38253
rect 5899 38197 5924 38253
rect 5980 38197 6005 38253
rect 6061 38197 6086 38253
rect 6142 38197 6167 38253
rect 6223 38197 6248 38253
rect 6304 38197 6329 38253
rect 6385 38197 6410 38253
rect 6466 38197 6491 38253
rect 6547 38197 6572 38253
rect 6628 38197 6653 38253
rect 6709 38197 6734 38253
rect 6790 38197 6815 38253
rect 6871 38197 6896 38253
rect 6952 38197 6977 38253
rect 7033 38197 7058 38253
rect 7114 38197 7139 38253
rect 7195 38197 7221 38253
rect 7277 38197 7303 38253
rect 7359 38197 7364 38253
rect 5186 38169 7364 38197
rect 5186 38113 5195 38169
rect 5251 38113 5276 38169
rect 5332 38113 5357 38169
rect 5413 38113 5438 38169
rect 5494 38113 5519 38169
rect 5575 38113 5600 38169
rect 5656 38113 5681 38169
rect 5737 38113 5762 38169
rect 5818 38113 5843 38169
rect 5899 38113 5924 38169
rect 5980 38113 6005 38169
rect 6061 38113 6086 38169
rect 6142 38113 6167 38169
rect 6223 38113 6248 38169
rect 6304 38113 6329 38169
rect 6385 38113 6410 38169
rect 6466 38113 6491 38169
rect 6547 38113 6572 38169
rect 6628 38113 6653 38169
rect 6709 38113 6734 38169
rect 6790 38113 6815 38169
rect 6871 38113 6896 38169
rect 6952 38113 6977 38169
rect 7033 38113 7058 38169
rect 7114 38113 7139 38169
rect 7195 38113 7221 38169
rect 7277 38113 7303 38169
rect 7359 38113 7364 38169
rect 5186 36294 7364 38113
rect 5186 36238 5195 36294
rect 5251 36238 5277 36294
rect 5333 36238 5359 36294
rect 5415 36238 5441 36294
rect 5497 36238 5523 36294
rect 5579 36238 5605 36294
rect 5661 36238 5687 36294
rect 5743 36238 5769 36294
rect 5825 36238 5851 36294
rect 5907 36238 5933 36294
rect 5989 36238 6015 36294
rect 6071 36238 6097 36294
rect 6153 36238 6179 36294
rect 6235 36238 6261 36294
rect 6317 36238 6343 36294
rect 6399 36238 6425 36294
rect 6481 36238 6507 36294
rect 6563 36238 6589 36294
rect 6645 36238 6671 36294
rect 6727 36238 6753 36294
rect 6809 36278 7364 36294
rect 6809 36238 6853 36278
rect 5186 36222 6853 36238
rect 6909 36222 6941 36278
rect 6997 36222 7029 36278
rect 7085 36222 7117 36278
rect 7173 36222 7205 36278
rect 7261 36222 7293 36278
rect 7349 36222 7364 36278
rect 5186 36214 7364 36222
rect 5186 36158 5195 36214
rect 5251 36158 5277 36214
rect 5333 36158 5359 36214
rect 5415 36158 5441 36214
rect 5497 36158 5523 36214
rect 5579 36158 5605 36214
rect 5661 36158 5687 36214
rect 5743 36158 5769 36214
rect 5825 36158 5851 36214
rect 5907 36158 5933 36214
rect 5989 36158 6015 36214
rect 6071 36158 6097 36214
rect 6153 36158 6179 36214
rect 6235 36158 6261 36214
rect 6317 36158 6343 36214
rect 6399 36158 6425 36214
rect 6481 36158 6507 36214
rect 6563 36158 6589 36214
rect 6645 36158 6671 36214
rect 6727 36158 6753 36214
rect 6809 36196 7364 36214
rect 6809 36158 6853 36196
rect 5186 36140 6853 36158
rect 6909 36140 6941 36196
rect 6997 36140 7029 36196
rect 7085 36140 7117 36196
rect 7173 36140 7205 36196
rect 7261 36140 7293 36196
rect 7349 36140 7364 36196
rect 5186 36134 7364 36140
rect 5186 36078 5195 36134
rect 5251 36078 5277 36134
rect 5333 36078 5359 36134
rect 5415 36078 5441 36134
rect 5497 36078 5523 36134
rect 5579 36078 5605 36134
rect 5661 36078 5687 36134
rect 5743 36078 5769 36134
rect 5825 36078 5851 36134
rect 5907 36078 5933 36134
rect 5989 36078 6015 36134
rect 6071 36078 6097 36134
rect 6153 36078 6179 36134
rect 6235 36078 6261 36134
rect 6317 36078 6343 36134
rect 6399 36078 6425 36134
rect 6481 36078 6507 36134
rect 6563 36078 6589 36134
rect 6645 36078 6671 36134
rect 6727 36078 6753 36134
rect 6809 36114 7364 36134
rect 6809 36078 6853 36114
rect 5186 36058 6853 36078
rect 6909 36058 6941 36114
rect 6997 36058 7029 36114
rect 7085 36058 7117 36114
rect 7173 36058 7205 36114
rect 7261 36058 7293 36114
rect 7349 36058 7364 36114
rect 5186 36054 7364 36058
rect 5186 35998 5195 36054
rect 5251 35998 5277 36054
rect 5333 35998 5359 36054
rect 5415 35998 5441 36054
rect 5497 35998 5523 36054
rect 5579 35998 5605 36054
rect 5661 35998 5687 36054
rect 5743 35998 5769 36054
rect 5825 35998 5851 36054
rect 5907 35998 5933 36054
rect 5989 35998 6015 36054
rect 6071 35998 6097 36054
rect 6153 35998 6179 36054
rect 6235 35998 6261 36054
rect 6317 35998 6343 36054
rect 6399 35998 6425 36054
rect 6481 35998 6507 36054
rect 6563 35998 6589 36054
rect 6645 35998 6671 36054
rect 6727 35998 6753 36054
rect 6809 36032 7364 36054
rect 6809 35998 6853 36032
rect 5186 35976 6853 35998
rect 6909 35976 6941 36032
rect 6997 35976 7029 36032
rect 7085 35976 7117 36032
rect 7173 35976 7205 36032
rect 7261 35976 7293 36032
rect 7349 35976 7364 36032
rect 5186 35974 7364 35976
rect 5186 35918 5195 35974
rect 5251 35918 5277 35974
rect 5333 35918 5359 35974
rect 5415 35918 5441 35974
rect 5497 35918 5523 35974
rect 5579 35918 5605 35974
rect 5661 35918 5687 35974
rect 5743 35918 5769 35974
rect 5825 35918 5851 35974
rect 5907 35918 5933 35974
rect 5989 35918 6015 35974
rect 6071 35918 6097 35974
rect 6153 35918 6179 35974
rect 6235 35918 6261 35974
rect 6317 35918 6343 35974
rect 6399 35918 6425 35974
rect 6481 35918 6507 35974
rect 6563 35918 6589 35974
rect 6645 35918 6671 35974
rect 6727 35918 6753 35974
rect 6809 35950 7364 35974
rect 6809 35918 6853 35950
rect 5186 35894 6853 35918
rect 6909 35894 6941 35950
rect 6997 35894 7029 35950
rect 7085 35894 7117 35950
rect 7173 35894 7205 35950
rect 7261 35894 7293 35950
rect 7349 35894 7364 35950
rect 5186 35838 5195 35894
rect 5251 35838 5277 35894
rect 5333 35838 5359 35894
rect 5415 35838 5441 35894
rect 5497 35838 5523 35894
rect 5579 35838 5605 35894
rect 5661 35838 5687 35894
rect 5743 35838 5769 35894
rect 5825 35838 5851 35894
rect 5907 35838 5933 35894
rect 5989 35838 6015 35894
rect 6071 35838 6097 35894
rect 6153 35838 6179 35894
rect 6235 35838 6261 35894
rect 6317 35838 6343 35894
rect 6399 35838 6425 35894
rect 6481 35838 6507 35894
rect 6563 35838 6589 35894
rect 6645 35838 6671 35894
rect 6727 35838 6753 35894
rect 6809 35868 7364 35894
rect 6809 35838 6853 35868
rect 5186 35814 6853 35838
rect 5186 35758 5195 35814
rect 5251 35758 5277 35814
rect 5333 35758 5359 35814
rect 5415 35758 5441 35814
rect 5497 35758 5523 35814
rect 5579 35758 5605 35814
rect 5661 35758 5687 35814
rect 5743 35758 5769 35814
rect 5825 35758 5851 35814
rect 5907 35758 5933 35814
rect 5989 35758 6015 35814
rect 6071 35758 6097 35814
rect 6153 35758 6179 35814
rect 6235 35758 6261 35814
rect 6317 35758 6343 35814
rect 6399 35758 6425 35814
rect 6481 35758 6507 35814
rect 6563 35758 6589 35814
rect 6645 35758 6671 35814
rect 6727 35758 6753 35814
rect 6809 35812 6853 35814
rect 6909 35812 6941 35868
rect 6997 35812 7029 35868
rect 7085 35812 7117 35868
rect 7173 35812 7205 35868
rect 7261 35812 7293 35868
rect 7349 35812 7364 35868
rect 6809 35786 7364 35812
rect 6809 35758 6853 35786
rect 5186 35734 6853 35758
rect 5186 35678 5195 35734
rect 5251 35678 5277 35734
rect 5333 35678 5359 35734
rect 5415 35678 5441 35734
rect 5497 35678 5523 35734
rect 5579 35678 5605 35734
rect 5661 35678 5687 35734
rect 5743 35678 5769 35734
rect 5825 35678 5851 35734
rect 5907 35678 5933 35734
rect 5989 35678 6015 35734
rect 6071 35678 6097 35734
rect 6153 35678 6179 35734
rect 6235 35678 6261 35734
rect 6317 35678 6343 35734
rect 6399 35678 6425 35734
rect 6481 35678 6507 35734
rect 6563 35678 6589 35734
rect 6645 35678 6671 35734
rect 6727 35678 6753 35734
rect 6809 35730 6853 35734
rect 6909 35730 6941 35786
rect 6997 35730 7029 35786
rect 7085 35730 7117 35786
rect 7173 35730 7205 35786
rect 7261 35730 7293 35786
rect 7349 35730 7364 35786
rect 6809 35704 7364 35730
rect 6809 35678 6853 35704
rect 5186 35654 6853 35678
rect 5186 35598 5195 35654
rect 5251 35598 5277 35654
rect 5333 35598 5359 35654
rect 5415 35598 5441 35654
rect 5497 35598 5523 35654
rect 5579 35598 5605 35654
rect 5661 35598 5687 35654
rect 5743 35598 5769 35654
rect 5825 35598 5851 35654
rect 5907 35598 5933 35654
rect 5989 35598 6015 35654
rect 6071 35598 6097 35654
rect 6153 35598 6179 35654
rect 6235 35598 6261 35654
rect 6317 35598 6343 35654
rect 6399 35598 6425 35654
rect 6481 35598 6507 35654
rect 6563 35598 6589 35654
rect 6645 35598 6671 35654
rect 6727 35598 6753 35654
rect 6809 35648 6853 35654
rect 6909 35648 6941 35704
rect 6997 35648 7029 35704
rect 7085 35648 7117 35704
rect 7173 35648 7205 35704
rect 7261 35648 7293 35704
rect 7349 35648 7364 35704
rect 6809 35622 7364 35648
rect 6809 35598 6853 35622
rect 5186 35574 6853 35598
rect 5186 35518 5195 35574
rect 5251 35518 5277 35574
rect 5333 35518 5359 35574
rect 5415 35518 5441 35574
rect 5497 35518 5523 35574
rect 5579 35518 5605 35574
rect 5661 35518 5687 35574
rect 5743 35518 5769 35574
rect 5825 35518 5851 35574
rect 5907 35518 5933 35574
rect 5989 35518 6015 35574
rect 6071 35518 6097 35574
rect 6153 35518 6179 35574
rect 6235 35518 6261 35574
rect 6317 35518 6343 35574
rect 6399 35518 6425 35574
rect 6481 35518 6507 35574
rect 6563 35518 6589 35574
rect 6645 35518 6671 35574
rect 6727 35518 6753 35574
rect 6809 35566 6853 35574
rect 6909 35566 6941 35622
rect 6997 35566 7029 35622
rect 7085 35566 7117 35622
rect 7173 35566 7205 35622
rect 7261 35566 7293 35622
rect 7349 35566 7364 35622
rect 6809 35539 7364 35566
rect 6809 35518 6853 35539
rect 5186 35494 6853 35518
rect 5186 35438 5195 35494
rect 5251 35438 5277 35494
rect 5333 35438 5359 35494
rect 5415 35438 5441 35494
rect 5497 35438 5523 35494
rect 5579 35438 5605 35494
rect 5661 35438 5687 35494
rect 5743 35438 5769 35494
rect 5825 35438 5851 35494
rect 5907 35438 5933 35494
rect 5989 35438 6015 35494
rect 6071 35438 6097 35494
rect 6153 35438 6179 35494
rect 6235 35438 6261 35494
rect 6317 35438 6343 35494
rect 6399 35438 6425 35494
rect 6481 35438 6507 35494
rect 6563 35438 6589 35494
rect 6645 35438 6671 35494
rect 6727 35438 6753 35494
rect 6809 35483 6853 35494
rect 6909 35483 6941 35539
rect 6997 35483 7029 35539
rect 7085 35483 7117 35539
rect 7173 35483 7205 35539
rect 7261 35483 7293 35539
rect 7349 35483 7364 35539
rect 6809 35456 7364 35483
rect 6809 35438 6853 35456
rect 5186 35414 6853 35438
rect 5186 35358 5195 35414
rect 5251 35358 5277 35414
rect 5333 35358 5359 35414
rect 5415 35358 5441 35414
rect 5497 35358 5523 35414
rect 5579 35358 5605 35414
rect 5661 35358 5687 35414
rect 5743 35358 5769 35414
rect 5825 35358 5851 35414
rect 5907 35358 5933 35414
rect 5989 35358 6015 35414
rect 6071 35358 6097 35414
rect 6153 35358 6179 35414
rect 6235 35358 6261 35414
rect 6317 35358 6343 35414
rect 6399 35358 6425 35414
rect 6481 35358 6507 35414
rect 6563 35358 6589 35414
rect 6645 35358 6671 35414
rect 6727 35358 6753 35414
rect 6809 35400 6853 35414
rect 6909 35400 6941 35456
rect 6997 35400 7029 35456
rect 7085 35400 7117 35456
rect 7173 35400 7205 35456
rect 7261 35400 7293 35456
rect 7349 35400 7364 35456
rect 6809 35373 7364 35400
rect 6809 35358 6853 35373
rect 5186 35334 6853 35358
rect 5186 35278 5195 35334
rect 5251 35278 5277 35334
rect 5333 35278 5359 35334
rect 5415 35278 5441 35334
rect 5497 35278 5523 35334
rect 5579 35278 5605 35334
rect 5661 35278 5687 35334
rect 5743 35278 5769 35334
rect 5825 35278 5851 35334
rect 5907 35278 5933 35334
rect 5989 35278 6015 35334
rect 6071 35278 6097 35334
rect 6153 35278 6179 35334
rect 6235 35278 6261 35334
rect 6317 35278 6343 35334
rect 6399 35278 6425 35334
rect 6481 35278 6507 35334
rect 6563 35278 6589 35334
rect 6645 35278 6671 35334
rect 6727 35278 6753 35334
rect 6809 35317 6853 35334
rect 6909 35317 6941 35373
rect 6997 35317 7029 35373
rect 7085 35317 7117 35373
rect 7173 35317 7205 35373
rect 7261 35317 7293 35373
rect 7349 35317 7364 35373
rect 6809 35290 7364 35317
rect 6809 35278 6853 35290
rect 5186 35254 6853 35278
rect 5186 35198 5195 35254
rect 5251 35198 5277 35254
rect 5333 35198 5359 35254
rect 5415 35198 5441 35254
rect 5497 35198 5523 35254
rect 5579 35198 5605 35254
rect 5661 35198 5687 35254
rect 5743 35198 5769 35254
rect 5825 35198 5851 35254
rect 5907 35198 5933 35254
rect 5989 35198 6015 35254
rect 6071 35198 6097 35254
rect 6153 35198 6179 35254
rect 6235 35198 6261 35254
rect 6317 35198 6343 35254
rect 6399 35198 6425 35254
rect 6481 35198 6507 35254
rect 6563 35198 6589 35254
rect 6645 35198 6671 35254
rect 6727 35198 6753 35254
rect 6809 35234 6853 35254
rect 6909 35234 6941 35290
rect 6997 35234 7029 35290
rect 7085 35234 7117 35290
rect 7173 35234 7205 35290
rect 7261 35234 7293 35290
rect 7349 35234 7364 35290
rect 6809 35207 7364 35234
rect 6809 35198 6853 35207
rect 5186 35174 6853 35198
rect 5186 35118 5195 35174
rect 5251 35118 5277 35174
rect 5333 35118 5359 35174
rect 5415 35118 5441 35174
rect 5497 35118 5523 35174
rect 5579 35118 5605 35174
rect 5661 35118 5687 35174
rect 5743 35118 5769 35174
rect 5825 35118 5851 35174
rect 5907 35118 5933 35174
rect 5989 35118 6015 35174
rect 6071 35118 6097 35174
rect 6153 35118 6179 35174
rect 6235 35118 6261 35174
rect 6317 35118 6343 35174
rect 6399 35118 6425 35174
rect 6481 35118 6507 35174
rect 6563 35118 6589 35174
rect 6645 35118 6671 35174
rect 6727 35118 6753 35174
rect 6809 35151 6853 35174
rect 6909 35151 6941 35207
rect 6997 35151 7029 35207
rect 7085 35151 7117 35207
rect 7173 35151 7205 35207
rect 7261 35151 7293 35207
rect 7349 35151 7364 35207
rect 6809 35124 7364 35151
rect 6809 35118 6853 35124
rect 5186 35094 6853 35118
rect 5186 35038 5195 35094
rect 5251 35038 5277 35094
rect 5333 35038 5359 35094
rect 5415 35038 5441 35094
rect 5497 35038 5523 35094
rect 5579 35038 5605 35094
rect 5661 35038 5687 35094
rect 5743 35038 5769 35094
rect 5825 35038 5851 35094
rect 5907 35038 5933 35094
rect 5989 35038 6015 35094
rect 6071 35038 6097 35094
rect 6153 35038 6179 35094
rect 6235 35038 6261 35094
rect 6317 35038 6343 35094
rect 6399 35038 6425 35094
rect 6481 35038 6507 35094
rect 6563 35038 6589 35094
rect 6645 35038 6671 35094
rect 6727 35038 6753 35094
rect 6809 35068 6853 35094
rect 6909 35068 6941 35124
rect 6997 35068 7029 35124
rect 7085 35068 7117 35124
rect 7173 35068 7205 35124
rect 7261 35068 7293 35124
rect 7349 35070 7364 35124
rect 7349 35068 7357 35070
rect 6809 35063 7357 35068
tri 7357 35063 7364 35070 nw
rect 7593 35070 9771 38004
tri 7593 35063 7600 35070 ne
rect 7600 35063 9771 35070
rect 6809 35038 7309 35063
rect 5186 35015 7309 35038
tri 7309 35015 7357 35063 nw
tri 7600 35015 7648 35063 ne
rect 7648 35015 9771 35063
rect 5186 35014 7213 35015
rect 5186 34958 5195 35014
rect 5251 34958 5277 35014
rect 5333 34958 5359 35014
rect 5415 34958 5441 35014
rect 5497 34958 5523 35014
rect 5579 34958 5605 35014
rect 5661 34958 5687 35014
rect 5743 34958 5769 35014
rect 5825 34958 5851 35014
rect 5907 34958 5933 35014
rect 5989 34958 6015 35014
rect 6071 34958 6097 35014
rect 6153 34958 6179 35014
rect 6235 34958 6261 35014
rect 6317 34958 6343 35014
rect 6399 34958 6425 35014
rect 6481 34958 6507 35014
rect 6563 34958 6589 35014
rect 6645 34958 6671 35014
rect 6727 34958 6753 35014
rect 6809 35010 7213 35014
rect 6809 34958 6847 35010
rect 5186 34954 6847 34958
rect 6903 34954 6989 35010
rect 7045 34980 7213 35010
rect 7045 34954 7102 34980
rect 5186 34934 7102 34954
rect 5186 34878 5195 34934
rect 5251 34878 5277 34934
rect 5333 34878 5359 34934
rect 5415 34878 5441 34934
rect 5497 34878 5523 34934
rect 5579 34878 5605 34934
rect 5661 34878 5687 34934
rect 5743 34878 5769 34934
rect 5825 34878 5851 34934
rect 5907 34878 5933 34934
rect 5989 34878 6015 34934
rect 6071 34878 6097 34934
rect 6153 34878 6179 34934
rect 6235 34878 6261 34934
rect 6317 34878 6343 34934
rect 6399 34878 6425 34934
rect 6481 34878 6507 34934
rect 6563 34878 6589 34934
rect 6645 34878 6671 34934
rect 6727 34878 6753 34934
rect 6809 34924 7102 34934
rect 7158 34924 7213 34980
rect 6809 34923 7213 34924
rect 6809 34878 6847 34923
rect 5186 34867 6847 34878
rect 6903 34867 6989 34923
rect 7045 34919 7213 34923
tri 7213 34919 7309 35015 nw
tri 7648 34919 7744 35015 ne
rect 7744 34919 9771 35015
rect 7045 34867 7068 34919
rect 5186 34854 7068 34867
rect 5186 34798 5195 34854
rect 5251 34798 5277 34854
rect 5333 34798 5359 34854
rect 5415 34798 5441 34854
rect 5497 34798 5523 34854
rect 5579 34798 5605 34854
rect 5661 34798 5687 34854
rect 5743 34798 5769 34854
rect 5825 34798 5851 34854
rect 5907 34798 5933 34854
rect 5989 34798 6015 34854
rect 6071 34798 6097 34854
rect 6153 34798 6179 34854
rect 6235 34798 6261 34854
rect 6317 34798 6343 34854
rect 6399 34798 6425 34854
rect 6481 34798 6507 34854
rect 6563 34798 6589 34854
rect 6645 34798 6671 34854
rect 6727 34798 6753 34854
rect 6809 34835 7068 34854
rect 6809 34798 6847 34835
rect 5186 34779 6847 34798
rect 6903 34779 6989 34835
rect 7045 34779 7068 34835
rect 5186 34774 7068 34779
tri 7068 34774 7213 34919 nw
tri 7744 34774 7889 34919 ne
rect 7889 34774 9771 34919
rect 5186 34718 5195 34774
rect 5251 34718 5277 34774
rect 5333 34718 5359 34774
rect 5415 34718 5441 34774
rect 5497 34718 5523 34774
rect 5579 34718 5605 34774
rect 5661 34718 5687 34774
rect 5743 34718 5769 34774
rect 5825 34718 5851 34774
rect 5907 34718 5933 34774
rect 5989 34718 6015 34774
rect 6071 34718 6097 34774
rect 6153 34718 6179 34774
rect 6235 34718 6261 34774
rect 6317 34718 6343 34774
rect 6399 34718 6425 34774
rect 6481 34718 6507 34774
rect 6563 34718 6589 34774
rect 6645 34718 6671 34774
rect 6727 34718 6753 34774
rect 6809 34749 7043 34774
tri 7043 34749 7068 34774 nw
tri 7889 34749 7914 34774 ne
rect 7914 34749 9771 34774
rect 6809 34718 6928 34749
rect 5186 34695 6928 34718
rect 5186 34694 6847 34695
rect 5186 34638 5195 34694
rect 5251 34638 5277 34694
rect 5333 34638 5359 34694
rect 5415 34638 5441 34694
rect 5497 34638 5523 34694
rect 5579 34638 5605 34694
rect 5661 34638 5687 34694
rect 5743 34638 5769 34694
rect 5825 34638 5851 34694
rect 5907 34638 5933 34694
rect 5989 34638 6015 34694
rect 6071 34638 6097 34694
rect 6153 34638 6179 34694
rect 6235 34638 6261 34694
rect 6317 34638 6343 34694
rect 6399 34638 6425 34694
rect 6481 34638 6507 34694
rect 6563 34638 6589 34694
rect 6645 34638 6671 34694
rect 6727 34638 6753 34694
rect 6809 34639 6847 34694
rect 6903 34639 6928 34695
rect 6809 34638 6928 34639
rect 5186 34634 6928 34638
tri 6928 34634 7043 34749 nw
tri 7914 34634 8029 34749 ne
rect 8029 34634 9771 34749
rect 5186 34614 6845 34634
rect 5186 34558 5195 34614
rect 5251 34558 5277 34614
rect 5333 34558 5359 34614
rect 5415 34558 5441 34614
rect 5497 34558 5523 34614
rect 5579 34558 5605 34614
rect 5661 34558 5687 34614
rect 5743 34558 5769 34614
rect 5825 34558 5851 34614
rect 5907 34558 5933 34614
rect 5989 34558 6015 34614
rect 6071 34558 6097 34614
rect 6153 34558 6179 34614
rect 6235 34558 6261 34614
rect 6317 34558 6343 34614
rect 6399 34558 6425 34614
rect 6481 34558 6507 34614
rect 6563 34558 6589 34614
rect 6645 34558 6671 34614
rect 6727 34558 6753 34614
rect 6809 34558 6845 34614
rect 5186 34551 6845 34558
tri 6845 34551 6928 34634 nw
tri 8029 34551 8112 34634 ne
rect 8112 34551 9771 34634
rect 5186 34229 6523 34551
tri 6523 34229 6845 34551 nw
tri 8112 34529 8134 34551 ne
rect 8134 34529 9771 34551
tri 8134 34229 8434 34529 ne
rect 8434 34229 9771 34529
rect 9955 35045 12298 38008
rect 9955 34529 11857 35045
tri 11857 34604 12298 35045 nw
tri 9955 34229 10255 34529 ne
rect 10255 34229 11857 34529
rect 3100 34173 4647 34229
tri 4647 34173 4703 34229 nw
rect 5186 34173 6467 34229
tri 6467 34173 6523 34229 nw
tri 8434 34173 8490 34229 ne
rect 8490 34173 8580 34229
rect 8636 34173 8661 34229
rect 8717 34173 8742 34229
rect 8798 34173 8823 34229
rect 8879 34173 8904 34229
rect 8960 34173 8985 34229
rect 9041 34173 9066 34229
rect 3100 34149 4623 34173
tri 4623 34149 4647 34173 nw
rect 5186 34149 6443 34173
tri 6443 34149 6467 34173 nw
tri 8490 34149 8514 34173 ne
rect 8514 34149 9066 34173
rect 3100 34093 4567 34149
tri 4567 34093 4623 34149 nw
rect 5186 34093 6387 34149
tri 6387 34093 6443 34149 nw
tri 8514 34093 8570 34149 ne
rect 8570 34093 8580 34149
rect 8636 34093 8661 34149
rect 8717 34093 8742 34149
rect 8798 34093 8823 34149
rect 8879 34093 8904 34149
rect 8960 34093 8985 34149
rect 9041 34093 9066 34149
rect 3100 34092 4566 34093
tri 4566 34092 4567 34093 nw
rect 3100 34069 4543 34092
tri 4543 34069 4566 34092 nw
rect 3100 34013 4487 34069
tri 4487 34013 4543 34069 nw
rect 3100 33989 4463 34013
tri 4463 33989 4487 34013 nw
rect 3100 33933 4407 33989
tri 4407 33933 4463 33989 nw
rect 3100 33909 4383 33933
tri 4383 33909 4407 33933 nw
rect 3100 33853 4327 33909
tri 4327 33853 4383 33909 nw
rect 3100 33829 4303 33853
tri 4303 33829 4327 33853 nw
rect 3100 31694 4300 33829
tri 4300 33826 4303 33829 nw
rect 3100 31638 3109 31694
rect 3165 31638 3190 31694
rect 3246 31638 3271 31694
rect 3327 31638 3352 31694
rect 3408 31638 3433 31694
rect 3489 31638 3514 31694
rect 3100 31614 3514 31638
rect 3100 31558 3109 31614
rect 3165 31558 3190 31614
rect 3246 31558 3271 31614
rect 3327 31558 3352 31614
rect 3408 31558 3433 31614
rect 3489 31558 3514 31614
rect 3100 31534 3514 31558
rect 3100 31478 3109 31534
rect 3165 31478 3190 31534
rect 3246 31478 3271 31534
rect 3327 31478 3352 31534
rect 3408 31478 3433 31534
rect 3489 31478 3514 31534
rect 3100 31454 3514 31478
rect 3100 31398 3109 31454
rect 3165 31398 3190 31454
rect 3246 31398 3271 31454
rect 3327 31398 3352 31454
rect 3408 31398 3433 31454
rect 3489 31398 3514 31454
rect 3100 31374 3514 31398
rect 3100 31318 3109 31374
rect 3165 31318 3190 31374
rect 3246 31318 3271 31374
rect 3327 31318 3352 31374
rect 3408 31318 3433 31374
rect 3489 31318 3514 31374
rect 3100 31294 3514 31318
rect 3100 31238 3109 31294
rect 3165 31238 3190 31294
rect 3246 31238 3271 31294
rect 3327 31238 3352 31294
rect 3408 31238 3433 31294
rect 3489 31238 3514 31294
rect 3100 31214 3514 31238
rect 3100 31158 3109 31214
rect 3165 31158 3190 31214
rect 3246 31158 3271 31214
rect 3327 31158 3352 31214
rect 3408 31158 3433 31214
rect 3489 31158 3514 31214
rect 3100 31134 3514 31158
rect 3100 31078 3109 31134
rect 3165 31078 3190 31134
rect 3246 31078 3271 31134
rect 3327 31078 3352 31134
rect 3408 31078 3433 31134
rect 3489 31078 3514 31134
rect 3100 31054 3514 31078
rect 3100 30998 3109 31054
rect 3165 30998 3190 31054
rect 3246 30998 3271 31054
rect 3327 30998 3352 31054
rect 3408 30998 3433 31054
rect 3489 30998 3514 31054
rect 3100 30974 3514 30998
rect 3100 30918 3109 30974
rect 3165 30918 3190 30974
rect 3246 30918 3271 30974
rect 3327 30918 3352 30974
rect 3408 30918 3433 30974
rect 3489 30918 3514 30974
rect 3100 30894 3514 30918
rect 3100 30838 3109 30894
rect 3165 30838 3190 30894
rect 3246 30838 3271 30894
rect 3327 30838 3352 30894
rect 3408 30838 3433 30894
rect 3489 30838 3514 30894
rect 3100 30814 3514 30838
rect 3100 30758 3109 30814
rect 3165 30758 3190 30814
rect 3246 30758 3271 30814
rect 3327 30758 3352 30814
rect 3408 30758 3433 30814
rect 3489 30758 3514 30814
rect 3100 30734 3514 30758
rect 3100 30678 3109 30734
rect 3165 30678 3190 30734
rect 3246 30678 3271 30734
rect 3327 30678 3352 30734
rect 3408 30678 3433 30734
rect 3489 30678 3514 30734
rect 3100 30654 3514 30678
rect 3100 30598 3109 30654
rect 3165 30598 3190 30654
rect 3246 30598 3271 30654
rect 3327 30598 3352 30654
rect 3408 30598 3433 30654
rect 3489 30598 3514 30654
rect 3100 30574 3514 30598
rect 3100 30518 3109 30574
rect 3165 30518 3190 30574
rect 3246 30518 3271 30574
rect 3327 30518 3352 30574
rect 3408 30518 3433 30574
rect 3489 30518 3514 30574
rect 3100 30494 3514 30518
rect 3100 30438 3109 30494
rect 3165 30438 3190 30494
rect 3246 30438 3271 30494
rect 3327 30438 3352 30494
rect 3408 30438 3433 30494
rect 3489 30438 3514 30494
rect 3100 30414 3514 30438
rect 3100 30358 3109 30414
rect 3165 30358 3190 30414
rect 3246 30358 3271 30414
rect 3327 30358 3352 30414
rect 3408 30358 3433 30414
rect 3489 30358 3514 30414
rect 3100 30334 3514 30358
rect 3100 30278 3109 30334
rect 3165 30278 3190 30334
rect 3246 30278 3271 30334
rect 3327 30278 3352 30334
rect 3408 30278 3433 30334
rect 3489 30278 3514 30334
rect 3100 30254 3514 30278
rect 3100 30198 3109 30254
rect 3165 30198 3190 30254
rect 3246 30198 3271 30254
rect 3327 30198 3352 30254
rect 3408 30198 3433 30254
rect 3489 30198 3514 30254
rect 3100 30174 3514 30198
rect 3100 30118 3109 30174
rect 3165 30118 3190 30174
rect 3246 30118 3271 30174
rect 3327 30118 3352 30174
rect 3408 30118 3433 30174
rect 3489 30118 3514 30174
rect 3100 30094 3514 30118
rect 3100 30038 3109 30094
rect 3165 30038 3190 30094
rect 3246 30038 3271 30094
rect 3327 30038 3352 30094
rect 3408 30038 3433 30094
rect 3489 30038 3514 30094
rect 3100 30014 3514 30038
rect 3100 29958 3109 30014
rect 3165 29958 3190 30014
rect 3246 29958 3271 30014
rect 3327 29958 3352 30014
rect 3408 29958 3433 30014
rect 3489 29958 3514 30014
rect 4290 29958 4300 31694
rect 3100 27094 4300 29958
rect 3100 27038 3109 27094
rect 3165 27038 3190 27094
rect 3246 27038 3271 27094
rect 3327 27038 3352 27094
rect 3408 27038 3433 27094
rect 3489 27038 3514 27094
rect 3100 27014 3514 27038
rect 3100 26958 3109 27014
rect 3165 26958 3190 27014
rect 3246 26958 3271 27014
rect 3327 26958 3352 27014
rect 3408 26958 3433 27014
rect 3489 26958 3514 27014
rect 3100 26934 3514 26958
rect 3100 26878 3109 26934
rect 3165 26878 3190 26934
rect 3246 26878 3271 26934
rect 3327 26878 3352 26934
rect 3408 26878 3433 26934
rect 3489 26878 3514 26934
rect 3100 26854 3514 26878
rect 3100 26798 3109 26854
rect 3165 26798 3190 26854
rect 3246 26798 3271 26854
rect 3327 26798 3352 26854
rect 3408 26798 3433 26854
rect 3489 26798 3514 26854
rect 3100 26774 3514 26798
rect 3100 26718 3109 26774
rect 3165 26718 3190 26774
rect 3246 26718 3271 26774
rect 3327 26718 3352 26774
rect 3408 26718 3433 26774
rect 3489 26718 3514 26774
rect 3100 26694 3514 26718
rect 3100 26638 3109 26694
rect 3165 26638 3190 26694
rect 3246 26638 3271 26694
rect 3327 26638 3352 26694
rect 3408 26638 3433 26694
rect 3489 26638 3514 26694
rect 3100 26614 3514 26638
rect 3100 26558 3109 26614
rect 3165 26558 3190 26614
rect 3246 26558 3271 26614
rect 3327 26558 3352 26614
rect 3408 26558 3433 26614
rect 3489 26558 3514 26614
rect 3100 26534 3514 26558
rect 3100 26478 3109 26534
rect 3165 26478 3190 26534
rect 3246 26478 3271 26534
rect 3327 26478 3352 26534
rect 3408 26478 3433 26534
rect 3489 26478 3514 26534
rect 3100 26454 3514 26478
rect 3100 26398 3109 26454
rect 3165 26398 3190 26454
rect 3246 26398 3271 26454
rect 3327 26398 3352 26454
rect 3408 26398 3433 26454
rect 3489 26398 3514 26454
rect 3100 26374 3514 26398
rect 3100 26318 3109 26374
rect 3165 26318 3190 26374
rect 3246 26318 3271 26374
rect 3327 26318 3352 26374
rect 3408 26318 3433 26374
rect 3489 26318 3514 26374
rect 3100 26294 3514 26318
rect 3100 26238 3109 26294
rect 3165 26238 3190 26294
rect 3246 26238 3271 26294
rect 3327 26238 3352 26294
rect 3408 26238 3433 26294
rect 3489 26238 3514 26294
rect 3100 26214 3514 26238
rect 3100 26158 3109 26214
rect 3165 26158 3190 26214
rect 3246 26158 3271 26214
rect 3327 26158 3352 26214
rect 3408 26158 3433 26214
rect 3489 26158 3514 26214
rect 3100 26134 3514 26158
rect 3100 26078 3109 26134
rect 3165 26078 3190 26134
rect 3246 26078 3271 26134
rect 3327 26078 3352 26134
rect 3408 26078 3433 26134
rect 3489 26078 3514 26134
rect 3100 26054 3514 26078
rect 3100 25998 3109 26054
rect 3165 25998 3190 26054
rect 3246 25998 3271 26054
rect 3327 25998 3352 26054
rect 3408 25998 3433 26054
rect 3489 25998 3514 26054
rect 3100 25974 3514 25998
rect 3100 25918 3109 25974
rect 3165 25918 3190 25974
rect 3246 25918 3271 25974
rect 3327 25918 3352 25974
rect 3408 25918 3433 25974
rect 3489 25918 3514 25974
rect 3100 25894 3514 25918
rect 3100 25838 3109 25894
rect 3165 25838 3190 25894
rect 3246 25838 3271 25894
rect 3327 25838 3352 25894
rect 3408 25838 3433 25894
rect 3489 25838 3514 25894
rect 3100 25814 3514 25838
rect 3100 25758 3109 25814
rect 3165 25758 3190 25814
rect 3246 25758 3271 25814
rect 3327 25758 3352 25814
rect 3408 25758 3433 25814
rect 3489 25758 3514 25814
rect 3100 25734 3514 25758
rect 3100 25678 3109 25734
rect 3165 25678 3190 25734
rect 3246 25678 3271 25734
rect 3327 25678 3352 25734
rect 3408 25678 3433 25734
rect 3489 25678 3514 25734
rect 3100 25654 3514 25678
rect 3100 25598 3109 25654
rect 3165 25598 3190 25654
rect 3246 25598 3271 25654
rect 3327 25598 3352 25654
rect 3408 25598 3433 25654
rect 3489 25598 3514 25654
rect 3100 25574 3514 25598
rect 3100 25518 3109 25574
rect 3165 25518 3190 25574
rect 3246 25518 3271 25574
rect 3327 25518 3352 25574
rect 3408 25518 3433 25574
rect 3489 25518 3514 25574
rect 3100 25494 3514 25518
rect 3100 25438 3109 25494
rect 3165 25438 3190 25494
rect 3246 25438 3271 25494
rect 3327 25438 3352 25494
rect 3408 25438 3433 25494
rect 3489 25438 3514 25494
rect 3100 25414 3514 25438
rect 3100 25358 3109 25414
rect 3165 25358 3190 25414
rect 3246 25358 3271 25414
rect 3327 25358 3352 25414
rect 3408 25358 3433 25414
rect 3489 25358 3514 25414
rect 4290 25358 4300 27094
rect 3100 22494 4300 25358
rect 3100 22438 3109 22494
rect 3165 22438 3190 22494
rect 3246 22438 3271 22494
rect 3327 22438 3352 22494
rect 3408 22438 3433 22494
rect 3489 22438 3514 22494
rect 3100 22414 3514 22438
rect 3100 22358 3109 22414
rect 3165 22358 3190 22414
rect 3246 22358 3271 22414
rect 3327 22358 3352 22414
rect 3408 22358 3433 22414
rect 3489 22358 3514 22414
rect 3100 22334 3514 22358
rect 3100 22278 3109 22334
rect 3165 22278 3190 22334
rect 3246 22278 3271 22334
rect 3327 22278 3352 22334
rect 3408 22278 3433 22334
rect 3489 22278 3514 22334
rect 3100 22254 3514 22278
rect 3100 22198 3109 22254
rect 3165 22198 3190 22254
rect 3246 22198 3271 22254
rect 3327 22198 3352 22254
rect 3408 22198 3433 22254
rect 3489 22198 3514 22254
rect 3100 22174 3514 22198
rect 3100 22118 3109 22174
rect 3165 22118 3190 22174
rect 3246 22118 3271 22174
rect 3327 22118 3352 22174
rect 3408 22118 3433 22174
rect 3489 22118 3514 22174
rect 3100 22094 3514 22118
rect 3100 22038 3109 22094
rect 3165 22038 3190 22094
rect 3246 22038 3271 22094
rect 3327 22038 3352 22094
rect 3408 22038 3433 22094
rect 3489 22038 3514 22094
rect 3100 22014 3514 22038
rect 3100 21958 3109 22014
rect 3165 21958 3190 22014
rect 3246 21958 3271 22014
rect 3327 21958 3352 22014
rect 3408 21958 3433 22014
rect 3489 21958 3514 22014
rect 3100 21934 3514 21958
rect 3100 21878 3109 21934
rect 3165 21878 3190 21934
rect 3246 21878 3271 21934
rect 3327 21878 3352 21934
rect 3408 21878 3433 21934
rect 3489 21878 3514 21934
rect 3100 21854 3514 21878
rect 3100 21798 3109 21854
rect 3165 21798 3190 21854
rect 3246 21798 3271 21854
rect 3327 21798 3352 21854
rect 3408 21798 3433 21854
rect 3489 21798 3514 21854
rect 3100 21774 3514 21798
rect 3100 21718 3109 21774
rect 3165 21718 3190 21774
rect 3246 21718 3271 21774
rect 3327 21718 3352 21774
rect 3408 21718 3433 21774
rect 3489 21718 3514 21774
rect 3100 21694 3514 21718
rect 3100 21638 3109 21694
rect 3165 21638 3190 21694
rect 3246 21638 3271 21694
rect 3327 21638 3352 21694
rect 3408 21638 3433 21694
rect 3489 21638 3514 21694
rect 3100 21614 3514 21638
rect 3100 21558 3109 21614
rect 3165 21558 3190 21614
rect 3246 21558 3271 21614
rect 3327 21558 3352 21614
rect 3408 21558 3433 21614
rect 3489 21558 3514 21614
rect 3100 21534 3514 21558
rect 3100 21478 3109 21534
rect 3165 21478 3190 21534
rect 3246 21478 3271 21534
rect 3327 21478 3352 21534
rect 3408 21478 3433 21534
rect 3489 21478 3514 21534
rect 3100 21454 3514 21478
rect 3100 21398 3109 21454
rect 3165 21398 3190 21454
rect 3246 21398 3271 21454
rect 3327 21398 3352 21454
rect 3408 21398 3433 21454
rect 3489 21398 3514 21454
rect 3100 21374 3514 21398
rect 3100 21318 3109 21374
rect 3165 21318 3190 21374
rect 3246 21318 3271 21374
rect 3327 21318 3352 21374
rect 3408 21318 3433 21374
rect 3489 21318 3514 21374
rect 3100 21294 3514 21318
rect 3100 21238 3109 21294
rect 3165 21238 3190 21294
rect 3246 21238 3271 21294
rect 3327 21238 3352 21294
rect 3408 21238 3433 21294
rect 3489 21238 3514 21294
rect 3100 21214 3514 21238
rect 3100 21158 3109 21214
rect 3165 21158 3190 21214
rect 3246 21158 3271 21214
rect 3327 21158 3352 21214
rect 3408 21158 3433 21214
rect 3489 21158 3514 21214
rect 3100 21134 3514 21158
rect 3100 21078 3109 21134
rect 3165 21078 3190 21134
rect 3246 21078 3271 21134
rect 3327 21078 3352 21134
rect 3408 21078 3433 21134
rect 3489 21078 3514 21134
rect 3100 21054 3514 21078
rect 3100 20998 3109 21054
rect 3165 20998 3190 21054
rect 3246 20998 3271 21054
rect 3327 20998 3352 21054
rect 3408 20998 3433 21054
rect 3489 20998 3514 21054
rect 3100 20974 3514 20998
rect 3100 20918 3109 20974
rect 3165 20918 3190 20974
rect 3246 20918 3271 20974
rect 3327 20918 3352 20974
rect 3408 20918 3433 20974
rect 3489 20918 3514 20974
rect 3100 20894 3514 20918
rect 3100 20838 3109 20894
rect 3165 20838 3190 20894
rect 3246 20838 3271 20894
rect 3327 20838 3352 20894
rect 3408 20838 3433 20894
rect 3489 20838 3514 20894
rect 3100 20814 3514 20838
rect 3100 20758 3109 20814
rect 3165 20758 3190 20814
rect 3246 20758 3271 20814
rect 3327 20758 3352 20814
rect 3408 20758 3433 20814
rect 3489 20758 3514 20814
rect 4290 20918 4300 22494
rect 5186 31694 6386 34093
tri 6386 34092 6387 34093 nw
tri 8570 34092 8571 34093 ne
rect 5186 31638 5195 31694
rect 5251 31638 5276 31694
rect 5332 31638 5357 31694
rect 5413 31638 5438 31694
rect 5494 31638 5519 31694
rect 5575 31638 5600 31694
rect 5186 31614 5600 31638
rect 5186 31558 5195 31614
rect 5251 31558 5276 31614
rect 5332 31558 5357 31614
rect 5413 31558 5438 31614
rect 5494 31558 5519 31614
rect 5575 31558 5600 31614
rect 5186 31534 5600 31558
rect 5186 31478 5195 31534
rect 5251 31478 5276 31534
rect 5332 31478 5357 31534
rect 5413 31478 5438 31534
rect 5494 31478 5519 31534
rect 5575 31478 5600 31534
rect 5186 31454 5600 31478
rect 5186 31398 5195 31454
rect 5251 31398 5276 31454
rect 5332 31398 5357 31454
rect 5413 31398 5438 31454
rect 5494 31398 5519 31454
rect 5575 31398 5600 31454
rect 5186 31374 5600 31398
rect 5186 31318 5195 31374
rect 5251 31318 5276 31374
rect 5332 31318 5357 31374
rect 5413 31318 5438 31374
rect 5494 31318 5519 31374
rect 5575 31318 5600 31374
rect 5186 31294 5600 31318
rect 5186 31238 5195 31294
rect 5251 31238 5276 31294
rect 5332 31238 5357 31294
rect 5413 31238 5438 31294
rect 5494 31238 5519 31294
rect 5575 31238 5600 31294
rect 5186 31214 5600 31238
rect 5186 31158 5195 31214
rect 5251 31158 5276 31214
rect 5332 31158 5357 31214
rect 5413 31158 5438 31214
rect 5494 31158 5519 31214
rect 5575 31158 5600 31214
rect 5186 31134 5600 31158
rect 5186 31078 5195 31134
rect 5251 31078 5276 31134
rect 5332 31078 5357 31134
rect 5413 31078 5438 31134
rect 5494 31078 5519 31134
rect 5575 31078 5600 31134
rect 5186 31054 5600 31078
rect 5186 30998 5195 31054
rect 5251 30998 5276 31054
rect 5332 30998 5357 31054
rect 5413 30998 5438 31054
rect 5494 30998 5519 31054
rect 5575 30998 5600 31054
rect 5186 30974 5600 30998
rect 5186 30918 5195 30974
rect 5251 30918 5276 30974
rect 5332 30918 5357 30974
rect 5413 30918 5438 30974
rect 5494 30918 5519 30974
rect 5575 30918 5600 30974
rect 5186 30894 5600 30918
rect 5186 30838 5195 30894
rect 5251 30838 5276 30894
rect 5332 30838 5357 30894
rect 5413 30838 5438 30894
rect 5494 30838 5519 30894
rect 5575 30838 5600 30894
rect 5186 30814 5600 30838
rect 5186 30758 5195 30814
rect 5251 30758 5276 30814
rect 5332 30758 5357 30814
rect 5413 30758 5438 30814
rect 5494 30758 5519 30814
rect 5575 30758 5600 30814
rect 5186 30734 5600 30758
rect 5186 30678 5195 30734
rect 5251 30678 5276 30734
rect 5332 30678 5357 30734
rect 5413 30678 5438 30734
rect 5494 30678 5519 30734
rect 5575 30678 5600 30734
rect 5186 30654 5600 30678
rect 5186 30598 5195 30654
rect 5251 30598 5276 30654
rect 5332 30598 5357 30654
rect 5413 30598 5438 30654
rect 5494 30598 5519 30654
rect 5575 30598 5600 30654
rect 5186 30574 5600 30598
rect 5186 30518 5195 30574
rect 5251 30518 5276 30574
rect 5332 30518 5357 30574
rect 5413 30518 5438 30574
rect 5494 30518 5519 30574
rect 5575 30518 5600 30574
rect 5186 30494 5600 30518
rect 5186 30438 5195 30494
rect 5251 30438 5276 30494
rect 5332 30438 5357 30494
rect 5413 30438 5438 30494
rect 5494 30438 5519 30494
rect 5575 30438 5600 30494
rect 5186 30414 5600 30438
rect 5186 30358 5195 30414
rect 5251 30358 5276 30414
rect 5332 30358 5357 30414
rect 5413 30358 5438 30414
rect 5494 30358 5519 30414
rect 5575 30358 5600 30414
rect 5186 30334 5600 30358
rect 5186 30278 5195 30334
rect 5251 30278 5276 30334
rect 5332 30278 5357 30334
rect 5413 30278 5438 30334
rect 5494 30278 5519 30334
rect 5575 30278 5600 30334
rect 5186 30254 5600 30278
rect 5186 30198 5195 30254
rect 5251 30198 5276 30254
rect 5332 30198 5357 30254
rect 5413 30198 5438 30254
rect 5494 30198 5519 30254
rect 5575 30198 5600 30254
rect 5186 30174 5600 30198
rect 5186 30118 5195 30174
rect 5251 30118 5276 30174
rect 5332 30118 5357 30174
rect 5413 30118 5438 30174
rect 5494 30118 5519 30174
rect 5575 30118 5600 30174
rect 5186 30094 5600 30118
rect 5186 30038 5195 30094
rect 5251 30038 5276 30094
rect 5332 30038 5357 30094
rect 5413 30038 5438 30094
rect 5494 30038 5519 30094
rect 5575 30038 5600 30094
rect 5186 30014 5600 30038
rect 5186 29958 5195 30014
rect 5251 29958 5276 30014
rect 5332 29958 5357 30014
rect 5413 29958 5438 30014
rect 5494 29958 5519 30014
rect 5575 29958 5600 30014
rect 6376 29958 6386 31694
rect 5186 27094 6386 29958
rect 5186 27038 5195 27094
rect 5251 27038 5276 27094
rect 5332 27038 5357 27094
rect 5413 27038 5438 27094
rect 5494 27038 5519 27094
rect 5575 27038 5600 27094
rect 5186 27014 5600 27038
rect 5186 26958 5195 27014
rect 5251 26958 5276 27014
rect 5332 26958 5357 27014
rect 5413 26958 5438 27014
rect 5494 26958 5519 27014
rect 5575 26958 5600 27014
rect 5186 26934 5600 26958
rect 5186 26878 5195 26934
rect 5251 26878 5276 26934
rect 5332 26878 5357 26934
rect 5413 26878 5438 26934
rect 5494 26878 5519 26934
rect 5575 26878 5600 26934
rect 5186 26854 5600 26878
rect 5186 26798 5195 26854
rect 5251 26798 5276 26854
rect 5332 26798 5357 26854
rect 5413 26798 5438 26854
rect 5494 26798 5519 26854
rect 5575 26798 5600 26854
rect 5186 26774 5600 26798
rect 5186 26718 5195 26774
rect 5251 26718 5276 26774
rect 5332 26718 5357 26774
rect 5413 26718 5438 26774
rect 5494 26718 5519 26774
rect 5575 26718 5600 26774
rect 5186 26694 5600 26718
rect 5186 26638 5195 26694
rect 5251 26638 5276 26694
rect 5332 26638 5357 26694
rect 5413 26638 5438 26694
rect 5494 26638 5519 26694
rect 5575 26638 5600 26694
rect 5186 26614 5600 26638
rect 5186 26558 5195 26614
rect 5251 26558 5276 26614
rect 5332 26558 5357 26614
rect 5413 26558 5438 26614
rect 5494 26558 5519 26614
rect 5575 26558 5600 26614
rect 5186 26534 5600 26558
rect 5186 26478 5195 26534
rect 5251 26478 5276 26534
rect 5332 26478 5357 26534
rect 5413 26478 5438 26534
rect 5494 26478 5519 26534
rect 5575 26478 5600 26534
rect 5186 26454 5600 26478
rect 5186 26398 5195 26454
rect 5251 26398 5276 26454
rect 5332 26398 5357 26454
rect 5413 26398 5438 26454
rect 5494 26398 5519 26454
rect 5575 26398 5600 26454
rect 5186 26374 5600 26398
rect 5186 26318 5195 26374
rect 5251 26318 5276 26374
rect 5332 26318 5357 26374
rect 5413 26318 5438 26374
rect 5494 26318 5519 26374
rect 5575 26318 5600 26374
rect 5186 26294 5600 26318
rect 5186 26238 5195 26294
rect 5251 26238 5276 26294
rect 5332 26238 5357 26294
rect 5413 26238 5438 26294
rect 5494 26238 5519 26294
rect 5575 26238 5600 26294
rect 5186 26214 5600 26238
rect 5186 26158 5195 26214
rect 5251 26158 5276 26214
rect 5332 26158 5357 26214
rect 5413 26158 5438 26214
rect 5494 26158 5519 26214
rect 5575 26158 5600 26214
rect 5186 26134 5600 26158
rect 5186 26078 5195 26134
rect 5251 26078 5276 26134
rect 5332 26078 5357 26134
rect 5413 26078 5438 26134
rect 5494 26078 5519 26134
rect 5575 26078 5600 26134
rect 5186 26054 5600 26078
rect 5186 25998 5195 26054
rect 5251 25998 5276 26054
rect 5332 25998 5357 26054
rect 5413 25998 5438 26054
rect 5494 25998 5519 26054
rect 5575 25998 5600 26054
rect 5186 25974 5600 25998
rect 5186 25918 5195 25974
rect 5251 25918 5276 25974
rect 5332 25918 5357 25974
rect 5413 25918 5438 25974
rect 5494 25918 5519 25974
rect 5575 25918 5600 25974
rect 5186 25894 5600 25918
rect 5186 25838 5195 25894
rect 5251 25838 5276 25894
rect 5332 25838 5357 25894
rect 5413 25838 5438 25894
rect 5494 25838 5519 25894
rect 5575 25838 5600 25894
rect 5186 25814 5600 25838
rect 5186 25758 5195 25814
rect 5251 25758 5276 25814
rect 5332 25758 5357 25814
rect 5413 25758 5438 25814
rect 5494 25758 5519 25814
rect 5575 25758 5600 25814
rect 5186 25734 5600 25758
rect 5186 25678 5195 25734
rect 5251 25678 5276 25734
rect 5332 25678 5357 25734
rect 5413 25678 5438 25734
rect 5494 25678 5519 25734
rect 5575 25678 5600 25734
rect 5186 25654 5600 25678
rect 5186 25598 5195 25654
rect 5251 25598 5276 25654
rect 5332 25598 5357 25654
rect 5413 25598 5438 25654
rect 5494 25598 5519 25654
rect 5575 25598 5600 25654
rect 5186 25574 5600 25598
rect 5186 25518 5195 25574
rect 5251 25518 5276 25574
rect 5332 25518 5357 25574
rect 5413 25518 5438 25574
rect 5494 25518 5519 25574
rect 5575 25518 5600 25574
rect 5186 25494 5600 25518
rect 5186 25438 5195 25494
rect 5251 25438 5276 25494
rect 5332 25438 5357 25494
rect 5413 25438 5438 25494
rect 5494 25438 5519 25494
rect 5575 25438 5600 25494
rect 5186 25414 5600 25438
rect 5186 25358 5195 25414
rect 5251 25358 5276 25414
rect 5332 25358 5357 25414
rect 5413 25358 5438 25414
rect 5494 25358 5519 25414
rect 5575 25358 5600 25414
rect 6376 25358 6386 27094
rect 5186 22494 6386 25358
rect 5186 22438 5195 22494
rect 5251 22438 5276 22494
rect 5332 22438 5357 22494
rect 5413 22438 5438 22494
rect 5494 22438 5519 22494
rect 5575 22438 5600 22494
rect 5186 22414 5600 22438
rect 5186 22358 5195 22414
rect 5251 22358 5276 22414
rect 5332 22358 5357 22414
rect 5413 22358 5438 22414
rect 5494 22358 5519 22414
rect 5575 22358 5600 22414
rect 5186 22334 5600 22358
rect 5186 22278 5195 22334
rect 5251 22278 5276 22334
rect 5332 22278 5357 22334
rect 5413 22278 5438 22334
rect 5494 22278 5519 22334
rect 5575 22278 5600 22334
rect 5186 22254 5600 22278
rect 5186 22198 5195 22254
rect 5251 22198 5276 22254
rect 5332 22198 5357 22254
rect 5413 22198 5438 22254
rect 5494 22198 5519 22254
rect 5575 22198 5600 22254
rect 5186 22174 5600 22198
rect 5186 22118 5195 22174
rect 5251 22118 5276 22174
rect 5332 22118 5357 22174
rect 5413 22118 5438 22174
rect 5494 22118 5519 22174
rect 5575 22118 5600 22174
rect 5186 22094 5600 22118
rect 5186 22038 5195 22094
rect 5251 22038 5276 22094
rect 5332 22038 5357 22094
rect 5413 22038 5438 22094
rect 5494 22038 5519 22094
rect 5575 22038 5600 22094
rect 5186 22014 5600 22038
rect 5186 21958 5195 22014
rect 5251 21958 5276 22014
rect 5332 21958 5357 22014
rect 5413 21958 5438 22014
rect 5494 21958 5519 22014
rect 5575 21958 5600 22014
rect 5186 21934 5600 21958
rect 5186 21878 5195 21934
rect 5251 21878 5276 21934
rect 5332 21878 5357 21934
rect 5413 21878 5438 21934
rect 5494 21878 5519 21934
rect 5575 21878 5600 21934
rect 5186 21854 5600 21878
rect 5186 21798 5195 21854
rect 5251 21798 5276 21854
rect 5332 21798 5357 21854
rect 5413 21798 5438 21854
rect 5494 21798 5519 21854
rect 5575 21798 5600 21854
rect 5186 21774 5600 21798
rect 5186 21718 5195 21774
rect 5251 21718 5276 21774
rect 5332 21718 5357 21774
rect 5413 21718 5438 21774
rect 5494 21718 5519 21774
rect 5575 21718 5600 21774
rect 5186 21694 5600 21718
rect 5186 21638 5195 21694
rect 5251 21638 5276 21694
rect 5332 21638 5357 21694
rect 5413 21638 5438 21694
rect 5494 21638 5519 21694
rect 5575 21638 5600 21694
rect 5186 21614 5600 21638
rect 5186 21558 5195 21614
rect 5251 21558 5276 21614
rect 5332 21558 5357 21614
rect 5413 21558 5438 21614
rect 5494 21558 5519 21614
rect 5575 21558 5600 21614
rect 5186 21534 5600 21558
rect 5186 21478 5195 21534
rect 5251 21478 5276 21534
rect 5332 21478 5357 21534
rect 5413 21478 5438 21534
rect 5494 21478 5519 21534
rect 5575 21478 5600 21534
rect 5186 21454 5600 21478
rect 5186 21398 5195 21454
rect 5251 21398 5276 21454
rect 5332 21398 5357 21454
rect 5413 21398 5438 21454
rect 5494 21398 5519 21454
rect 5575 21398 5600 21454
rect 5186 21374 5600 21398
rect 5186 21318 5195 21374
rect 5251 21318 5276 21374
rect 5332 21318 5357 21374
rect 5413 21318 5438 21374
rect 5494 21318 5519 21374
rect 5575 21318 5600 21374
rect 5186 21294 5600 21318
rect 5186 21238 5195 21294
rect 5251 21238 5276 21294
rect 5332 21238 5357 21294
rect 5413 21238 5438 21294
rect 5494 21238 5519 21294
rect 5575 21238 5600 21294
rect 5186 21214 5600 21238
rect 5186 21158 5195 21214
rect 5251 21158 5276 21214
rect 5332 21158 5357 21214
rect 5413 21158 5438 21214
rect 5494 21158 5519 21214
rect 5575 21158 5600 21214
rect 5186 21134 5600 21158
rect 5186 21078 5195 21134
rect 5251 21078 5276 21134
rect 5332 21078 5357 21134
rect 5413 21078 5438 21134
rect 5494 21078 5519 21134
rect 5575 21078 5600 21134
rect 5186 21054 5600 21078
rect 5186 20998 5195 21054
rect 5251 20998 5276 21054
rect 5332 20998 5357 21054
rect 5413 20998 5438 21054
rect 5494 20998 5519 21054
rect 5575 20998 5600 21054
rect 5186 20974 5600 20998
tri 4300 20918 4318 20936 sw
rect 5186 20918 5195 20974
rect 5251 20918 5276 20974
rect 5332 20918 5357 20974
rect 5413 20918 5438 20974
rect 5494 20918 5519 20974
rect 5575 20918 5600 20974
rect 4290 20894 4318 20918
tri 4318 20894 4342 20918 sw
rect 5186 20894 5600 20918
rect 4290 20838 4342 20894
tri 4342 20838 4398 20894 sw
rect 5186 20838 5195 20894
rect 5251 20838 5276 20894
rect 5332 20838 5357 20894
rect 5413 20838 5438 20894
rect 5494 20838 5519 20894
rect 5575 20838 5600 20894
rect 4290 20814 4398 20838
tri 4398 20814 4422 20838 sw
rect 5186 20814 5600 20838
rect 4290 20758 4422 20814
tri 4422 20758 4478 20814 sw
rect 5186 20758 5195 20814
rect 5251 20758 5276 20814
rect 5332 20758 5357 20814
rect 5413 20758 5438 20814
rect 5494 20758 5519 20814
rect 5575 20758 5600 20814
rect 6376 20758 6386 22494
rect 8571 34069 9066 34093
rect 8571 34013 8580 34069
rect 8636 34013 8661 34069
rect 8717 34013 8742 34069
rect 8798 34013 8823 34069
rect 8879 34013 8904 34069
rect 8960 34013 8985 34069
rect 9041 34013 9066 34069
rect 8571 33989 9066 34013
rect 8571 33933 8580 33989
rect 8636 33933 8661 33989
rect 8717 33933 8742 33989
rect 8798 33933 8823 33989
rect 8879 33933 8904 33989
rect 8960 33933 8985 33989
rect 9041 33933 9066 33989
rect 8571 33909 9066 33933
rect 8571 33853 8580 33909
rect 8636 33853 8661 33909
rect 8717 33853 8742 33909
rect 8798 33853 8823 33909
rect 8879 33853 8904 33909
rect 8960 33853 8985 33909
rect 9041 33853 9066 33909
rect 8571 33829 9066 33853
rect 8571 33773 8580 33829
rect 8636 33773 8661 33829
rect 8717 33773 8742 33829
rect 8798 33773 8823 33829
rect 8879 33773 8904 33829
rect 8960 33773 8985 33829
rect 9041 33773 9066 33829
rect 8571 33749 9066 33773
rect 8571 33693 8580 33749
rect 8636 33693 8661 33749
rect 8717 33693 8742 33749
rect 8798 33693 8823 33749
rect 8879 33693 8904 33749
rect 8960 33693 8985 33749
rect 9041 33693 9066 33749
rect 8571 33669 9066 33693
rect 8571 33613 8580 33669
rect 8636 33613 8661 33669
rect 8717 33613 8742 33669
rect 8798 33613 8823 33669
rect 8879 33613 8904 33669
rect 8960 33613 8985 33669
rect 9041 33613 9066 33669
rect 8571 33589 9066 33613
rect 8571 33533 8580 33589
rect 8636 33533 8661 33589
rect 8717 33533 8742 33589
rect 8798 33533 8823 33589
rect 8879 33533 8904 33589
rect 8960 33533 8985 33589
rect 9041 33533 9066 33589
rect 8571 33509 9066 33533
rect 8571 33453 8580 33509
rect 8636 33453 8661 33509
rect 8717 33453 8742 33509
rect 8798 33453 8823 33509
rect 8879 33453 8904 33509
rect 8960 33453 8985 33509
rect 9041 33453 9066 33509
rect 8571 33429 9066 33453
rect 8571 33373 8580 33429
rect 8636 33373 8661 33429
rect 8717 33373 8742 33429
rect 8798 33373 8823 33429
rect 8879 33373 8904 33429
rect 8960 33373 8985 33429
rect 9041 33373 9066 33429
rect 8571 33349 9066 33373
rect 8571 33293 8580 33349
rect 8636 33293 8661 33349
rect 8717 33293 8742 33349
rect 8798 33293 8823 33349
rect 8879 33293 8904 33349
rect 8960 33293 8985 33349
rect 9041 33293 9066 33349
rect 8571 33269 9066 33293
rect 8571 33213 8580 33269
rect 8636 33213 8661 33269
rect 8717 33213 8742 33269
rect 8798 33213 8823 33269
rect 8879 33213 8904 33269
rect 8960 33213 8985 33269
rect 9041 33213 9066 33269
rect 8571 33189 9066 33213
rect 8571 33133 8580 33189
rect 8636 33133 8661 33189
rect 8717 33133 8742 33189
rect 8798 33133 8823 33189
rect 8879 33133 8904 33189
rect 8960 33133 8985 33189
rect 9041 33133 9066 33189
rect 8571 33109 9066 33133
rect 8571 33053 8580 33109
rect 8636 33053 8661 33109
rect 8717 33053 8742 33109
rect 8798 33053 8823 33109
rect 8879 33053 8904 33109
rect 8960 33053 8985 33109
rect 9041 33053 9066 33109
rect 8571 33029 9066 33053
rect 8571 32973 8580 33029
rect 8636 32973 8661 33029
rect 8717 32973 8742 33029
rect 8798 32973 8823 33029
rect 8879 32973 8904 33029
rect 8960 32973 8985 33029
rect 9041 32973 9066 33029
rect 8571 32949 9066 32973
rect 8571 32893 8580 32949
rect 8636 32893 8661 32949
rect 8717 32893 8742 32949
rect 8798 32893 8823 32949
rect 8879 32893 8904 32949
rect 8960 32893 8985 32949
rect 9041 32893 9066 32949
rect 8571 32869 9066 32893
rect 8571 32813 8580 32869
rect 8636 32813 8661 32869
rect 8717 32813 8742 32869
rect 8798 32813 8823 32869
rect 8879 32813 8904 32869
rect 8960 32813 8985 32869
rect 9041 32813 9066 32869
rect 8571 32789 9066 32813
rect 8571 32733 8580 32789
rect 8636 32733 8661 32789
rect 8717 32733 8742 32789
rect 8798 32733 8823 32789
rect 8879 32733 8904 32789
rect 8960 32733 8985 32789
rect 9041 32733 9066 32789
rect 8571 32709 9066 32733
rect 8571 32653 8580 32709
rect 8636 32653 8661 32709
rect 8717 32653 8742 32709
rect 8798 32653 8823 32709
rect 8879 32653 8904 32709
rect 8960 32653 8985 32709
rect 9041 32653 9066 32709
rect 8571 32629 9066 32653
rect 8571 32573 8580 32629
rect 8636 32573 8661 32629
rect 8717 32573 8742 32629
rect 8798 32573 8823 32629
rect 8879 32573 8904 32629
rect 8960 32573 8985 32629
rect 9041 32573 9066 32629
rect 8571 32549 9066 32573
rect 8571 32493 8580 32549
rect 8636 32493 8661 32549
rect 8717 32493 8742 32549
rect 8798 32493 8823 32549
rect 8879 32493 8904 32549
rect 8960 32493 8985 32549
rect 9041 32493 9066 32549
rect 9762 32493 9771 34229
tri 10255 34173 10311 34229 ne
rect 10311 34173 10666 34229
rect 10722 34173 10747 34229
rect 10803 34173 10828 34229
rect 10884 34173 10909 34229
rect 10965 34173 10990 34229
rect 11046 34173 11071 34229
rect 11127 34173 11152 34229
tri 10311 34149 10335 34173 ne
rect 10335 34149 11152 34173
tri 10335 34093 10391 34149 ne
rect 10391 34093 10666 34149
rect 10722 34093 10747 34149
rect 10803 34093 10828 34149
rect 10884 34093 10909 34149
rect 10965 34093 10990 34149
rect 11046 34093 11071 34149
rect 11127 34093 11152 34149
tri 10391 34092 10392 34093 ne
rect 10392 34092 11152 34093
tri 10392 34069 10415 34092 ne
rect 10415 34069 11152 34092
tri 10415 34013 10471 34069 ne
rect 10471 34013 10666 34069
rect 10722 34013 10747 34069
rect 10803 34013 10828 34069
rect 10884 34013 10909 34069
rect 10965 34013 10990 34069
rect 11046 34013 11071 34069
rect 11127 34013 11152 34069
tri 10471 33989 10495 34013 ne
rect 10495 33989 11152 34013
tri 10495 33933 10551 33989 ne
rect 10551 33933 10666 33989
rect 10722 33933 10747 33989
rect 10803 33933 10828 33989
rect 10884 33933 10909 33989
rect 10965 33933 10990 33989
rect 11046 33933 11071 33989
rect 11127 33933 11152 33989
tri 10551 33909 10575 33933 ne
rect 10575 33909 11152 33933
tri 10575 33853 10631 33909 ne
rect 10631 33853 10666 33909
rect 10722 33853 10747 33909
rect 10803 33853 10828 33909
rect 10884 33853 10909 33909
rect 10965 33853 10990 33909
rect 11046 33853 11071 33909
rect 11127 33853 11152 33909
tri 10631 33829 10655 33853 ne
rect 10655 33829 11152 33853
tri 10655 33827 10657 33829 ne
rect 8571 29629 9771 32493
rect 8571 29573 8580 29629
rect 8636 29573 8661 29629
rect 8717 29573 8742 29629
rect 8798 29573 8823 29629
rect 8879 29573 8904 29629
rect 8960 29573 8985 29629
rect 9041 29573 9066 29629
rect 8571 29549 9066 29573
rect 8571 29493 8580 29549
rect 8636 29493 8661 29549
rect 8717 29493 8742 29549
rect 8798 29493 8823 29549
rect 8879 29493 8904 29549
rect 8960 29493 8985 29549
rect 9041 29493 9066 29549
rect 8571 29469 9066 29493
rect 8571 29413 8580 29469
rect 8636 29413 8661 29469
rect 8717 29413 8742 29469
rect 8798 29413 8823 29469
rect 8879 29413 8904 29469
rect 8960 29413 8985 29469
rect 9041 29413 9066 29469
rect 8571 29389 9066 29413
rect 8571 29333 8580 29389
rect 8636 29333 8661 29389
rect 8717 29333 8742 29389
rect 8798 29333 8823 29389
rect 8879 29333 8904 29389
rect 8960 29333 8985 29389
rect 9041 29333 9066 29389
rect 8571 29309 9066 29333
rect 8571 29253 8580 29309
rect 8636 29253 8661 29309
rect 8717 29253 8742 29309
rect 8798 29253 8823 29309
rect 8879 29253 8904 29309
rect 8960 29253 8985 29309
rect 9041 29253 9066 29309
rect 8571 29229 9066 29253
rect 8571 29173 8580 29229
rect 8636 29173 8661 29229
rect 8717 29173 8742 29229
rect 8798 29173 8823 29229
rect 8879 29173 8904 29229
rect 8960 29173 8985 29229
rect 9041 29173 9066 29229
rect 8571 29149 9066 29173
rect 8571 29093 8580 29149
rect 8636 29093 8661 29149
rect 8717 29093 8742 29149
rect 8798 29093 8823 29149
rect 8879 29093 8904 29149
rect 8960 29093 8985 29149
rect 9041 29093 9066 29149
rect 8571 29069 9066 29093
rect 8571 29013 8580 29069
rect 8636 29013 8661 29069
rect 8717 29013 8742 29069
rect 8798 29013 8823 29069
rect 8879 29013 8904 29069
rect 8960 29013 8985 29069
rect 9041 29013 9066 29069
rect 8571 28989 9066 29013
rect 8571 28933 8580 28989
rect 8636 28933 8661 28989
rect 8717 28933 8742 28989
rect 8798 28933 8823 28989
rect 8879 28933 8904 28989
rect 8960 28933 8985 28989
rect 9041 28933 9066 28989
rect 8571 28909 9066 28933
rect 8571 28853 8580 28909
rect 8636 28853 8661 28909
rect 8717 28853 8742 28909
rect 8798 28853 8823 28909
rect 8879 28853 8904 28909
rect 8960 28853 8985 28909
rect 9041 28853 9066 28909
rect 8571 28829 9066 28853
rect 8571 28773 8580 28829
rect 8636 28773 8661 28829
rect 8717 28773 8742 28829
rect 8798 28773 8823 28829
rect 8879 28773 8904 28829
rect 8960 28773 8985 28829
rect 9041 28773 9066 28829
rect 8571 28749 9066 28773
rect 8571 28693 8580 28749
rect 8636 28693 8661 28749
rect 8717 28693 8742 28749
rect 8798 28693 8823 28749
rect 8879 28693 8904 28749
rect 8960 28693 8985 28749
rect 9041 28693 9066 28749
rect 8571 28669 9066 28693
rect 8571 28613 8580 28669
rect 8636 28613 8661 28669
rect 8717 28613 8742 28669
rect 8798 28613 8823 28669
rect 8879 28613 8904 28669
rect 8960 28613 8985 28669
rect 9041 28613 9066 28669
rect 8571 28589 9066 28613
rect 8571 28533 8580 28589
rect 8636 28533 8661 28589
rect 8717 28533 8742 28589
rect 8798 28533 8823 28589
rect 8879 28533 8904 28589
rect 8960 28533 8985 28589
rect 9041 28533 9066 28589
rect 8571 28509 9066 28533
rect 8571 28453 8580 28509
rect 8636 28453 8661 28509
rect 8717 28453 8742 28509
rect 8798 28453 8823 28509
rect 8879 28453 8904 28509
rect 8960 28453 8985 28509
rect 9041 28453 9066 28509
rect 8571 28429 9066 28453
rect 8571 28373 8580 28429
rect 8636 28373 8661 28429
rect 8717 28373 8742 28429
rect 8798 28373 8823 28429
rect 8879 28373 8904 28429
rect 8960 28373 8985 28429
rect 9041 28373 9066 28429
rect 8571 28349 9066 28373
rect 8571 28293 8580 28349
rect 8636 28293 8661 28349
rect 8717 28293 8742 28349
rect 8798 28293 8823 28349
rect 8879 28293 8904 28349
rect 8960 28293 8985 28349
rect 9041 28293 9066 28349
rect 8571 28269 9066 28293
rect 8571 28213 8580 28269
rect 8636 28213 8661 28269
rect 8717 28213 8742 28269
rect 8798 28213 8823 28269
rect 8879 28213 8904 28269
rect 8960 28213 8985 28269
rect 9041 28213 9066 28269
rect 8571 28189 9066 28213
rect 8571 28133 8580 28189
rect 8636 28133 8661 28189
rect 8717 28133 8742 28189
rect 8798 28133 8823 28189
rect 8879 28133 8904 28189
rect 8960 28133 8985 28189
rect 9041 28133 9066 28189
rect 8571 28109 9066 28133
rect 8571 28053 8580 28109
rect 8636 28053 8661 28109
rect 8717 28053 8742 28109
rect 8798 28053 8823 28109
rect 8879 28053 8904 28109
rect 8960 28053 8985 28109
rect 9041 28053 9066 28109
rect 8571 28029 9066 28053
rect 8571 27973 8580 28029
rect 8636 27973 8661 28029
rect 8717 27973 8742 28029
rect 8798 27973 8823 28029
rect 8879 27973 8904 28029
rect 8960 27973 8985 28029
rect 9041 27973 9066 28029
rect 8571 27949 9066 27973
rect 8571 27893 8580 27949
rect 8636 27893 8661 27949
rect 8717 27893 8742 27949
rect 8798 27893 8823 27949
rect 8879 27893 8904 27949
rect 8960 27893 8985 27949
rect 9041 27893 9066 27949
rect 9762 27893 9771 29629
rect 8571 25029 9771 27893
rect 8571 24973 8580 25029
rect 8636 24973 8661 25029
rect 8717 24973 8742 25029
rect 8798 24973 8823 25029
rect 8879 24973 8904 25029
rect 8960 24973 8985 25029
rect 9041 24973 9066 25029
rect 8571 24949 9066 24973
rect 8571 24893 8580 24949
rect 8636 24893 8661 24949
rect 8717 24893 8742 24949
rect 8798 24893 8823 24949
rect 8879 24893 8904 24949
rect 8960 24893 8985 24949
rect 9041 24893 9066 24949
rect 8571 24869 9066 24893
rect 8571 24813 8580 24869
rect 8636 24813 8661 24869
rect 8717 24813 8742 24869
rect 8798 24813 8823 24869
rect 8879 24813 8904 24869
rect 8960 24813 8985 24869
rect 9041 24813 9066 24869
rect 8571 24789 9066 24813
rect 8571 24733 8580 24789
rect 8636 24733 8661 24789
rect 8717 24733 8742 24789
rect 8798 24733 8823 24789
rect 8879 24733 8904 24789
rect 8960 24733 8985 24789
rect 9041 24733 9066 24789
rect 8571 24709 9066 24733
rect 8571 24653 8580 24709
rect 8636 24653 8661 24709
rect 8717 24653 8742 24709
rect 8798 24653 8823 24709
rect 8879 24653 8904 24709
rect 8960 24653 8985 24709
rect 9041 24653 9066 24709
rect 8571 24629 9066 24653
rect 8571 24573 8580 24629
rect 8636 24573 8661 24629
rect 8717 24573 8742 24629
rect 8798 24573 8823 24629
rect 8879 24573 8904 24629
rect 8960 24573 8985 24629
rect 9041 24573 9066 24629
rect 8571 24549 9066 24573
rect 8571 24493 8580 24549
rect 8636 24493 8661 24549
rect 8717 24493 8742 24549
rect 8798 24493 8823 24549
rect 8879 24493 8904 24549
rect 8960 24493 8985 24549
rect 9041 24493 9066 24549
rect 8571 24469 9066 24493
rect 8571 24413 8580 24469
rect 8636 24413 8661 24469
rect 8717 24413 8742 24469
rect 8798 24413 8823 24469
rect 8879 24413 8904 24469
rect 8960 24413 8985 24469
rect 9041 24413 9066 24469
rect 8571 24389 9066 24413
rect 8571 24333 8580 24389
rect 8636 24333 8661 24389
rect 8717 24333 8742 24389
rect 8798 24333 8823 24389
rect 8879 24333 8904 24389
rect 8960 24333 8985 24389
rect 9041 24333 9066 24389
rect 8571 24309 9066 24333
rect 8571 24253 8580 24309
rect 8636 24253 8661 24309
rect 8717 24253 8742 24309
rect 8798 24253 8823 24309
rect 8879 24253 8904 24309
rect 8960 24253 8985 24309
rect 9041 24253 9066 24309
rect 8571 24229 9066 24253
rect 8571 24173 8580 24229
rect 8636 24173 8661 24229
rect 8717 24173 8742 24229
rect 8798 24173 8823 24229
rect 8879 24173 8904 24229
rect 8960 24173 8985 24229
rect 9041 24173 9066 24229
rect 8571 24149 9066 24173
rect 8571 24093 8580 24149
rect 8636 24093 8661 24149
rect 8717 24093 8742 24149
rect 8798 24093 8823 24149
rect 8879 24093 8904 24149
rect 8960 24093 8985 24149
rect 9041 24093 9066 24149
rect 8571 24069 9066 24093
rect 8571 24013 8580 24069
rect 8636 24013 8661 24069
rect 8717 24013 8742 24069
rect 8798 24013 8823 24069
rect 8879 24013 8904 24069
rect 8960 24013 8985 24069
rect 9041 24013 9066 24069
rect 8571 23989 9066 24013
rect 8571 23933 8580 23989
rect 8636 23933 8661 23989
rect 8717 23933 8742 23989
rect 8798 23933 8823 23989
rect 8879 23933 8904 23989
rect 8960 23933 8985 23989
rect 9041 23933 9066 23989
rect 8571 23909 9066 23933
rect 8571 23853 8580 23909
rect 8636 23853 8661 23909
rect 8717 23853 8742 23909
rect 8798 23853 8823 23909
rect 8879 23853 8904 23909
rect 8960 23853 8985 23909
rect 9041 23853 9066 23909
rect 8571 23829 9066 23853
rect 8571 23773 8580 23829
rect 8636 23773 8661 23829
rect 8717 23773 8742 23829
rect 8798 23773 8823 23829
rect 8879 23773 8904 23829
rect 8960 23773 8985 23829
rect 9041 23773 9066 23829
rect 8571 23749 9066 23773
rect 8571 23693 8580 23749
rect 8636 23693 8661 23749
rect 8717 23693 8742 23749
rect 8798 23693 8823 23749
rect 8879 23693 8904 23749
rect 8960 23693 8985 23749
rect 9041 23693 9066 23749
rect 8571 23669 9066 23693
rect 8571 23613 8580 23669
rect 8636 23613 8661 23669
rect 8717 23613 8742 23669
rect 8798 23613 8823 23669
rect 8879 23613 8904 23669
rect 8960 23613 8985 23669
rect 9041 23613 9066 23669
rect 8571 23589 9066 23613
rect 8571 23533 8580 23589
rect 8636 23533 8661 23589
rect 8717 23533 8742 23589
rect 8798 23533 8823 23589
rect 8879 23533 8904 23589
rect 8960 23533 8985 23589
rect 9041 23533 9066 23589
rect 8571 23509 9066 23533
rect 8571 23453 8580 23509
rect 8636 23453 8661 23509
rect 8717 23453 8742 23509
rect 8798 23453 8823 23509
rect 8879 23453 8904 23509
rect 8960 23453 8985 23509
rect 9041 23453 9066 23509
rect 8571 23429 9066 23453
rect 8571 23373 8580 23429
rect 8636 23373 8661 23429
rect 8717 23373 8742 23429
rect 8798 23373 8823 23429
rect 8879 23373 8904 23429
rect 8960 23373 8985 23429
rect 9041 23373 9066 23429
rect 8571 23349 9066 23373
rect 8571 23293 8580 23349
rect 8636 23293 8661 23349
rect 8717 23293 8742 23349
rect 8798 23293 8823 23349
rect 8879 23293 8904 23349
rect 8960 23293 8985 23349
rect 9041 23293 9066 23349
rect 9762 23293 9771 25029
tri 8535 22088 8571 22124 se
rect 8571 22088 9771 23293
rect 10657 33773 10666 33829
rect 10722 33773 10747 33829
rect 10803 33773 10828 33829
rect 10884 33773 10909 33829
rect 10965 33773 10990 33829
rect 11046 33773 11071 33829
rect 11127 33773 11152 33829
rect 10657 33749 11152 33773
rect 10657 33693 10666 33749
rect 10722 33693 10747 33749
rect 10803 33693 10828 33749
rect 10884 33693 10909 33749
rect 10965 33693 10990 33749
rect 11046 33693 11071 33749
rect 11127 33693 11152 33749
rect 10657 33669 11152 33693
rect 10657 33613 10666 33669
rect 10722 33613 10747 33669
rect 10803 33613 10828 33669
rect 10884 33613 10909 33669
rect 10965 33613 10990 33669
rect 11046 33613 11071 33669
rect 11127 33613 11152 33669
rect 10657 33589 11152 33613
rect 10657 33533 10666 33589
rect 10722 33533 10747 33589
rect 10803 33533 10828 33589
rect 10884 33533 10909 33589
rect 10965 33533 10990 33589
rect 11046 33533 11071 33589
rect 11127 33533 11152 33589
rect 10657 33509 11152 33533
rect 10657 33453 10666 33509
rect 10722 33453 10747 33509
rect 10803 33453 10828 33509
rect 10884 33453 10909 33509
rect 10965 33453 10990 33509
rect 11046 33453 11071 33509
rect 11127 33453 11152 33509
rect 10657 33429 11152 33453
rect 10657 33373 10666 33429
rect 10722 33373 10747 33429
rect 10803 33373 10828 33429
rect 10884 33373 10909 33429
rect 10965 33373 10990 33429
rect 11046 33373 11071 33429
rect 11127 33373 11152 33429
rect 10657 33349 11152 33373
rect 10657 33293 10666 33349
rect 10722 33293 10747 33349
rect 10803 33293 10828 33349
rect 10884 33293 10909 33349
rect 10965 33293 10990 33349
rect 11046 33293 11071 33349
rect 11127 33293 11152 33349
rect 10657 33269 11152 33293
rect 10657 33213 10666 33269
rect 10722 33213 10747 33269
rect 10803 33213 10828 33269
rect 10884 33213 10909 33269
rect 10965 33213 10990 33269
rect 11046 33213 11071 33269
rect 11127 33213 11152 33269
rect 10657 33189 11152 33213
rect 10657 33133 10666 33189
rect 10722 33133 10747 33189
rect 10803 33133 10828 33189
rect 10884 33133 10909 33189
rect 10965 33133 10990 33189
rect 11046 33133 11071 33189
rect 11127 33133 11152 33189
rect 10657 33109 11152 33133
rect 10657 33053 10666 33109
rect 10722 33053 10747 33109
rect 10803 33053 10828 33109
rect 10884 33053 10909 33109
rect 10965 33053 10990 33109
rect 11046 33053 11071 33109
rect 11127 33053 11152 33109
rect 10657 33029 11152 33053
rect 10657 32973 10666 33029
rect 10722 32973 10747 33029
rect 10803 32973 10828 33029
rect 10884 32973 10909 33029
rect 10965 32973 10990 33029
rect 11046 32973 11071 33029
rect 11127 32973 11152 33029
rect 10657 32949 11152 32973
rect 10657 32893 10666 32949
rect 10722 32893 10747 32949
rect 10803 32893 10828 32949
rect 10884 32893 10909 32949
rect 10965 32893 10990 32949
rect 11046 32893 11071 32949
rect 11127 32893 11152 32949
rect 10657 32869 11152 32893
rect 10657 32813 10666 32869
rect 10722 32813 10747 32869
rect 10803 32813 10828 32869
rect 10884 32813 10909 32869
rect 10965 32813 10990 32869
rect 11046 32813 11071 32869
rect 11127 32813 11152 32869
rect 10657 32789 11152 32813
rect 10657 32733 10666 32789
rect 10722 32733 10747 32789
rect 10803 32733 10828 32789
rect 10884 32733 10909 32789
rect 10965 32733 10990 32789
rect 11046 32733 11071 32789
rect 11127 32733 11152 32789
rect 10657 32709 11152 32733
rect 10657 32653 10666 32709
rect 10722 32653 10747 32709
rect 10803 32653 10828 32709
rect 10884 32653 10909 32709
rect 10965 32653 10990 32709
rect 11046 32653 11071 32709
rect 11127 32653 11152 32709
rect 10657 32629 11152 32653
rect 10657 32573 10666 32629
rect 10722 32573 10747 32629
rect 10803 32573 10828 32629
rect 10884 32573 10909 32629
rect 10965 32573 10990 32629
rect 11046 32573 11071 32629
rect 11127 32573 11152 32629
rect 10657 32549 11152 32573
rect 10657 32493 10666 32549
rect 10722 32493 10747 32549
rect 10803 32493 10828 32549
rect 10884 32493 10909 32549
rect 10965 32493 10990 32549
rect 11046 32493 11071 32549
rect 11127 32493 11152 32549
rect 11848 32493 11857 34229
rect 10657 29629 11857 32493
rect 10657 29573 10666 29629
rect 10722 29573 10747 29629
rect 10803 29573 10828 29629
rect 10884 29573 10909 29629
rect 10965 29573 10990 29629
rect 11046 29573 11071 29629
rect 11127 29573 11152 29629
rect 10657 29549 11152 29573
rect 10657 29493 10666 29549
rect 10722 29493 10747 29549
rect 10803 29493 10828 29549
rect 10884 29493 10909 29549
rect 10965 29493 10990 29549
rect 11046 29493 11071 29549
rect 11127 29493 11152 29549
rect 10657 29469 11152 29493
rect 10657 29413 10666 29469
rect 10722 29413 10747 29469
rect 10803 29413 10828 29469
rect 10884 29413 10909 29469
rect 10965 29413 10990 29469
rect 11046 29413 11071 29469
rect 11127 29413 11152 29469
rect 10657 29389 11152 29413
rect 10657 29333 10666 29389
rect 10722 29333 10747 29389
rect 10803 29333 10828 29389
rect 10884 29333 10909 29389
rect 10965 29333 10990 29389
rect 11046 29333 11071 29389
rect 11127 29333 11152 29389
rect 10657 29309 11152 29333
rect 10657 29253 10666 29309
rect 10722 29253 10747 29309
rect 10803 29253 10828 29309
rect 10884 29253 10909 29309
rect 10965 29253 10990 29309
rect 11046 29253 11071 29309
rect 11127 29253 11152 29309
rect 10657 29229 11152 29253
rect 10657 29173 10666 29229
rect 10722 29173 10747 29229
rect 10803 29173 10828 29229
rect 10884 29173 10909 29229
rect 10965 29173 10990 29229
rect 11046 29173 11071 29229
rect 11127 29173 11152 29229
rect 10657 29149 11152 29173
rect 10657 29093 10666 29149
rect 10722 29093 10747 29149
rect 10803 29093 10828 29149
rect 10884 29093 10909 29149
rect 10965 29093 10990 29149
rect 11046 29093 11071 29149
rect 11127 29093 11152 29149
rect 10657 29069 11152 29093
rect 10657 29013 10666 29069
rect 10722 29013 10747 29069
rect 10803 29013 10828 29069
rect 10884 29013 10909 29069
rect 10965 29013 10990 29069
rect 11046 29013 11071 29069
rect 11127 29013 11152 29069
rect 10657 28989 11152 29013
rect 10657 28933 10666 28989
rect 10722 28933 10747 28989
rect 10803 28933 10828 28989
rect 10884 28933 10909 28989
rect 10965 28933 10990 28989
rect 11046 28933 11071 28989
rect 11127 28933 11152 28989
rect 10657 28909 11152 28933
rect 10657 28853 10666 28909
rect 10722 28853 10747 28909
rect 10803 28853 10828 28909
rect 10884 28853 10909 28909
rect 10965 28853 10990 28909
rect 11046 28853 11071 28909
rect 11127 28853 11152 28909
rect 10657 28829 11152 28853
rect 10657 28773 10666 28829
rect 10722 28773 10747 28829
rect 10803 28773 10828 28829
rect 10884 28773 10909 28829
rect 10965 28773 10990 28829
rect 11046 28773 11071 28829
rect 11127 28773 11152 28829
rect 10657 28749 11152 28773
rect 10657 28693 10666 28749
rect 10722 28693 10747 28749
rect 10803 28693 10828 28749
rect 10884 28693 10909 28749
rect 10965 28693 10990 28749
rect 11046 28693 11071 28749
rect 11127 28693 11152 28749
rect 10657 28669 11152 28693
rect 10657 28613 10666 28669
rect 10722 28613 10747 28669
rect 10803 28613 10828 28669
rect 10884 28613 10909 28669
rect 10965 28613 10990 28669
rect 11046 28613 11071 28669
rect 11127 28613 11152 28669
rect 10657 28589 11152 28613
rect 10657 28533 10666 28589
rect 10722 28533 10747 28589
rect 10803 28533 10828 28589
rect 10884 28533 10909 28589
rect 10965 28533 10990 28589
rect 11046 28533 11071 28589
rect 11127 28533 11152 28589
rect 10657 28509 11152 28533
rect 10657 28453 10666 28509
rect 10722 28453 10747 28509
rect 10803 28453 10828 28509
rect 10884 28453 10909 28509
rect 10965 28453 10990 28509
rect 11046 28453 11071 28509
rect 11127 28453 11152 28509
rect 10657 28429 11152 28453
rect 10657 28373 10666 28429
rect 10722 28373 10747 28429
rect 10803 28373 10828 28429
rect 10884 28373 10909 28429
rect 10965 28373 10990 28429
rect 11046 28373 11071 28429
rect 11127 28373 11152 28429
rect 10657 28349 11152 28373
rect 10657 28293 10666 28349
rect 10722 28293 10747 28349
rect 10803 28293 10828 28349
rect 10884 28293 10909 28349
rect 10965 28293 10990 28349
rect 11046 28293 11071 28349
rect 11127 28293 11152 28349
rect 10657 28269 11152 28293
rect 10657 28213 10666 28269
rect 10722 28213 10747 28269
rect 10803 28213 10828 28269
rect 10884 28213 10909 28269
rect 10965 28213 10990 28269
rect 11046 28213 11071 28269
rect 11127 28213 11152 28269
rect 10657 28189 11152 28213
rect 10657 28133 10666 28189
rect 10722 28133 10747 28189
rect 10803 28133 10828 28189
rect 10884 28133 10909 28189
rect 10965 28133 10990 28189
rect 11046 28133 11071 28189
rect 11127 28133 11152 28189
rect 10657 28109 11152 28133
rect 10657 28053 10666 28109
rect 10722 28053 10747 28109
rect 10803 28053 10828 28109
rect 10884 28053 10909 28109
rect 10965 28053 10990 28109
rect 11046 28053 11071 28109
rect 11127 28053 11152 28109
rect 10657 28029 11152 28053
rect 10657 27973 10666 28029
rect 10722 27973 10747 28029
rect 10803 27973 10828 28029
rect 10884 27973 10909 28029
rect 10965 27973 10990 28029
rect 11046 27973 11071 28029
rect 11127 27973 11152 28029
rect 10657 27949 11152 27973
rect 10657 27893 10666 27949
rect 10722 27893 10747 27949
rect 10803 27893 10828 27949
rect 10884 27893 10909 27949
rect 10965 27893 10990 27949
rect 11046 27893 11071 27949
rect 11127 27893 11152 27949
rect 11848 27893 11857 29629
rect 10657 25029 11857 27893
rect 10657 24973 10666 25029
rect 10722 24973 10747 25029
rect 10803 24973 10828 25029
rect 10884 24973 10909 25029
rect 10965 24973 10990 25029
rect 11046 24973 11071 25029
rect 11127 24973 11152 25029
rect 10657 24949 11152 24973
rect 10657 24893 10666 24949
rect 10722 24893 10747 24949
rect 10803 24893 10828 24949
rect 10884 24893 10909 24949
rect 10965 24893 10990 24949
rect 11046 24893 11071 24949
rect 11127 24893 11152 24949
rect 10657 24869 11152 24893
rect 10657 24813 10666 24869
rect 10722 24813 10747 24869
rect 10803 24813 10828 24869
rect 10884 24813 10909 24869
rect 10965 24813 10990 24869
rect 11046 24813 11071 24869
rect 11127 24813 11152 24869
rect 10657 24789 11152 24813
rect 10657 24733 10666 24789
rect 10722 24733 10747 24789
rect 10803 24733 10828 24789
rect 10884 24733 10909 24789
rect 10965 24733 10990 24789
rect 11046 24733 11071 24789
rect 11127 24733 11152 24789
rect 10657 24709 11152 24733
rect 10657 24653 10666 24709
rect 10722 24653 10747 24709
rect 10803 24653 10828 24709
rect 10884 24653 10909 24709
rect 10965 24653 10990 24709
rect 11046 24653 11071 24709
rect 11127 24653 11152 24709
rect 10657 24629 11152 24653
rect 10657 24573 10666 24629
rect 10722 24573 10747 24629
rect 10803 24573 10828 24629
rect 10884 24573 10909 24629
rect 10965 24573 10990 24629
rect 11046 24573 11071 24629
rect 11127 24573 11152 24629
rect 10657 24549 11152 24573
rect 10657 24493 10666 24549
rect 10722 24493 10747 24549
rect 10803 24493 10828 24549
rect 10884 24493 10909 24549
rect 10965 24493 10990 24549
rect 11046 24493 11071 24549
rect 11127 24493 11152 24549
rect 10657 24469 11152 24493
rect 10657 24413 10666 24469
rect 10722 24413 10747 24469
rect 10803 24413 10828 24469
rect 10884 24413 10909 24469
rect 10965 24413 10990 24469
rect 11046 24413 11071 24469
rect 11127 24413 11152 24469
rect 10657 24389 11152 24413
rect 10657 24333 10666 24389
rect 10722 24333 10747 24389
rect 10803 24333 10828 24389
rect 10884 24333 10909 24389
rect 10965 24333 10990 24389
rect 11046 24333 11071 24389
rect 11127 24333 11152 24389
rect 10657 24309 11152 24333
rect 10657 24253 10666 24309
rect 10722 24253 10747 24309
rect 10803 24253 10828 24309
rect 10884 24253 10909 24309
rect 10965 24253 10990 24309
rect 11046 24253 11071 24309
rect 11127 24253 11152 24309
rect 10657 24229 11152 24253
rect 10657 24173 10666 24229
rect 10722 24173 10747 24229
rect 10803 24173 10828 24229
rect 10884 24173 10909 24229
rect 10965 24173 10990 24229
rect 11046 24173 11071 24229
rect 11127 24173 11152 24229
rect 10657 24149 11152 24173
rect 10657 24093 10666 24149
rect 10722 24093 10747 24149
rect 10803 24093 10828 24149
rect 10884 24093 10909 24149
rect 10965 24093 10990 24149
rect 11046 24093 11071 24149
rect 11127 24093 11152 24149
rect 10657 24069 11152 24093
rect 10657 24013 10666 24069
rect 10722 24013 10747 24069
rect 10803 24013 10828 24069
rect 10884 24013 10909 24069
rect 10965 24013 10990 24069
rect 11046 24013 11071 24069
rect 11127 24013 11152 24069
rect 10657 23989 11152 24013
rect 10657 23933 10666 23989
rect 10722 23933 10747 23989
rect 10803 23933 10828 23989
rect 10884 23933 10909 23989
rect 10965 23933 10990 23989
rect 11046 23933 11071 23989
rect 11127 23933 11152 23989
rect 10657 23909 11152 23933
rect 10657 23853 10666 23909
rect 10722 23853 10747 23909
rect 10803 23853 10828 23909
rect 10884 23853 10909 23909
rect 10965 23853 10990 23909
rect 11046 23853 11071 23909
rect 11127 23853 11152 23909
rect 10657 23829 11152 23853
rect 10657 23773 10666 23829
rect 10722 23773 10747 23829
rect 10803 23773 10828 23829
rect 10884 23773 10909 23829
rect 10965 23773 10990 23829
rect 11046 23773 11071 23829
rect 11127 23773 11152 23829
rect 10657 23749 11152 23773
rect 10657 23693 10666 23749
rect 10722 23693 10747 23749
rect 10803 23693 10828 23749
rect 10884 23693 10909 23749
rect 10965 23693 10990 23749
rect 11046 23693 11071 23749
rect 11127 23693 11152 23749
rect 10657 23669 11152 23693
rect 10657 23613 10666 23669
rect 10722 23613 10747 23669
rect 10803 23613 10828 23669
rect 10884 23613 10909 23669
rect 10965 23613 10990 23669
rect 11046 23613 11071 23669
rect 11127 23613 11152 23669
rect 10657 23589 11152 23613
rect 10657 23533 10666 23589
rect 10722 23533 10747 23589
rect 10803 23533 10828 23589
rect 10884 23533 10909 23589
rect 10965 23533 10990 23589
rect 11046 23533 11071 23589
rect 11127 23533 11152 23589
rect 10657 23509 11152 23533
rect 10657 23453 10666 23509
rect 10722 23453 10747 23509
rect 10803 23453 10828 23509
rect 10884 23453 10909 23509
rect 10965 23453 10990 23509
rect 11046 23453 11071 23509
rect 11127 23453 11152 23509
rect 10657 23429 11152 23453
rect 10657 23373 10666 23429
rect 10722 23373 10747 23429
rect 10803 23373 10828 23429
rect 10884 23373 10909 23429
rect 10965 23373 10990 23429
rect 11046 23373 11071 23429
rect 11127 23373 11152 23429
rect 10657 23349 11152 23373
rect 10657 23293 10666 23349
rect 10722 23293 10747 23349
rect 10803 23293 10828 23349
rect 10884 23293 10909 23349
rect 10965 23293 10990 23349
rect 11046 23293 11071 23349
rect 11127 23293 11152 23349
rect 11848 23293 11857 25029
tri 8077 21630 8535 22088 se
rect 8535 21630 9771 22088
tri 10199 21630 10657 22088 se
rect 10657 21630 11857 23293
tri 7578 21131 8077 21630 se
rect 8077 21202 9343 21630
tri 9343 21202 9771 21630 nw
tri 9771 21202 10199 21630 se
rect 10199 21592 11857 21630
rect 10199 21202 10766 21592
rect 8077 21131 9113 21202
rect 7578 20972 9113 21131
tri 9113 20972 9343 21202 nw
tri 9541 20972 9771 21202 se
rect 9771 20972 10766 21202
rect 3100 20478 4478 20758
tri 4478 20478 4758 20758 sw
rect 5186 20478 6386 20758
rect 3100 20440 4758 20478
tri 3100 20429 3111 20440 ne
rect 3111 20429 4758 20440
tri 4758 20429 4807 20478 sw
tri 5186 20429 5235 20478 ne
rect 5235 20429 6386 20478
tri 6386 20429 6929 20972 sw
rect 7578 20929 9070 20972
tri 9070 20929 9113 20972 nw
tri 9498 20929 9541 20972 se
rect 9541 20929 10766 20972
rect 7578 20501 8642 20929
tri 8642 20501 9070 20929 nw
tri 9070 20501 9498 20929 se
rect 9498 20501 10766 20929
tri 10766 20501 11857 21592 nw
rect 7578 20429 8570 20501
tri 8570 20429 8642 20501 nw
rect 9070 20429 10692 20501
tri 3111 20373 3167 20429 ne
rect 3167 20373 4807 20429
tri 4807 20373 4863 20429 sw
tri 5235 20373 5291 20429 ne
rect 5291 20373 6929 20429
tri 6929 20373 6985 20429 sw
rect 7578 20373 7640 20429
rect 7696 20373 7726 20429
rect 7782 20373 7812 20429
rect 7868 20373 7898 20429
rect 7954 20373 7984 20429
rect 8040 20373 8070 20429
rect 8126 20373 8156 20429
rect 8212 20373 8242 20429
rect 8298 20373 8327 20429
rect 8383 20373 8412 20429
rect 8468 20373 8497 20429
rect 8553 20373 8568 20429
tri 8568 20427 8570 20429 nw
tri 3167 20349 3191 20373 ne
rect 3191 20349 4863 20373
tri 4863 20349 4887 20373 sw
tri 5291 20349 5315 20373 ne
rect 5315 20349 6985 20373
tri 6985 20349 7009 20373 sw
rect 7578 20349 8568 20373
tri 3191 20293 3247 20349 ne
rect 3247 20293 4887 20349
tri 4887 20293 4943 20349 sw
tri 5315 20293 5371 20349 ne
rect 5371 20293 7009 20349
tri 7009 20293 7065 20349 sw
rect 7578 20293 7640 20349
rect 7696 20293 7726 20349
rect 7782 20293 7812 20349
rect 7868 20293 7898 20349
rect 7954 20293 7984 20349
rect 8040 20293 8070 20349
rect 8126 20293 8156 20349
rect 8212 20293 8242 20349
rect 8298 20293 8327 20349
rect 8383 20293 8412 20349
rect 8468 20293 8497 20349
rect 8553 20293 8568 20349
tri 3247 20269 3271 20293 ne
rect 3271 20269 4943 20293
tri 4943 20269 4967 20293 sw
tri 5371 20269 5395 20293 ne
rect 5395 20269 7065 20293
tri 7065 20269 7089 20293 sw
rect 7578 20269 8568 20293
tri 3271 20213 3327 20269 ne
rect 3327 20213 4967 20269
tri 4967 20213 5023 20269 sw
tri 5395 20213 5451 20269 ne
rect 5451 20213 7089 20269
tri 7089 20213 7145 20269 sw
rect 7578 20213 7640 20269
rect 7696 20213 7726 20269
rect 7782 20213 7812 20269
rect 7868 20213 7898 20269
rect 7954 20213 7984 20269
rect 8040 20213 8070 20269
rect 8126 20213 8156 20269
rect 8212 20213 8242 20269
rect 8298 20213 8327 20269
rect 8383 20213 8412 20269
rect 8468 20213 8497 20269
rect 8553 20213 8568 20269
tri 3327 20189 3351 20213 ne
rect 3351 20189 5023 20213
tri 5023 20189 5047 20213 sw
tri 5451 20189 5475 20213 ne
rect 5475 20189 7145 20213
tri 7145 20189 7169 20213 sw
rect 7578 20189 8568 20213
tri 3351 20133 3407 20189 ne
rect 3407 20133 5047 20189
tri 5047 20133 5103 20189 sw
tri 5475 20133 5531 20189 ne
rect 5531 20133 7169 20189
tri 7169 20133 7225 20189 sw
rect 7578 20133 7640 20189
rect 7696 20133 7726 20189
rect 7782 20133 7812 20189
rect 7868 20133 7898 20189
rect 7954 20133 7984 20189
rect 8040 20133 8070 20189
rect 8126 20133 8156 20189
rect 8212 20133 8242 20189
rect 8298 20133 8327 20189
rect 8383 20133 8412 20189
rect 8468 20133 8497 20189
rect 8553 20133 8568 20189
tri 3407 20109 3431 20133 ne
rect 3431 20109 5103 20133
tri 5103 20109 5127 20133 sw
tri 5531 20109 5555 20133 ne
rect 5555 20109 7225 20133
tri 7225 20109 7249 20133 sw
rect 7578 20109 8568 20133
tri 3431 20053 3487 20109 ne
rect 3487 20053 5127 20109
tri 5127 20053 5183 20109 sw
tri 5555 20053 5611 20109 ne
rect 5611 20053 7249 20109
tri 7249 20053 7305 20109 sw
rect 7578 20053 7640 20109
rect 7696 20053 7726 20109
rect 7782 20053 7812 20109
rect 7868 20053 7898 20109
rect 7954 20053 7984 20109
rect 8040 20053 8070 20109
rect 8126 20053 8156 20109
rect 8212 20053 8242 20109
rect 8298 20053 8327 20109
rect 8383 20053 8412 20109
rect 8468 20053 8497 20109
rect 8553 20053 8568 20109
rect 9070 20373 9079 20429
rect 9135 20373 9170 20429
rect 9226 20373 9260 20429
rect 9316 20373 9350 20429
rect 9406 20373 9440 20429
rect 9496 20373 9530 20429
rect 9586 20373 9620 20429
rect 9676 20373 9710 20429
rect 9766 20427 10692 20429
tri 10692 20427 10766 20501 nw
rect 9766 20373 10322 20427
rect 9070 20349 10322 20373
rect 9070 20293 9079 20349
rect 9135 20293 9170 20349
rect 9226 20293 9260 20349
rect 9316 20293 9350 20349
rect 9406 20293 9440 20349
rect 9496 20293 9530 20349
rect 9586 20293 9620 20349
rect 9676 20293 9710 20349
rect 9766 20293 10322 20349
rect 9070 20269 10322 20293
rect 9070 20213 9079 20269
rect 9135 20213 9170 20269
rect 9226 20213 9260 20269
rect 9316 20213 9350 20269
rect 9406 20213 9440 20269
rect 9496 20213 9530 20269
rect 9586 20213 9620 20269
rect 9676 20213 9710 20269
rect 9766 20213 10322 20269
rect 9070 20189 10322 20213
rect 9070 20133 9079 20189
rect 9135 20133 9170 20189
rect 9226 20133 9260 20189
rect 9316 20133 9350 20189
rect 9406 20133 9440 20189
rect 9496 20133 9530 20189
rect 9586 20133 9620 20189
rect 9676 20133 9710 20189
rect 9766 20133 10322 20189
rect 9070 20109 10322 20133
tri 8568 20053 8572 20057 sw
rect 9070 20053 9079 20109
rect 9135 20053 9170 20109
rect 9226 20053 9260 20109
rect 9316 20053 9350 20109
rect 9406 20053 9440 20109
rect 9496 20053 9530 20109
rect 9586 20053 9620 20109
rect 9676 20053 9710 20109
rect 9766 20057 10322 20109
tri 10322 20057 10692 20427 nw
rect 9766 20053 10311 20057
tri 3487 20050 3490 20053 ne
rect 3490 20050 5183 20053
tri 5183 20050 5186 20053 sw
tri 5611 20050 5614 20053 ne
rect 5614 20050 7305 20053
tri 3490 20029 3511 20050 ne
rect 3511 20029 5186 20050
tri 5186 20029 5207 20050 sw
tri 5614 20029 5635 20050 ne
rect 5635 20029 7305 20050
tri 7305 20029 7329 20053 sw
rect 7578 20046 8572 20053
tri 8572 20046 8579 20053 sw
rect 9070 20046 10311 20053
tri 10311 20046 10322 20057 nw
rect 7578 20029 8579 20046
tri 8579 20029 8596 20046 sw
tri 9053 20029 9070 20046 se
rect 9070 20029 10208 20046
tri 3511 19973 3567 20029 ne
rect 3567 19979 5207 20029
tri 5207 19979 5257 20029 sw
tri 5635 19979 5685 20029 ne
rect 5685 19979 7329 20029
tri 7329 19979 7379 20029 sw
rect 3567 19973 5257 19979
tri 5257 19973 5263 19979 sw
tri 5685 19973 5691 19979 ne
rect 5691 19973 7379 19979
tri 3567 19949 3591 19973 ne
rect 3591 19949 5263 19973
tri 5263 19949 5287 19973 sw
tri 5691 19949 5715 19973 ne
rect 5715 19949 7379 19973
tri 3591 19893 3647 19949 ne
rect 3647 19893 5287 19949
tri 5287 19893 5343 19949 sw
tri 5715 19893 5771 19949 ne
rect 5771 19893 7379 19949
tri 3647 19869 3671 19893 ne
rect 3671 19869 5343 19893
tri 5343 19869 5367 19893 sw
tri 5771 19869 5795 19893 ne
rect 5795 19869 7379 19893
tri 3671 19813 3727 19869 ne
rect 3727 19813 5367 19869
tri 5367 19813 5423 19869 sw
tri 5795 19813 5851 19869 ne
rect 5851 19813 7379 19869
tri 3727 19789 3751 19813 ne
rect 3751 19789 5423 19813
tri 5423 19789 5447 19813 sw
tri 5851 19789 5875 19813 ne
rect 5875 19789 7379 19813
tri 3751 19733 3807 19789 ne
rect 3807 19759 5447 19789
tri 5447 19759 5477 19789 sw
tri 5875 19759 5905 19789 ne
rect 5905 19759 7379 19789
rect 3807 19733 5477 19759
tri 5477 19733 5503 19759 sw
tri 5905 19733 5931 19759 ne
rect 5931 19733 7379 19759
tri 3807 19709 3831 19733 ne
rect 3831 19709 5503 19733
tri 5503 19709 5527 19733 sw
tri 5931 19709 5955 19733 ne
rect 5955 19709 7379 19733
tri 3831 19653 3887 19709 ne
rect 3887 19653 5527 19709
tri 5527 19653 5583 19709 sw
tri 5955 19653 6011 19709 ne
rect 6011 19653 7379 19709
tri 3887 19629 3911 19653 ne
rect 3911 19629 5583 19653
tri 5583 19629 5607 19653 sw
tri 6011 19629 6035 19653 ne
rect 6035 19629 7379 19653
tri 3911 19573 3967 19629 ne
rect 3967 19573 5607 19629
tri 5607 19573 5663 19629 sw
tri 6035 19573 6091 19629 ne
rect 6091 19573 7379 19629
tri 3967 19549 3991 19573 ne
rect 3991 19549 5663 19573
tri 5663 19549 5687 19573 sw
tri 6091 19549 6115 19573 ne
rect 6115 19549 7379 19573
tri 3991 19493 4047 19549 ne
rect 4047 19493 5687 19549
tri 5687 19493 5743 19549 sw
tri 6115 19493 6171 19549 ne
rect 6171 19493 7379 19549
tri 4047 19469 4071 19493 ne
rect 4071 19469 5743 19493
tri 5743 19469 5767 19493 sw
tri 6171 19469 6195 19493 ne
rect 6195 19469 7379 19493
tri 4071 19413 4127 19469 ne
rect 4127 19413 5767 19469
tri 5767 19413 5823 19469 sw
tri 6195 19413 6251 19469 ne
rect 6251 19413 7379 19469
tri 4127 19389 4151 19413 ne
rect 4151 19389 5823 19413
tri 5823 19389 5847 19413 sw
tri 6251 19389 6275 19413 ne
rect 6275 19389 7379 19413
tri 4151 19333 4207 19389 ne
rect 4207 19333 5847 19389
tri 5847 19333 5903 19389 sw
tri 6275 19333 6331 19389 ne
rect 6331 19333 7379 19389
tri 4207 19331 4209 19333 ne
rect 4209 19331 5903 19333
tri 5903 19331 5905 19333 sw
tri 6331 19331 6333 19333 ne
rect 6333 19331 7379 19333
tri 4209 19309 4231 19331 ne
rect 4231 19309 5905 19331
tri 6333 19309 6355 19331 ne
rect 6355 19309 7379 19331
tri 4231 19278 4262 19309 ne
rect 4262 19278 5905 19309
tri 6355 19278 6386 19309 ne
rect 6386 19278 7379 19309
tri 4262 19275 4265 19278 ne
rect 4265 19275 5905 19278
tri 6386 19275 6389 19278 ne
tri 4265 19253 4287 19275 ne
rect 4287 19253 5905 19275
tri 4287 19240 4300 19253 ne
rect 4300 19240 5905 19253
tri 4300 19229 4311 19240 ne
rect 4311 19229 5905 19240
tri 4311 19173 4367 19229 ne
rect 4367 19173 5905 19229
tri 4367 19149 4391 19173 ne
rect 4391 19149 5905 19173
tri 4391 19093 4447 19149 ne
rect 4447 19093 5905 19149
tri 4447 19069 4471 19093 ne
rect 4471 19069 5905 19093
tri 4471 19013 4527 19069 ne
rect 4527 19013 5905 19069
tri 4527 18989 4551 19013 ne
rect 4551 18989 5905 19013
tri 4551 18933 4607 18989 ne
rect 4607 18933 5905 18989
tri 4607 18909 4631 18933 ne
rect 4631 18909 5905 18933
tri 4631 18853 4687 18909 ne
rect 4687 18853 5905 18909
tri 4687 18829 4711 18853 ne
rect 4711 18829 5905 18853
tri 4711 18791 4749 18829 ne
rect 4749 18508 5905 18829
tri 4749 18478 4779 18508 ne
rect 4779 18478 5905 18508
tri 5905 18478 6047 18620 sw
tri 6247 18478 6389 18620 se
rect 6389 18478 7379 19278
tri 4779 18078 5179 18478 ne
rect 5179 17894 7379 18478
rect 5179 17838 5188 17894
rect 5244 17838 5270 17894
rect 5326 17838 5352 17894
rect 5408 17838 5434 17894
rect 5490 17838 5516 17894
rect 5572 17838 5598 17894
rect 5654 17838 5680 17894
rect 5736 17838 5762 17894
rect 5818 17838 5844 17894
rect 5900 17838 5926 17894
rect 5982 17838 6008 17894
rect 6064 17838 6090 17894
rect 6146 17838 6172 17894
rect 6228 17838 6254 17894
rect 6310 17838 6336 17894
rect 6392 17838 6418 17894
rect 6474 17838 6500 17894
rect 6556 17838 6582 17894
rect 6638 17838 6664 17894
rect 6720 17838 6746 17894
rect 6802 17838 6828 17894
rect 6884 17838 6909 17894
rect 6965 17838 6990 17894
rect 7046 17838 7071 17894
rect 7127 17838 7152 17894
rect 7208 17838 7233 17894
rect 7289 17838 7314 17894
rect 7370 17838 7379 17894
rect 5179 17814 7379 17838
rect 5179 17758 5188 17814
rect 5244 17758 5270 17814
rect 5326 17758 5352 17814
rect 5408 17758 5434 17814
rect 5490 17758 5516 17814
rect 5572 17758 5598 17814
rect 5654 17758 5680 17814
rect 5736 17758 5762 17814
rect 5818 17758 5844 17814
rect 5900 17758 5926 17814
rect 5982 17758 6008 17814
rect 6064 17758 6090 17814
rect 6146 17758 6172 17814
rect 6228 17758 6254 17814
rect 6310 17758 6336 17814
rect 6392 17758 6418 17814
rect 6474 17758 6500 17814
rect 6556 17758 6582 17814
rect 6638 17758 6664 17814
rect 6720 17758 6746 17814
rect 6802 17758 6828 17814
rect 6884 17758 6909 17814
rect 6965 17758 6990 17814
rect 7046 17758 7071 17814
rect 7127 17758 7152 17814
rect 7208 17758 7233 17814
rect 7289 17758 7314 17814
rect 7370 17758 7379 17814
rect 5179 17734 7379 17758
rect 5179 17678 5188 17734
rect 5244 17678 5270 17734
rect 5326 17678 5352 17734
rect 5408 17678 5434 17734
rect 5490 17678 5516 17734
rect 5572 17678 5598 17734
rect 5654 17678 5680 17734
rect 5736 17678 5762 17734
rect 5818 17678 5844 17734
rect 5900 17678 5926 17734
rect 5982 17678 6008 17734
rect 6064 17678 6090 17734
rect 6146 17678 6172 17734
rect 6228 17678 6254 17734
rect 6310 17678 6336 17734
rect 6392 17678 6418 17734
rect 6474 17678 6500 17734
rect 6556 17678 6582 17734
rect 6638 17678 6664 17734
rect 6720 17678 6746 17734
rect 6802 17678 6828 17734
rect 6884 17678 6909 17734
rect 6965 17678 6990 17734
rect 7046 17678 7071 17734
rect 7127 17678 7152 17734
rect 7208 17678 7233 17734
rect 7289 17678 7314 17734
rect 7370 17678 7379 17734
rect 5179 17654 7379 17678
rect 5179 17598 5188 17654
rect 5244 17598 5270 17654
rect 5326 17598 5352 17654
rect 5408 17598 5434 17654
rect 5490 17598 5516 17654
rect 5572 17598 5598 17654
rect 5654 17598 5680 17654
rect 5736 17598 5762 17654
rect 5818 17598 5844 17654
rect 5900 17598 5926 17654
rect 5982 17598 6008 17654
rect 6064 17598 6090 17654
rect 6146 17598 6172 17654
rect 6228 17598 6254 17654
rect 6310 17598 6336 17654
rect 6392 17598 6418 17654
rect 6474 17598 6500 17654
rect 6556 17598 6582 17654
rect 6638 17598 6664 17654
rect 6720 17598 6746 17654
rect 6802 17598 6828 17654
rect 6884 17598 6909 17654
rect 6965 17598 6990 17654
rect 7046 17598 7071 17654
rect 7127 17598 7152 17654
rect 7208 17598 7233 17654
rect 7289 17598 7314 17654
rect 7370 17598 7379 17654
rect 5179 17574 7379 17598
rect 5179 17518 5188 17574
rect 5244 17518 5270 17574
rect 5326 17518 5352 17574
rect 5408 17518 5434 17574
rect 5490 17518 5516 17574
rect 5572 17518 5598 17574
rect 5654 17518 5680 17574
rect 5736 17518 5762 17574
rect 5818 17518 5844 17574
rect 5900 17518 5926 17574
rect 5982 17518 6008 17574
rect 6064 17518 6090 17574
rect 6146 17518 6172 17574
rect 6228 17518 6254 17574
rect 6310 17518 6336 17574
rect 6392 17518 6418 17574
rect 6474 17518 6500 17574
rect 6556 17518 6582 17574
rect 6638 17518 6664 17574
rect 6720 17518 6746 17574
rect 6802 17518 6828 17574
rect 6884 17518 6909 17574
rect 6965 17518 6990 17574
rect 7046 17518 7071 17574
rect 7127 17518 7152 17574
rect 7208 17518 7233 17574
rect 7289 17518 7314 17574
rect 7370 17518 7379 17574
rect 5179 17494 7379 17518
rect 5179 17438 5188 17494
rect 5244 17438 5270 17494
rect 5326 17438 5352 17494
rect 5408 17438 5434 17494
rect 5490 17438 5516 17494
rect 5572 17438 5598 17494
rect 5654 17438 5680 17494
rect 5736 17438 5762 17494
rect 5818 17438 5844 17494
rect 5900 17438 5926 17494
rect 5982 17438 6008 17494
rect 6064 17438 6090 17494
rect 6146 17438 6172 17494
rect 6228 17438 6254 17494
rect 6310 17438 6336 17494
rect 6392 17438 6418 17494
rect 6474 17438 6500 17494
rect 6556 17438 6582 17494
rect 6638 17438 6664 17494
rect 6720 17438 6746 17494
rect 6802 17438 6828 17494
rect 6884 17438 6909 17494
rect 6965 17438 6990 17494
rect 7046 17438 7071 17494
rect 7127 17438 7152 17494
rect 7208 17438 7233 17494
rect 7289 17438 7314 17494
rect 7370 17438 7379 17494
rect 5179 17414 7379 17438
rect 5179 17358 5188 17414
rect 5244 17358 5270 17414
rect 5326 17358 5352 17414
rect 5408 17358 5434 17414
rect 5490 17358 5516 17414
rect 5572 17358 5598 17414
rect 5654 17358 5680 17414
rect 5736 17358 5762 17414
rect 5818 17358 5844 17414
rect 5900 17358 5926 17414
rect 5982 17358 6008 17414
rect 6064 17358 6090 17414
rect 6146 17358 6172 17414
rect 6228 17358 6254 17414
rect 6310 17358 6336 17414
rect 6392 17358 6418 17414
rect 6474 17358 6500 17414
rect 6556 17358 6582 17414
rect 6638 17358 6664 17414
rect 6720 17358 6746 17414
rect 6802 17358 6828 17414
rect 6884 17358 6909 17414
rect 6965 17358 6990 17414
rect 7046 17358 7071 17414
rect 7127 17358 7152 17414
rect 7208 17358 7233 17414
rect 7289 17358 7314 17414
rect 7370 17358 7379 17414
rect 5179 17334 7379 17358
rect 5179 17278 5188 17334
rect 5244 17278 5270 17334
rect 5326 17278 5352 17334
rect 5408 17278 5434 17334
rect 5490 17278 5516 17334
rect 5572 17278 5598 17334
rect 5654 17278 5680 17334
rect 5736 17278 5762 17334
rect 5818 17278 5844 17334
rect 5900 17278 5926 17334
rect 5982 17278 6008 17334
rect 6064 17278 6090 17334
rect 6146 17278 6172 17334
rect 6228 17278 6254 17334
rect 6310 17278 6336 17334
rect 6392 17278 6418 17334
rect 6474 17278 6500 17334
rect 6556 17278 6582 17334
rect 6638 17278 6664 17334
rect 6720 17278 6746 17334
rect 6802 17278 6828 17334
rect 6884 17278 6909 17334
rect 6965 17278 6990 17334
rect 7046 17278 7071 17334
rect 7127 17278 7152 17334
rect 7208 17278 7233 17334
rect 7289 17278 7314 17334
rect 7370 17278 7379 17334
rect 5179 17254 7379 17278
rect 5179 17198 5188 17254
rect 5244 17198 5270 17254
rect 5326 17198 5352 17254
rect 5408 17198 5434 17254
rect 5490 17198 5516 17254
rect 5572 17198 5598 17254
rect 5654 17198 5680 17254
rect 5736 17198 5762 17254
rect 5818 17198 5844 17254
rect 5900 17198 5926 17254
rect 5982 17198 6008 17254
rect 6064 17198 6090 17254
rect 6146 17198 6172 17254
rect 6228 17198 6254 17254
rect 6310 17198 6336 17254
rect 6392 17198 6418 17254
rect 6474 17198 6500 17254
rect 6556 17198 6582 17254
rect 6638 17198 6664 17254
rect 6720 17198 6746 17254
rect 6802 17198 6828 17254
rect 6884 17198 6909 17254
rect 6965 17198 6990 17254
rect 7046 17198 7071 17254
rect 7127 17198 7152 17254
rect 7208 17198 7233 17254
rect 7289 17198 7314 17254
rect 7370 17198 7379 17254
rect 5179 17174 7379 17198
rect 5179 17118 5188 17174
rect 5244 17118 5270 17174
rect 5326 17118 5352 17174
rect 5408 17118 5434 17174
rect 5490 17118 5516 17174
rect 5572 17118 5598 17174
rect 5654 17118 5680 17174
rect 5736 17118 5762 17174
rect 5818 17118 5844 17174
rect 5900 17118 5926 17174
rect 5982 17118 6008 17174
rect 6064 17118 6090 17174
rect 6146 17118 6172 17174
rect 6228 17118 6254 17174
rect 6310 17118 6336 17174
rect 6392 17118 6418 17174
rect 6474 17118 6500 17174
rect 6556 17118 6582 17174
rect 6638 17118 6664 17174
rect 6720 17118 6746 17174
rect 6802 17118 6828 17174
rect 6884 17118 6909 17174
rect 6965 17118 6990 17174
rect 7046 17118 7071 17174
rect 7127 17118 7152 17174
rect 7208 17118 7233 17174
rect 7289 17118 7314 17174
rect 7370 17118 7379 17174
rect 5179 17094 7379 17118
rect 5179 17038 5188 17094
rect 5244 17038 5270 17094
rect 5326 17038 5352 17094
rect 5408 17038 5434 17094
rect 5490 17038 5516 17094
rect 5572 17038 5598 17094
rect 5654 17038 5680 17094
rect 5736 17038 5762 17094
rect 5818 17038 5844 17094
rect 5900 17038 5926 17094
rect 5982 17038 6008 17094
rect 6064 17038 6090 17094
rect 6146 17038 6172 17094
rect 6228 17038 6254 17094
rect 6310 17038 6336 17094
rect 6392 17038 6418 17094
rect 6474 17038 6500 17094
rect 6556 17038 6582 17094
rect 6638 17038 6664 17094
rect 6720 17038 6746 17094
rect 6802 17038 6828 17094
rect 6884 17038 6909 17094
rect 6965 17038 6990 17094
rect 7046 17038 7071 17094
rect 7127 17038 7152 17094
rect 7208 17038 7233 17094
rect 7289 17038 7314 17094
rect 7370 17038 7379 17094
rect 5179 17014 7379 17038
rect 5179 16958 5188 17014
rect 5244 16958 5270 17014
rect 5326 16958 5352 17014
rect 5408 16958 5434 17014
rect 5490 16958 5516 17014
rect 5572 16958 5598 17014
rect 5654 16958 5680 17014
rect 5736 16958 5762 17014
rect 5818 16958 5844 17014
rect 5900 16958 5926 17014
rect 5982 16958 6008 17014
rect 6064 16958 6090 17014
rect 6146 16958 6172 17014
rect 6228 16958 6254 17014
rect 6310 16958 6336 17014
rect 6392 16958 6418 17014
rect 6474 16958 6500 17014
rect 6556 16958 6582 17014
rect 6638 16958 6664 17014
rect 6720 16958 6746 17014
rect 6802 16958 6828 17014
rect 6884 16958 6909 17014
rect 6965 16958 6990 17014
rect 7046 16958 7071 17014
rect 7127 16958 7152 17014
rect 7208 16958 7233 17014
rect 7289 16958 7314 17014
rect 7370 16958 7379 17014
rect 5179 16934 7379 16958
rect 5179 16878 5188 16934
rect 5244 16878 5270 16934
rect 5326 16878 5352 16934
rect 5408 16878 5434 16934
rect 5490 16878 5516 16934
rect 5572 16878 5598 16934
rect 5654 16878 5680 16934
rect 5736 16878 5762 16934
rect 5818 16878 5844 16934
rect 5900 16878 5926 16934
rect 5982 16878 6008 16934
rect 6064 16878 6090 16934
rect 6146 16878 6172 16934
rect 6228 16878 6254 16934
rect 6310 16878 6336 16934
rect 6392 16878 6418 16934
rect 6474 16878 6500 16934
rect 6556 16878 6582 16934
rect 6638 16878 6664 16934
rect 6720 16878 6746 16934
rect 6802 16878 6828 16934
rect 6884 16878 6909 16934
rect 6965 16878 6990 16934
rect 7046 16878 7071 16934
rect 7127 16878 7152 16934
rect 7208 16878 7233 16934
rect 7289 16878 7314 16934
rect 7370 16878 7379 16934
rect 5179 16854 7379 16878
rect 5179 16798 5188 16854
rect 5244 16798 5270 16854
rect 5326 16798 5352 16854
rect 5408 16798 5434 16854
rect 5490 16798 5516 16854
rect 5572 16798 5598 16854
rect 5654 16798 5680 16854
rect 5736 16798 5762 16854
rect 5818 16798 5844 16854
rect 5900 16798 5926 16854
rect 5982 16798 6008 16854
rect 6064 16798 6090 16854
rect 6146 16798 6172 16854
rect 6228 16798 6254 16854
rect 6310 16798 6336 16854
rect 6392 16798 6418 16854
rect 6474 16798 6500 16854
rect 6556 16798 6582 16854
rect 6638 16798 6664 16854
rect 6720 16798 6746 16854
rect 6802 16798 6828 16854
rect 6884 16798 6909 16854
rect 6965 16798 6990 16854
rect 7046 16798 7071 16854
rect 7127 16798 7152 16854
rect 7208 16798 7233 16854
rect 7289 16798 7314 16854
rect 7370 16798 7379 16854
rect 5179 16774 7379 16798
rect 5179 16718 5188 16774
rect 5244 16718 5270 16774
rect 5326 16718 5352 16774
rect 5408 16718 5434 16774
rect 5490 16718 5516 16774
rect 5572 16718 5598 16774
rect 5654 16718 5680 16774
rect 5736 16718 5762 16774
rect 5818 16718 5844 16774
rect 5900 16718 5926 16774
rect 5982 16718 6008 16774
rect 6064 16718 6090 16774
rect 6146 16718 6172 16774
rect 6228 16718 6254 16774
rect 6310 16718 6336 16774
rect 6392 16718 6418 16774
rect 6474 16718 6500 16774
rect 6556 16718 6582 16774
rect 6638 16718 6664 16774
rect 6720 16718 6746 16774
rect 6802 16718 6828 16774
rect 6884 16718 6909 16774
rect 6965 16718 6990 16774
rect 7046 16718 7071 16774
rect 7127 16718 7152 16774
rect 7208 16718 7233 16774
rect 7289 16718 7314 16774
rect 7370 16718 7379 16774
rect 5179 16694 7379 16718
rect 5179 16638 5188 16694
rect 5244 16638 5270 16694
rect 5326 16638 5352 16694
rect 5408 16638 5434 16694
rect 5490 16638 5516 16694
rect 5572 16638 5598 16694
rect 5654 16638 5680 16694
rect 5736 16638 5762 16694
rect 5818 16638 5844 16694
rect 5900 16638 5926 16694
rect 5982 16638 6008 16694
rect 6064 16638 6090 16694
rect 6146 16638 6172 16694
rect 6228 16638 6254 16694
rect 6310 16638 6336 16694
rect 6392 16638 6418 16694
rect 6474 16638 6500 16694
rect 6556 16638 6582 16694
rect 6638 16638 6664 16694
rect 6720 16638 6746 16694
rect 6802 16638 6828 16694
rect 6884 16638 6909 16694
rect 6965 16638 6990 16694
rect 7046 16638 7071 16694
rect 7127 16638 7152 16694
rect 7208 16638 7233 16694
rect 7289 16638 7314 16694
rect 7370 16638 7379 16694
rect 5179 16614 7379 16638
rect 5179 16558 5188 16614
rect 5244 16558 5270 16614
rect 5326 16558 5352 16614
rect 5408 16558 5434 16614
rect 5490 16558 5516 16614
rect 5572 16558 5598 16614
rect 5654 16558 5680 16614
rect 5736 16558 5762 16614
rect 5818 16558 5844 16614
rect 5900 16558 5926 16614
rect 5982 16558 6008 16614
rect 6064 16558 6090 16614
rect 6146 16558 6172 16614
rect 6228 16558 6254 16614
rect 6310 16558 6336 16614
rect 6392 16558 6418 16614
rect 6474 16558 6500 16614
rect 6556 16558 6582 16614
rect 6638 16558 6664 16614
rect 6720 16558 6746 16614
rect 6802 16558 6828 16614
rect 6884 16558 6909 16614
rect 6965 16558 6990 16614
rect 7046 16558 7071 16614
rect 7127 16558 7152 16614
rect 7208 16558 7233 16614
rect 7289 16558 7314 16614
rect 7370 16558 7379 16614
rect 5179 16534 7379 16558
rect 5179 16478 5188 16534
rect 5244 16478 5270 16534
rect 5326 16478 5352 16534
rect 5408 16478 5434 16534
rect 5490 16478 5516 16534
rect 5572 16478 5598 16534
rect 5654 16478 5680 16534
rect 5736 16478 5762 16534
rect 5818 16478 5844 16534
rect 5900 16478 5926 16534
rect 5982 16478 6008 16534
rect 6064 16478 6090 16534
rect 6146 16478 6172 16534
rect 6228 16478 6254 16534
rect 6310 16478 6336 16534
rect 6392 16478 6418 16534
rect 6474 16478 6500 16534
rect 6556 16478 6582 16534
rect 6638 16478 6664 16534
rect 6720 16478 6746 16534
rect 6802 16478 6828 16534
rect 6884 16478 6909 16534
rect 6965 16478 6990 16534
rect 7046 16478 7071 16534
rect 7127 16478 7152 16534
rect 7208 16478 7233 16534
rect 7289 16478 7314 16534
rect 7370 16478 7379 16534
rect 5179 16454 7379 16478
rect 5179 16398 5188 16454
rect 5244 16398 5270 16454
rect 5326 16398 5352 16454
rect 5408 16398 5434 16454
rect 5490 16398 5516 16454
rect 5572 16398 5598 16454
rect 5654 16398 5680 16454
rect 5736 16398 5762 16454
rect 5818 16398 5844 16454
rect 5900 16398 5926 16454
rect 5982 16398 6008 16454
rect 6064 16398 6090 16454
rect 6146 16398 6172 16454
rect 6228 16398 6254 16454
rect 6310 16398 6336 16454
rect 6392 16398 6418 16454
rect 6474 16398 6500 16454
rect 6556 16398 6582 16454
rect 6638 16398 6664 16454
rect 6720 16398 6746 16454
rect 6802 16398 6828 16454
rect 6884 16398 6909 16454
rect 6965 16398 6990 16454
rect 7046 16398 7071 16454
rect 7127 16398 7152 16454
rect 7208 16398 7233 16454
rect 7289 16398 7314 16454
rect 7370 16398 7379 16454
rect 5179 16374 7379 16398
rect 5179 16318 5188 16374
rect 5244 16318 5270 16374
rect 5326 16318 5352 16374
rect 5408 16318 5434 16374
rect 5490 16318 5516 16374
rect 5572 16318 5598 16374
rect 5654 16318 5680 16374
rect 5736 16318 5762 16374
rect 5818 16318 5844 16374
rect 5900 16318 5926 16374
rect 5982 16318 6008 16374
rect 6064 16318 6090 16374
rect 6146 16318 6172 16374
rect 6228 16318 6254 16374
rect 6310 16318 6336 16374
rect 6392 16318 6418 16374
rect 6474 16318 6500 16374
rect 6556 16318 6582 16374
rect 6638 16318 6664 16374
rect 6720 16318 6746 16374
rect 6802 16318 6828 16374
rect 6884 16318 6909 16374
rect 6965 16318 6990 16374
rect 7046 16318 7071 16374
rect 7127 16318 7152 16374
rect 7208 16318 7233 16374
rect 7289 16318 7314 16374
rect 7370 16318 7379 16374
rect 5179 16294 7379 16318
rect 5179 16238 5188 16294
rect 5244 16238 5270 16294
rect 5326 16238 5352 16294
rect 5408 16238 5434 16294
rect 5490 16238 5516 16294
rect 5572 16238 5598 16294
rect 5654 16238 5680 16294
rect 5736 16238 5762 16294
rect 5818 16238 5844 16294
rect 5900 16238 5926 16294
rect 5982 16238 6008 16294
rect 6064 16238 6090 16294
rect 6146 16238 6172 16294
rect 6228 16238 6254 16294
rect 6310 16238 6336 16294
rect 6392 16238 6418 16294
rect 6474 16238 6500 16294
rect 6556 16238 6582 16294
rect 6638 16238 6664 16294
rect 6720 16238 6746 16294
rect 6802 16238 6828 16294
rect 6884 16238 6909 16294
rect 6965 16238 6990 16294
rect 7046 16238 7071 16294
rect 7127 16238 7152 16294
rect 7208 16238 7233 16294
rect 7289 16238 7314 16294
rect 7370 16238 7379 16294
rect 5179 16214 7379 16238
rect 5179 16158 5188 16214
rect 5244 16158 5270 16214
rect 5326 16158 5352 16214
rect 5408 16158 5434 16214
rect 5490 16158 5516 16214
rect 5572 16158 5598 16214
rect 5654 16158 5680 16214
rect 5736 16158 5762 16214
rect 5818 16158 5844 16214
rect 5900 16158 5926 16214
rect 5982 16158 6008 16214
rect 6064 16158 6090 16214
rect 6146 16158 6172 16214
rect 6228 16158 6254 16214
rect 6310 16158 6336 16214
rect 6392 16158 6418 16214
rect 6474 16158 6500 16214
rect 6556 16158 6582 16214
rect 6638 16158 6664 16214
rect 6720 16158 6746 16214
rect 6802 16158 6828 16214
rect 6884 16158 6909 16214
rect 6965 16158 6990 16214
rect 7046 16158 7071 16214
rect 7127 16158 7152 16214
rect 7208 16158 7233 16214
rect 7289 16158 7314 16214
rect 7370 16158 7379 16214
rect 5179 13294 7379 16158
rect 5179 13238 5188 13294
rect 5244 13238 5270 13294
rect 5326 13238 5352 13294
rect 5408 13238 5434 13294
rect 5490 13238 5516 13294
rect 5572 13238 5598 13294
rect 5654 13238 5680 13294
rect 5736 13238 5762 13294
rect 5818 13238 5844 13294
rect 5900 13238 5926 13294
rect 5982 13238 6008 13294
rect 6064 13238 6090 13294
rect 6146 13238 6172 13294
rect 6228 13238 6254 13294
rect 6310 13238 6336 13294
rect 6392 13238 6418 13294
rect 6474 13238 6500 13294
rect 6556 13238 6582 13294
rect 6638 13238 6664 13294
rect 6720 13238 6746 13294
rect 6802 13238 6828 13294
rect 6884 13238 6909 13294
rect 6965 13238 6990 13294
rect 7046 13238 7071 13294
rect 7127 13238 7152 13294
rect 7208 13238 7233 13294
rect 7289 13238 7314 13294
rect 7370 13238 7379 13294
rect 5179 13214 7379 13238
rect 5179 13158 5188 13214
rect 5244 13158 5270 13214
rect 5326 13158 5352 13214
rect 5408 13158 5434 13214
rect 5490 13158 5516 13214
rect 5572 13158 5598 13214
rect 5654 13158 5680 13214
rect 5736 13158 5762 13214
rect 5818 13158 5844 13214
rect 5900 13158 5926 13214
rect 5982 13158 6008 13214
rect 6064 13158 6090 13214
rect 6146 13158 6172 13214
rect 6228 13158 6254 13214
rect 6310 13158 6336 13214
rect 6392 13158 6418 13214
rect 6474 13158 6500 13214
rect 6556 13158 6582 13214
rect 6638 13158 6664 13214
rect 6720 13158 6746 13214
rect 6802 13158 6828 13214
rect 6884 13158 6909 13214
rect 6965 13158 6990 13214
rect 7046 13158 7071 13214
rect 7127 13158 7152 13214
rect 7208 13158 7233 13214
rect 7289 13158 7314 13214
rect 7370 13158 7379 13214
rect 5179 13134 7379 13158
rect 5179 13078 5188 13134
rect 5244 13078 5270 13134
rect 5326 13078 5352 13134
rect 5408 13078 5434 13134
rect 5490 13078 5516 13134
rect 5572 13078 5598 13134
rect 5654 13078 5680 13134
rect 5736 13078 5762 13134
rect 5818 13078 5844 13134
rect 5900 13078 5926 13134
rect 5982 13078 6008 13134
rect 6064 13078 6090 13134
rect 6146 13078 6172 13134
rect 6228 13078 6254 13134
rect 6310 13078 6336 13134
rect 6392 13078 6418 13134
rect 6474 13078 6500 13134
rect 6556 13078 6582 13134
rect 6638 13078 6664 13134
rect 6720 13078 6746 13134
rect 6802 13078 6828 13134
rect 6884 13078 6909 13134
rect 6965 13078 6990 13134
rect 7046 13078 7071 13134
rect 7127 13078 7152 13134
rect 7208 13078 7233 13134
rect 7289 13078 7314 13134
rect 7370 13078 7379 13134
rect 5179 13054 7379 13078
rect 5179 12998 5188 13054
rect 5244 12998 5270 13054
rect 5326 12998 5352 13054
rect 5408 12998 5434 13054
rect 5490 12998 5516 13054
rect 5572 12998 5598 13054
rect 5654 12998 5680 13054
rect 5736 12998 5762 13054
rect 5818 12998 5844 13054
rect 5900 12998 5926 13054
rect 5982 12998 6008 13054
rect 6064 12998 6090 13054
rect 6146 12998 6172 13054
rect 6228 12998 6254 13054
rect 6310 12998 6336 13054
rect 6392 12998 6418 13054
rect 6474 12998 6500 13054
rect 6556 12998 6582 13054
rect 6638 12998 6664 13054
rect 6720 12998 6746 13054
rect 6802 12998 6828 13054
rect 6884 12998 6909 13054
rect 6965 12998 6990 13054
rect 7046 12998 7071 13054
rect 7127 12998 7152 13054
rect 7208 12998 7233 13054
rect 7289 12998 7314 13054
rect 7370 12998 7379 13054
rect 5179 12974 7379 12998
rect 5179 12918 5188 12974
rect 5244 12918 5270 12974
rect 5326 12918 5352 12974
rect 5408 12918 5434 12974
rect 5490 12918 5516 12974
rect 5572 12918 5598 12974
rect 5654 12918 5680 12974
rect 5736 12918 5762 12974
rect 5818 12918 5844 12974
rect 5900 12918 5926 12974
rect 5982 12918 6008 12974
rect 6064 12918 6090 12974
rect 6146 12918 6172 12974
rect 6228 12918 6254 12974
rect 6310 12918 6336 12974
rect 6392 12918 6418 12974
rect 6474 12918 6500 12974
rect 6556 12918 6582 12974
rect 6638 12918 6664 12974
rect 6720 12918 6746 12974
rect 6802 12918 6828 12974
rect 6884 12918 6909 12974
rect 6965 12918 6990 12974
rect 7046 12918 7071 12974
rect 7127 12918 7152 12974
rect 7208 12918 7233 12974
rect 7289 12918 7314 12974
rect 7370 12918 7379 12974
rect 5179 12894 7379 12918
rect 5179 12838 5188 12894
rect 5244 12838 5270 12894
rect 5326 12838 5352 12894
rect 5408 12838 5434 12894
rect 5490 12838 5516 12894
rect 5572 12838 5598 12894
rect 5654 12838 5680 12894
rect 5736 12838 5762 12894
rect 5818 12838 5844 12894
rect 5900 12838 5926 12894
rect 5982 12838 6008 12894
rect 6064 12838 6090 12894
rect 6146 12838 6172 12894
rect 6228 12838 6254 12894
rect 6310 12838 6336 12894
rect 6392 12838 6418 12894
rect 6474 12838 6500 12894
rect 6556 12838 6582 12894
rect 6638 12838 6664 12894
rect 6720 12838 6746 12894
rect 6802 12838 6828 12894
rect 6884 12838 6909 12894
rect 6965 12838 6990 12894
rect 7046 12838 7071 12894
rect 7127 12838 7152 12894
rect 7208 12838 7233 12894
rect 7289 12838 7314 12894
rect 7370 12838 7379 12894
rect 5179 12814 7379 12838
rect 5179 12758 5188 12814
rect 5244 12758 5270 12814
rect 5326 12758 5352 12814
rect 5408 12758 5434 12814
rect 5490 12758 5516 12814
rect 5572 12758 5598 12814
rect 5654 12758 5680 12814
rect 5736 12758 5762 12814
rect 5818 12758 5844 12814
rect 5900 12758 5926 12814
rect 5982 12758 6008 12814
rect 6064 12758 6090 12814
rect 6146 12758 6172 12814
rect 6228 12758 6254 12814
rect 6310 12758 6336 12814
rect 6392 12758 6418 12814
rect 6474 12758 6500 12814
rect 6556 12758 6582 12814
rect 6638 12758 6664 12814
rect 6720 12758 6746 12814
rect 6802 12758 6828 12814
rect 6884 12758 6909 12814
rect 6965 12758 6990 12814
rect 7046 12758 7071 12814
rect 7127 12758 7152 12814
rect 7208 12758 7233 12814
rect 7289 12758 7314 12814
rect 7370 12758 7379 12814
rect 5179 12734 7379 12758
rect 5179 12678 5188 12734
rect 5244 12678 5270 12734
rect 5326 12678 5352 12734
rect 5408 12678 5434 12734
rect 5490 12678 5516 12734
rect 5572 12678 5598 12734
rect 5654 12678 5680 12734
rect 5736 12678 5762 12734
rect 5818 12678 5844 12734
rect 5900 12678 5926 12734
rect 5982 12678 6008 12734
rect 6064 12678 6090 12734
rect 6146 12678 6172 12734
rect 6228 12678 6254 12734
rect 6310 12678 6336 12734
rect 6392 12678 6418 12734
rect 6474 12678 6500 12734
rect 6556 12678 6582 12734
rect 6638 12678 6664 12734
rect 6720 12678 6746 12734
rect 6802 12678 6828 12734
rect 6884 12678 6909 12734
rect 6965 12678 6990 12734
rect 7046 12678 7071 12734
rect 7127 12678 7152 12734
rect 7208 12678 7233 12734
rect 7289 12678 7314 12734
rect 7370 12678 7379 12734
rect 5179 12654 7379 12678
rect 5179 12598 5188 12654
rect 5244 12598 5270 12654
rect 5326 12598 5352 12654
rect 5408 12598 5434 12654
rect 5490 12598 5516 12654
rect 5572 12598 5598 12654
rect 5654 12598 5680 12654
rect 5736 12598 5762 12654
rect 5818 12598 5844 12654
rect 5900 12598 5926 12654
rect 5982 12598 6008 12654
rect 6064 12598 6090 12654
rect 6146 12598 6172 12654
rect 6228 12598 6254 12654
rect 6310 12598 6336 12654
rect 6392 12598 6418 12654
rect 6474 12598 6500 12654
rect 6556 12598 6582 12654
rect 6638 12598 6664 12654
rect 6720 12598 6746 12654
rect 6802 12598 6828 12654
rect 6884 12598 6909 12654
rect 6965 12598 6990 12654
rect 7046 12598 7071 12654
rect 7127 12598 7152 12654
rect 7208 12598 7233 12654
rect 7289 12598 7314 12654
rect 7370 12598 7379 12654
rect 5179 12574 7379 12598
rect 5179 12518 5188 12574
rect 5244 12518 5270 12574
rect 5326 12518 5352 12574
rect 5408 12518 5434 12574
rect 5490 12518 5516 12574
rect 5572 12518 5598 12574
rect 5654 12518 5680 12574
rect 5736 12518 5762 12574
rect 5818 12518 5844 12574
rect 5900 12518 5926 12574
rect 5982 12518 6008 12574
rect 6064 12518 6090 12574
rect 6146 12518 6172 12574
rect 6228 12518 6254 12574
rect 6310 12518 6336 12574
rect 6392 12518 6418 12574
rect 6474 12518 6500 12574
rect 6556 12518 6582 12574
rect 6638 12518 6664 12574
rect 6720 12518 6746 12574
rect 6802 12518 6828 12574
rect 6884 12518 6909 12574
rect 6965 12518 6990 12574
rect 7046 12518 7071 12574
rect 7127 12518 7152 12574
rect 7208 12518 7233 12574
rect 7289 12518 7314 12574
rect 7370 12518 7379 12574
rect 5179 12494 7379 12518
rect 5179 12438 5188 12494
rect 5244 12438 5270 12494
rect 5326 12438 5352 12494
rect 5408 12438 5434 12494
rect 5490 12438 5516 12494
rect 5572 12438 5598 12494
rect 5654 12438 5680 12494
rect 5736 12438 5762 12494
rect 5818 12438 5844 12494
rect 5900 12438 5926 12494
rect 5982 12438 6008 12494
rect 6064 12438 6090 12494
rect 6146 12438 6172 12494
rect 6228 12438 6254 12494
rect 6310 12438 6336 12494
rect 6392 12438 6418 12494
rect 6474 12438 6500 12494
rect 6556 12438 6582 12494
rect 6638 12438 6664 12494
rect 6720 12438 6746 12494
rect 6802 12438 6828 12494
rect 6884 12438 6909 12494
rect 6965 12438 6990 12494
rect 7046 12438 7071 12494
rect 7127 12438 7152 12494
rect 7208 12438 7233 12494
rect 7289 12438 7314 12494
rect 7370 12438 7379 12494
rect 5179 12414 7379 12438
rect 5179 12358 5188 12414
rect 5244 12358 5270 12414
rect 5326 12358 5352 12414
rect 5408 12358 5434 12414
rect 5490 12358 5516 12414
rect 5572 12358 5598 12414
rect 5654 12358 5680 12414
rect 5736 12358 5762 12414
rect 5818 12358 5844 12414
rect 5900 12358 5926 12414
rect 5982 12358 6008 12414
rect 6064 12358 6090 12414
rect 6146 12358 6172 12414
rect 6228 12358 6254 12414
rect 6310 12358 6336 12414
rect 6392 12358 6418 12414
rect 6474 12358 6500 12414
rect 6556 12358 6582 12414
rect 6638 12358 6664 12414
rect 6720 12358 6746 12414
rect 6802 12358 6828 12414
rect 6884 12358 6909 12414
rect 6965 12358 6990 12414
rect 7046 12358 7071 12414
rect 7127 12358 7152 12414
rect 7208 12358 7233 12414
rect 7289 12358 7314 12414
rect 7370 12358 7379 12414
rect 5179 12334 7379 12358
rect 5179 12278 5188 12334
rect 5244 12278 5270 12334
rect 5326 12278 5352 12334
rect 5408 12278 5434 12334
rect 5490 12278 5516 12334
rect 5572 12278 5598 12334
rect 5654 12278 5680 12334
rect 5736 12278 5762 12334
rect 5818 12278 5844 12334
rect 5900 12278 5926 12334
rect 5982 12278 6008 12334
rect 6064 12278 6090 12334
rect 6146 12278 6172 12334
rect 6228 12278 6254 12334
rect 6310 12278 6336 12334
rect 6392 12278 6418 12334
rect 6474 12278 6500 12334
rect 6556 12278 6582 12334
rect 6638 12278 6664 12334
rect 6720 12278 6746 12334
rect 6802 12278 6828 12334
rect 6884 12278 6909 12334
rect 6965 12278 6990 12334
rect 7046 12278 7071 12334
rect 7127 12278 7152 12334
rect 7208 12278 7233 12334
rect 7289 12278 7314 12334
rect 7370 12278 7379 12334
rect 5179 12254 7379 12278
rect 5179 12198 5188 12254
rect 5244 12198 5270 12254
rect 5326 12198 5352 12254
rect 5408 12198 5434 12254
rect 5490 12198 5516 12254
rect 5572 12198 5598 12254
rect 5654 12198 5680 12254
rect 5736 12198 5762 12254
rect 5818 12198 5844 12254
rect 5900 12198 5926 12254
rect 5982 12198 6008 12254
rect 6064 12198 6090 12254
rect 6146 12198 6172 12254
rect 6228 12198 6254 12254
rect 6310 12198 6336 12254
rect 6392 12198 6418 12254
rect 6474 12198 6500 12254
rect 6556 12198 6582 12254
rect 6638 12198 6664 12254
rect 6720 12198 6746 12254
rect 6802 12198 6828 12254
rect 6884 12198 6909 12254
rect 6965 12198 6990 12254
rect 7046 12198 7071 12254
rect 7127 12198 7152 12254
rect 7208 12198 7233 12254
rect 7289 12198 7314 12254
rect 7370 12198 7379 12254
rect 5179 12174 7379 12198
rect 5179 12118 5188 12174
rect 5244 12118 5270 12174
rect 5326 12118 5352 12174
rect 5408 12118 5434 12174
rect 5490 12118 5516 12174
rect 5572 12118 5598 12174
rect 5654 12118 5680 12174
rect 5736 12118 5762 12174
rect 5818 12118 5844 12174
rect 5900 12118 5926 12174
rect 5982 12118 6008 12174
rect 6064 12118 6090 12174
rect 6146 12118 6172 12174
rect 6228 12118 6254 12174
rect 6310 12118 6336 12174
rect 6392 12118 6418 12174
rect 6474 12118 6500 12174
rect 6556 12118 6582 12174
rect 6638 12118 6664 12174
rect 6720 12118 6746 12174
rect 6802 12118 6828 12174
rect 6884 12118 6909 12174
rect 6965 12118 6990 12174
rect 7046 12118 7071 12174
rect 7127 12118 7152 12174
rect 7208 12118 7233 12174
rect 7289 12118 7314 12174
rect 7370 12118 7379 12174
rect 5179 12094 7379 12118
rect 5179 12038 5188 12094
rect 5244 12038 5270 12094
rect 5326 12038 5352 12094
rect 5408 12038 5434 12094
rect 5490 12038 5516 12094
rect 5572 12038 5598 12094
rect 5654 12038 5680 12094
rect 5736 12038 5762 12094
rect 5818 12038 5844 12094
rect 5900 12038 5926 12094
rect 5982 12038 6008 12094
rect 6064 12038 6090 12094
rect 6146 12038 6172 12094
rect 6228 12038 6254 12094
rect 6310 12038 6336 12094
rect 6392 12038 6418 12094
rect 6474 12038 6500 12094
rect 6556 12038 6582 12094
rect 6638 12038 6664 12094
rect 6720 12038 6746 12094
rect 6802 12038 6828 12094
rect 6884 12038 6909 12094
rect 6965 12038 6990 12094
rect 7046 12038 7071 12094
rect 7127 12038 7152 12094
rect 7208 12038 7233 12094
rect 7289 12038 7314 12094
rect 7370 12038 7379 12094
rect 5179 12014 7379 12038
rect 5179 11958 5188 12014
rect 5244 11958 5270 12014
rect 5326 11958 5352 12014
rect 5408 11958 5434 12014
rect 5490 11958 5516 12014
rect 5572 11958 5598 12014
rect 5654 11958 5680 12014
rect 5736 11958 5762 12014
rect 5818 11958 5844 12014
rect 5900 11958 5926 12014
rect 5982 11958 6008 12014
rect 6064 11958 6090 12014
rect 6146 11958 6172 12014
rect 6228 11958 6254 12014
rect 6310 11958 6336 12014
rect 6392 11958 6418 12014
rect 6474 11958 6500 12014
rect 6556 11958 6582 12014
rect 6638 11958 6664 12014
rect 6720 11958 6746 12014
rect 6802 11958 6828 12014
rect 6884 11958 6909 12014
rect 6965 11958 6990 12014
rect 7046 11958 7071 12014
rect 7127 11958 7152 12014
rect 7208 11958 7233 12014
rect 7289 11958 7314 12014
rect 7370 11958 7379 12014
rect 5179 11934 7379 11958
rect 5179 11878 5188 11934
rect 5244 11878 5270 11934
rect 5326 11878 5352 11934
rect 5408 11878 5434 11934
rect 5490 11878 5516 11934
rect 5572 11878 5598 11934
rect 5654 11878 5680 11934
rect 5736 11878 5762 11934
rect 5818 11878 5844 11934
rect 5900 11878 5926 11934
rect 5982 11878 6008 11934
rect 6064 11878 6090 11934
rect 6146 11878 6172 11934
rect 6228 11878 6254 11934
rect 6310 11878 6336 11934
rect 6392 11878 6418 11934
rect 6474 11878 6500 11934
rect 6556 11878 6582 11934
rect 6638 11878 6664 11934
rect 6720 11878 6746 11934
rect 6802 11878 6828 11934
rect 6884 11878 6909 11934
rect 6965 11878 6990 11934
rect 7046 11878 7071 11934
rect 7127 11878 7152 11934
rect 7208 11878 7233 11934
rect 7289 11878 7314 11934
rect 7370 11878 7379 11934
rect 5179 11854 7379 11878
rect 5179 11798 5188 11854
rect 5244 11798 5270 11854
rect 5326 11798 5352 11854
rect 5408 11798 5434 11854
rect 5490 11798 5516 11854
rect 5572 11798 5598 11854
rect 5654 11798 5680 11854
rect 5736 11798 5762 11854
rect 5818 11798 5844 11854
rect 5900 11798 5926 11854
rect 5982 11798 6008 11854
rect 6064 11798 6090 11854
rect 6146 11798 6172 11854
rect 6228 11798 6254 11854
rect 6310 11798 6336 11854
rect 6392 11798 6418 11854
rect 6474 11798 6500 11854
rect 6556 11798 6582 11854
rect 6638 11798 6664 11854
rect 6720 11798 6746 11854
rect 6802 11798 6828 11854
rect 6884 11798 6909 11854
rect 6965 11798 6990 11854
rect 7046 11798 7071 11854
rect 7127 11798 7152 11854
rect 7208 11798 7233 11854
rect 7289 11798 7314 11854
rect 7370 11798 7379 11854
rect 5179 11774 7379 11798
rect 5179 11718 5188 11774
rect 5244 11718 5270 11774
rect 5326 11718 5352 11774
rect 5408 11718 5434 11774
rect 5490 11718 5516 11774
rect 5572 11718 5598 11774
rect 5654 11718 5680 11774
rect 5736 11718 5762 11774
rect 5818 11718 5844 11774
rect 5900 11718 5926 11774
rect 5982 11718 6008 11774
rect 6064 11718 6090 11774
rect 6146 11718 6172 11774
rect 6228 11718 6254 11774
rect 6310 11718 6336 11774
rect 6392 11718 6418 11774
rect 6474 11718 6500 11774
rect 6556 11718 6582 11774
rect 6638 11718 6664 11774
rect 6720 11718 6746 11774
rect 6802 11718 6828 11774
rect 6884 11718 6909 11774
rect 6965 11718 6990 11774
rect 7046 11718 7071 11774
rect 7127 11718 7152 11774
rect 7208 11718 7233 11774
rect 7289 11718 7314 11774
rect 7370 11718 7379 11774
rect 5179 11694 7379 11718
rect 5179 11638 5188 11694
rect 5244 11638 5270 11694
rect 5326 11638 5352 11694
rect 5408 11638 5434 11694
rect 5490 11638 5516 11694
rect 5572 11638 5598 11694
rect 5654 11638 5680 11694
rect 5736 11638 5762 11694
rect 5818 11638 5844 11694
rect 5900 11638 5926 11694
rect 5982 11638 6008 11694
rect 6064 11638 6090 11694
rect 6146 11638 6172 11694
rect 6228 11638 6254 11694
rect 6310 11638 6336 11694
rect 6392 11638 6418 11694
rect 6474 11638 6500 11694
rect 6556 11638 6582 11694
rect 6638 11638 6664 11694
rect 6720 11638 6746 11694
rect 6802 11638 6828 11694
rect 6884 11638 6909 11694
rect 6965 11638 6990 11694
rect 7046 11638 7071 11694
rect 7127 11638 7152 11694
rect 7208 11638 7233 11694
rect 7289 11638 7314 11694
rect 7370 11638 7379 11694
rect 5179 11614 7379 11638
rect 5179 11558 5188 11614
rect 5244 11558 5270 11614
rect 5326 11558 5352 11614
rect 5408 11558 5434 11614
rect 5490 11558 5516 11614
rect 5572 11558 5598 11614
rect 5654 11558 5680 11614
rect 5736 11558 5762 11614
rect 5818 11558 5844 11614
rect 5900 11558 5926 11614
rect 5982 11558 6008 11614
rect 6064 11558 6090 11614
rect 6146 11558 6172 11614
rect 6228 11558 6254 11614
rect 6310 11558 6336 11614
rect 6392 11558 6418 11614
rect 6474 11558 6500 11614
rect 6556 11558 6582 11614
rect 6638 11558 6664 11614
rect 6720 11558 6746 11614
rect 6802 11558 6828 11614
rect 6884 11558 6909 11614
rect 6965 11558 6990 11614
rect 7046 11558 7071 11614
rect 7127 11558 7152 11614
rect 7208 11558 7233 11614
rect 7289 11558 7314 11614
rect 7370 11558 7379 11614
rect 5179 5101 7379 11558
rect 5179 5045 5191 5101
rect 5247 5045 5273 5101
rect 5329 5045 5355 5101
rect 5411 5045 5437 5101
rect 5493 5045 5519 5101
rect 5575 5045 5601 5101
rect 5657 5045 5683 5101
rect 5739 5045 5765 5101
rect 5821 5045 5847 5101
rect 5903 5045 5929 5101
rect 5985 5045 6011 5101
rect 6067 5045 6093 5101
rect 6149 5045 6175 5101
rect 6231 5045 6257 5101
rect 6313 5045 6339 5101
rect 6395 5045 6421 5101
rect 6477 5045 6503 5101
rect 6559 5045 6585 5101
rect 6641 5045 6666 5101
rect 6722 5045 6747 5101
rect 6803 5045 6828 5101
rect 6884 5045 6909 5101
rect 6965 5045 6990 5101
rect 7046 5045 7071 5101
rect 7127 5045 7152 5101
rect 7208 5045 7233 5101
rect 7289 5045 7314 5101
rect 7370 5045 7379 5101
rect 5179 5021 7379 5045
rect 5179 4965 5191 5021
rect 5247 4965 5273 5021
rect 5329 4965 5355 5021
rect 5411 4965 5437 5021
rect 5493 4965 5519 5021
rect 5575 4965 5601 5021
rect 5657 4965 5683 5021
rect 5739 4965 5765 5021
rect 5821 4965 5847 5021
rect 5903 4965 5929 5021
rect 5985 4965 6011 5021
rect 6067 4965 6093 5021
rect 6149 4965 6175 5021
rect 6231 4965 6257 5021
rect 6313 4965 6339 5021
rect 6395 4965 6421 5021
rect 6477 4965 6503 5021
rect 6559 4965 6585 5021
rect 6641 4965 6666 5021
rect 6722 4965 6747 5021
rect 6803 4965 6828 5021
rect 6884 4965 6909 5021
rect 6965 4965 6990 5021
rect 7046 4965 7071 5021
rect 7127 4965 7152 5021
rect 7208 4965 7233 5021
rect 7289 4965 7314 5021
rect 7370 4965 7379 5021
rect 5179 4941 7379 4965
rect 5179 4885 5191 4941
rect 5247 4885 5273 4941
rect 5329 4885 5355 4941
rect 5411 4885 5437 4941
rect 5493 4885 5519 4941
rect 5575 4885 5601 4941
rect 5657 4885 5683 4941
rect 5739 4885 5765 4941
rect 5821 4885 5847 4941
rect 5903 4885 5929 4941
rect 5985 4885 6011 4941
rect 6067 4885 6093 4941
rect 6149 4885 6175 4941
rect 6231 4885 6257 4941
rect 6313 4885 6339 4941
rect 6395 4885 6421 4941
rect 6477 4885 6503 4941
rect 6559 4885 6585 4941
rect 6641 4885 6666 4941
rect 6722 4885 6747 4941
rect 6803 4885 6828 4941
rect 6884 4885 6909 4941
rect 6965 4885 6990 4941
rect 7046 4885 7071 4941
rect 7127 4885 7152 4941
rect 7208 4885 7233 4941
rect 7289 4885 7314 4941
rect 7370 4885 7379 4941
rect 5179 4861 7379 4885
rect 5179 4805 5191 4861
rect 5247 4805 5273 4861
rect 5329 4805 5355 4861
rect 5411 4805 5437 4861
rect 5493 4805 5519 4861
rect 5575 4805 5601 4861
rect 5657 4805 5683 4861
rect 5739 4805 5765 4861
rect 5821 4805 5847 4861
rect 5903 4805 5929 4861
rect 5985 4805 6011 4861
rect 6067 4805 6093 4861
rect 6149 4805 6175 4861
rect 6231 4805 6257 4861
rect 6313 4805 6339 4861
rect 6395 4805 6421 4861
rect 6477 4805 6503 4861
rect 6559 4805 6585 4861
rect 6641 4805 6666 4861
rect 6722 4805 6747 4861
rect 6803 4805 6828 4861
rect 6884 4805 6909 4861
rect 6965 4805 6990 4861
rect 7046 4805 7071 4861
rect 7127 4805 7152 4861
rect 7208 4805 7233 4861
rect 7289 4805 7314 4861
rect 7370 4805 7379 4861
rect 5179 4781 7379 4805
rect 5179 4725 5191 4781
rect 5247 4725 5273 4781
rect 5329 4725 5355 4781
rect 5411 4725 5437 4781
rect 5493 4725 5519 4781
rect 5575 4725 5601 4781
rect 5657 4725 5683 4781
rect 5739 4725 5765 4781
rect 5821 4725 5847 4781
rect 5903 4725 5929 4781
rect 5985 4725 6011 4781
rect 6067 4725 6093 4781
rect 6149 4725 6175 4781
rect 6231 4725 6257 4781
rect 6313 4725 6339 4781
rect 6395 4725 6421 4781
rect 6477 4725 6503 4781
rect 6559 4725 6585 4781
rect 6641 4725 6666 4781
rect 6722 4725 6747 4781
rect 6803 4725 6828 4781
rect 6884 4725 6909 4781
rect 6965 4725 6990 4781
rect 7046 4725 7071 4781
rect 7127 4725 7152 4781
rect 7208 4725 7233 4781
rect 7289 4725 7314 4781
rect 7370 4725 7379 4781
rect 5179 4701 7379 4725
rect 5179 4645 5191 4701
rect 5247 4645 5273 4701
rect 5329 4645 5355 4701
rect 5411 4645 5437 4701
rect 5493 4645 5519 4701
rect 5575 4645 5601 4701
rect 5657 4645 5683 4701
rect 5739 4645 5765 4701
rect 5821 4645 5847 4701
rect 5903 4645 5929 4701
rect 5985 4645 6011 4701
rect 6067 4645 6093 4701
rect 6149 4645 6175 4701
rect 6231 4645 6257 4701
rect 6313 4645 6339 4701
rect 6395 4645 6421 4701
rect 6477 4645 6503 4701
rect 6559 4645 6585 4701
rect 6641 4645 6666 4701
rect 6722 4645 6747 4701
rect 6803 4645 6828 4701
rect 6884 4645 6909 4701
rect 6965 4645 6990 4701
rect 7046 4645 7071 4701
rect 7127 4645 7152 4701
rect 7208 4645 7233 4701
rect 7289 4645 7314 4701
rect 7370 4645 7379 4701
rect 5179 4621 7379 4645
rect 5179 4565 5191 4621
rect 5247 4565 5273 4621
rect 5329 4565 5355 4621
rect 5411 4565 5437 4621
rect 5493 4565 5519 4621
rect 5575 4565 5601 4621
rect 5657 4565 5683 4621
rect 5739 4565 5765 4621
rect 5821 4565 5847 4621
rect 5903 4565 5929 4621
rect 5985 4565 6011 4621
rect 6067 4565 6093 4621
rect 6149 4565 6175 4621
rect 6231 4565 6257 4621
rect 6313 4565 6339 4621
rect 6395 4565 6421 4621
rect 6477 4565 6503 4621
rect 6559 4565 6585 4621
rect 6641 4565 6666 4621
rect 6722 4565 6747 4621
rect 6803 4565 6828 4621
rect 6884 4565 6909 4621
rect 6965 4565 6990 4621
rect 7046 4565 7071 4621
rect 7127 4565 7152 4621
rect 7208 4565 7233 4621
rect 7289 4565 7314 4621
rect 7370 4565 7379 4621
rect 5179 4541 7379 4565
rect 5179 4485 5191 4541
rect 5247 4485 5273 4541
rect 5329 4485 5355 4541
rect 5411 4485 5437 4541
rect 5493 4485 5519 4541
rect 5575 4485 5601 4541
rect 5657 4485 5683 4541
rect 5739 4485 5765 4541
rect 5821 4485 5847 4541
rect 5903 4485 5929 4541
rect 5985 4485 6011 4541
rect 6067 4485 6093 4541
rect 6149 4485 6175 4541
rect 6231 4485 6257 4541
rect 6313 4485 6339 4541
rect 6395 4485 6421 4541
rect 6477 4485 6503 4541
rect 6559 4485 6585 4541
rect 6641 4485 6666 4541
rect 6722 4485 6747 4541
rect 6803 4485 6828 4541
rect 6884 4485 6909 4541
rect 6965 4485 6990 4541
rect 7046 4485 7071 4541
rect 7127 4485 7152 4541
rect 7208 4485 7233 4541
rect 7289 4485 7314 4541
rect 7370 4485 7379 4541
rect 5179 4461 7379 4485
rect 5179 4405 5191 4461
rect 5247 4405 5273 4461
rect 5329 4405 5355 4461
rect 5411 4405 5437 4461
rect 5493 4405 5519 4461
rect 5575 4405 5601 4461
rect 5657 4405 5683 4461
rect 5739 4405 5765 4461
rect 5821 4405 5847 4461
rect 5903 4405 5929 4461
rect 5985 4405 6011 4461
rect 6067 4405 6093 4461
rect 6149 4405 6175 4461
rect 6231 4405 6257 4461
rect 6313 4405 6339 4461
rect 6395 4405 6421 4461
rect 6477 4405 6503 4461
rect 6559 4405 6585 4461
rect 6641 4405 6666 4461
rect 6722 4405 6747 4461
rect 6803 4405 6828 4461
rect 6884 4405 6909 4461
rect 6965 4405 6990 4461
rect 7046 4405 7071 4461
rect 7127 4405 7152 4461
rect 7208 4405 7233 4461
rect 7289 4405 7314 4461
rect 7370 4405 7379 4461
rect 5179 4381 7379 4405
rect 5179 4325 5191 4381
rect 5247 4325 5273 4381
rect 5329 4325 5355 4381
rect 5411 4325 5437 4381
rect 5493 4325 5519 4381
rect 5575 4325 5601 4381
rect 5657 4325 5683 4381
rect 5739 4325 5765 4381
rect 5821 4325 5847 4381
rect 5903 4325 5929 4381
rect 5985 4325 6011 4381
rect 6067 4325 6093 4381
rect 6149 4325 6175 4381
rect 6231 4325 6257 4381
rect 6313 4325 6339 4381
rect 6395 4325 6421 4381
rect 6477 4325 6503 4381
rect 6559 4325 6585 4381
rect 6641 4325 6666 4381
rect 6722 4325 6747 4381
rect 6803 4325 6828 4381
rect 6884 4325 6909 4381
rect 6965 4325 6990 4381
rect 7046 4325 7071 4381
rect 7127 4325 7152 4381
rect 7208 4325 7233 4381
rect 7289 4325 7314 4381
rect 7370 4325 7379 4381
rect 5179 4301 7379 4325
rect 5179 4245 5191 4301
rect 5247 4245 5273 4301
rect 5329 4245 5355 4301
rect 5411 4245 5437 4301
rect 5493 4245 5519 4301
rect 5575 4245 5601 4301
rect 5657 4245 5683 4301
rect 5739 4245 5765 4301
rect 5821 4245 5847 4301
rect 5903 4245 5929 4301
rect 5985 4245 6011 4301
rect 6067 4245 6093 4301
rect 6149 4245 6175 4301
rect 6231 4245 6257 4301
rect 6313 4245 6339 4301
rect 6395 4245 6421 4301
rect 6477 4245 6503 4301
rect 6559 4245 6585 4301
rect 6641 4245 6666 4301
rect 6722 4245 6747 4301
rect 6803 4245 6828 4301
rect 6884 4245 6909 4301
rect 6965 4245 6990 4301
rect 7046 4245 7071 4301
rect 7127 4245 7152 4301
rect 7208 4245 7233 4301
rect 7289 4245 7314 4301
rect 7370 4245 7379 4301
rect 5179 4221 7379 4245
rect 5179 4165 5191 4221
rect 5247 4165 5273 4221
rect 5329 4165 5355 4221
rect 5411 4165 5437 4221
rect 5493 4165 5519 4221
rect 5575 4165 5601 4221
rect 5657 4165 5683 4221
rect 5739 4165 5765 4221
rect 5821 4165 5847 4221
rect 5903 4165 5929 4221
rect 5985 4165 6011 4221
rect 6067 4165 6093 4221
rect 6149 4165 6175 4221
rect 6231 4165 6257 4221
rect 6313 4165 6339 4221
rect 6395 4165 6421 4221
rect 6477 4165 6503 4221
rect 6559 4165 6585 4221
rect 6641 4165 6666 4221
rect 6722 4165 6747 4221
rect 6803 4165 6828 4221
rect 6884 4165 6909 4221
rect 6965 4165 6990 4221
rect 7046 4165 7071 4221
rect 7127 4165 7152 4221
rect 7208 4165 7233 4221
rect 7289 4165 7314 4221
rect 7370 4165 7379 4221
rect 5179 4141 7379 4165
rect 5179 4085 5191 4141
rect 5247 4085 5273 4141
rect 5329 4085 5355 4141
rect 5411 4085 5437 4141
rect 5493 4085 5519 4141
rect 5575 4085 5601 4141
rect 5657 4085 5683 4141
rect 5739 4085 5765 4141
rect 5821 4085 5847 4141
rect 5903 4085 5929 4141
rect 5985 4085 6011 4141
rect 6067 4085 6093 4141
rect 6149 4085 6175 4141
rect 6231 4085 6257 4141
rect 6313 4085 6339 4141
rect 6395 4085 6421 4141
rect 6477 4085 6503 4141
rect 6559 4085 6585 4141
rect 6641 4085 6666 4141
rect 6722 4085 6747 4141
rect 6803 4085 6828 4141
rect 6884 4085 6909 4141
rect 6965 4085 6990 4141
rect 7046 4085 7071 4141
rect 7127 4085 7152 4141
rect 7208 4085 7233 4141
rect 7289 4085 7314 4141
rect 7370 4085 7379 4141
rect 5179 4061 7379 4085
rect 5179 4005 5191 4061
rect 5247 4005 5273 4061
rect 5329 4005 5355 4061
rect 5411 4005 5437 4061
rect 5493 4005 5519 4061
rect 5575 4005 5601 4061
rect 5657 4005 5683 4061
rect 5739 4005 5765 4061
rect 5821 4005 5847 4061
rect 5903 4005 5929 4061
rect 5985 4005 6011 4061
rect 6067 4005 6093 4061
rect 6149 4005 6175 4061
rect 6231 4005 6257 4061
rect 6313 4005 6339 4061
rect 6395 4005 6421 4061
rect 6477 4005 6503 4061
rect 6559 4005 6585 4061
rect 6641 4005 6666 4061
rect 6722 4005 6747 4061
rect 6803 4005 6828 4061
rect 6884 4005 6909 4061
rect 6965 4005 6990 4061
rect 7046 4005 7071 4061
rect 7127 4005 7152 4061
rect 7208 4005 7233 4061
rect 7289 4005 7314 4061
rect 7370 4005 7379 4061
rect 5179 3981 7379 4005
rect 5179 3925 5191 3981
rect 5247 3925 5273 3981
rect 5329 3925 5355 3981
rect 5411 3925 5437 3981
rect 5493 3925 5519 3981
rect 5575 3925 5601 3981
rect 5657 3925 5683 3981
rect 5739 3925 5765 3981
rect 5821 3925 5847 3981
rect 5903 3925 5929 3981
rect 5985 3925 6011 3981
rect 6067 3925 6093 3981
rect 6149 3925 6175 3981
rect 6231 3925 6257 3981
rect 6313 3925 6339 3981
rect 6395 3925 6421 3981
rect 6477 3925 6503 3981
rect 6559 3925 6585 3981
rect 6641 3925 6666 3981
rect 6722 3925 6747 3981
rect 6803 3925 6828 3981
rect 6884 3925 6909 3981
rect 6965 3925 6990 3981
rect 7046 3925 7071 3981
rect 7127 3925 7152 3981
rect 7208 3925 7233 3981
rect 7289 3925 7314 3981
rect 7370 3925 7379 3981
rect 5179 3901 7379 3925
rect 5179 3845 5191 3901
rect 5247 3845 5273 3901
rect 5329 3845 5355 3901
rect 5411 3845 5437 3901
rect 5493 3845 5519 3901
rect 5575 3845 5601 3901
rect 5657 3845 5683 3901
rect 5739 3845 5765 3901
rect 5821 3845 5847 3901
rect 5903 3845 5929 3901
rect 5985 3845 6011 3901
rect 6067 3845 6093 3901
rect 6149 3845 6175 3901
rect 6231 3845 6257 3901
rect 6313 3845 6339 3901
rect 6395 3845 6421 3901
rect 6477 3845 6503 3901
rect 6559 3845 6585 3901
rect 6641 3845 6666 3901
rect 6722 3845 6747 3901
rect 6803 3845 6828 3901
rect 6884 3845 6909 3901
rect 6965 3845 6990 3901
rect 7046 3845 7071 3901
rect 7127 3845 7152 3901
rect 7208 3845 7233 3901
rect 7289 3845 7314 3901
rect 7370 3845 7379 3901
rect 5179 3821 7379 3845
rect 5179 3765 5191 3821
rect 5247 3765 5273 3821
rect 5329 3765 5355 3821
rect 5411 3765 5437 3821
rect 5493 3765 5519 3821
rect 5575 3765 5601 3821
rect 5657 3765 5683 3821
rect 5739 3765 5765 3821
rect 5821 3765 5847 3821
rect 5903 3765 5929 3821
rect 5985 3765 6011 3821
rect 6067 3765 6093 3821
rect 6149 3765 6175 3821
rect 6231 3765 6257 3821
rect 6313 3765 6339 3821
rect 6395 3765 6421 3821
rect 6477 3765 6503 3821
rect 6559 3765 6585 3821
rect 6641 3765 6666 3821
rect 6722 3765 6747 3821
rect 6803 3765 6828 3821
rect 6884 3765 6909 3821
rect 6965 3765 6990 3821
rect 7046 3765 7071 3821
rect 7127 3765 7152 3821
rect 7208 3765 7233 3821
rect 7289 3765 7314 3821
rect 7370 3765 7379 3821
rect 5179 3741 7379 3765
rect 5179 3685 5191 3741
rect 5247 3685 5273 3741
rect 5329 3685 5355 3741
rect 5411 3685 5437 3741
rect 5493 3685 5519 3741
rect 5575 3685 5601 3741
rect 5657 3685 5683 3741
rect 5739 3685 5765 3741
rect 5821 3685 5847 3741
rect 5903 3685 5929 3741
rect 5985 3685 6011 3741
rect 6067 3685 6093 3741
rect 6149 3685 6175 3741
rect 6231 3685 6257 3741
rect 6313 3685 6339 3741
rect 6395 3685 6421 3741
rect 6477 3685 6503 3741
rect 6559 3685 6585 3741
rect 6641 3685 6666 3741
rect 6722 3685 6747 3741
rect 6803 3685 6828 3741
rect 6884 3685 6909 3741
rect 6965 3685 6990 3741
rect 7046 3685 7071 3741
rect 7127 3685 7152 3741
rect 7208 3685 7233 3741
rect 7289 3685 7314 3741
rect 7370 3685 7379 3741
rect 5179 3661 7379 3685
rect 5179 3605 5191 3661
rect 5247 3605 5273 3661
rect 5329 3605 5355 3661
rect 5411 3605 5437 3661
rect 5493 3605 5519 3661
rect 5575 3605 5601 3661
rect 5657 3605 5683 3661
rect 5739 3605 5765 3661
rect 5821 3605 5847 3661
rect 5903 3605 5929 3661
rect 5985 3605 6011 3661
rect 6067 3605 6093 3661
rect 6149 3605 6175 3661
rect 6231 3605 6257 3661
rect 6313 3605 6339 3661
rect 6395 3605 6421 3661
rect 6477 3605 6503 3661
rect 6559 3605 6585 3661
rect 6641 3605 6666 3661
rect 6722 3605 6747 3661
rect 6803 3605 6828 3661
rect 6884 3605 6909 3661
rect 6965 3605 6990 3661
rect 7046 3605 7071 3661
rect 7127 3605 7152 3661
rect 7208 3605 7233 3661
rect 7289 3605 7314 3661
rect 7370 3605 7379 3661
rect 5179 3581 7379 3605
rect 5179 3525 5191 3581
rect 5247 3525 5273 3581
rect 5329 3525 5355 3581
rect 5411 3525 5437 3581
rect 5493 3525 5519 3581
rect 5575 3525 5601 3581
rect 5657 3525 5683 3581
rect 5739 3525 5765 3581
rect 5821 3525 5847 3581
rect 5903 3525 5929 3581
rect 5985 3525 6011 3581
rect 6067 3525 6093 3581
rect 6149 3525 6175 3581
rect 6231 3525 6257 3581
rect 6313 3525 6339 3581
rect 6395 3525 6421 3581
rect 6477 3525 6503 3581
rect 6559 3525 6585 3581
rect 6641 3525 6666 3581
rect 6722 3525 6747 3581
rect 6803 3525 6828 3581
rect 6884 3525 6909 3581
rect 6965 3525 6990 3581
rect 7046 3525 7071 3581
rect 7127 3525 7152 3581
rect 7208 3525 7233 3581
rect 7289 3525 7314 3581
rect 7370 3525 7379 3581
rect 5179 3501 7379 3525
rect 5179 3445 5191 3501
rect 5247 3445 5273 3501
rect 5329 3445 5355 3501
rect 5411 3445 5437 3501
rect 5493 3445 5519 3501
rect 5575 3445 5601 3501
rect 5657 3445 5683 3501
rect 5739 3445 5765 3501
rect 5821 3445 5847 3501
rect 5903 3445 5929 3501
rect 5985 3445 6011 3501
rect 6067 3445 6093 3501
rect 6149 3445 6175 3501
rect 6231 3445 6257 3501
rect 6313 3445 6339 3501
rect 6395 3445 6421 3501
rect 6477 3445 6503 3501
rect 6559 3445 6585 3501
rect 6641 3445 6666 3501
rect 6722 3445 6747 3501
rect 6803 3445 6828 3501
rect 6884 3445 6909 3501
rect 6965 3445 6990 3501
rect 7046 3445 7071 3501
rect 7127 3445 7152 3501
rect 7208 3445 7233 3501
rect 7289 3445 7314 3501
rect 7370 3445 7379 3501
rect 5179 3421 7379 3445
rect 5179 3365 5191 3421
rect 5247 3365 5273 3421
rect 5329 3365 5355 3421
rect 5411 3365 5437 3421
rect 5493 3365 5519 3421
rect 5575 3365 5601 3421
rect 5657 3365 5683 3421
rect 5739 3365 5765 3421
rect 5821 3365 5847 3421
rect 5903 3365 5929 3421
rect 5985 3365 6011 3421
rect 6067 3365 6093 3421
rect 6149 3365 6175 3421
rect 6231 3365 6257 3421
rect 6313 3365 6339 3421
rect 6395 3365 6421 3421
rect 6477 3365 6503 3421
rect 6559 3365 6585 3421
rect 6641 3365 6666 3421
rect 6722 3365 6747 3421
rect 6803 3365 6828 3421
rect 6884 3365 6909 3421
rect 6965 3365 6990 3421
rect 7046 3365 7071 3421
rect 7127 3365 7152 3421
rect 7208 3365 7233 3421
rect 7289 3365 7314 3421
rect 7370 3365 7379 3421
rect 5179 3341 7379 3365
rect 5179 3285 5191 3341
rect 5247 3285 5273 3341
rect 5329 3285 5355 3341
rect 5411 3285 5437 3341
rect 5493 3285 5519 3341
rect 5575 3285 5601 3341
rect 5657 3285 5683 3341
rect 5739 3285 5765 3341
rect 5821 3285 5847 3341
rect 5903 3285 5929 3341
rect 5985 3285 6011 3341
rect 6067 3285 6093 3341
rect 6149 3285 6175 3341
rect 6231 3285 6257 3341
rect 6313 3285 6339 3341
rect 6395 3285 6421 3341
rect 6477 3285 6503 3341
rect 6559 3285 6585 3341
rect 6641 3285 6666 3341
rect 6722 3285 6747 3341
rect 6803 3285 6828 3341
rect 6884 3285 6909 3341
rect 6965 3285 6990 3341
rect 7046 3285 7071 3341
rect 7127 3285 7152 3341
rect 7208 3285 7233 3341
rect 7289 3285 7314 3341
rect 7370 3285 7379 3341
rect 5179 3261 7379 3285
rect 5179 3205 5191 3261
rect 5247 3205 5273 3261
rect 5329 3205 5355 3261
rect 5411 3205 5437 3261
rect 5493 3205 5519 3261
rect 5575 3205 5601 3261
rect 5657 3205 5683 3261
rect 5739 3205 5765 3261
rect 5821 3205 5847 3261
rect 5903 3205 5929 3261
rect 5985 3205 6011 3261
rect 6067 3205 6093 3261
rect 6149 3205 6175 3261
rect 6231 3205 6257 3261
rect 6313 3205 6339 3261
rect 6395 3205 6421 3261
rect 6477 3205 6503 3261
rect 6559 3205 6585 3261
rect 6641 3205 6666 3261
rect 6722 3205 6747 3261
rect 6803 3205 6828 3261
rect 6884 3205 6909 3261
rect 6965 3205 6990 3261
rect 7046 3205 7071 3261
rect 7127 3205 7152 3261
rect 7208 3205 7233 3261
rect 7289 3205 7314 3261
rect 7370 3205 7379 3261
rect 5179 3181 7379 3205
rect 5179 3125 5191 3181
rect 5247 3125 5273 3181
rect 5329 3125 5355 3181
rect 5411 3125 5437 3181
rect 5493 3125 5519 3181
rect 5575 3125 5601 3181
rect 5657 3125 5683 3181
rect 5739 3125 5765 3181
rect 5821 3125 5847 3181
rect 5903 3125 5929 3181
rect 5985 3125 6011 3181
rect 6067 3125 6093 3181
rect 6149 3125 6175 3181
rect 6231 3125 6257 3181
rect 6313 3125 6339 3181
rect 6395 3125 6421 3181
rect 6477 3125 6503 3181
rect 6559 3125 6585 3181
rect 6641 3125 6666 3181
rect 6722 3125 6747 3181
rect 6803 3125 6828 3181
rect 6884 3125 6909 3181
rect 6965 3125 6990 3181
rect 7046 3125 7071 3181
rect 7127 3125 7152 3181
rect 7208 3125 7233 3181
rect 7289 3125 7314 3181
rect 7370 3125 7379 3181
rect 5179 3101 7379 3125
rect 5179 3045 5191 3101
rect 5247 3045 5273 3101
rect 5329 3045 5355 3101
rect 5411 3045 5437 3101
rect 5493 3045 5519 3101
rect 5575 3045 5601 3101
rect 5657 3045 5683 3101
rect 5739 3045 5765 3101
rect 5821 3045 5847 3101
rect 5903 3045 5929 3101
rect 5985 3045 6011 3101
rect 6067 3045 6093 3101
rect 6149 3045 6175 3101
rect 6231 3045 6257 3101
rect 6313 3045 6339 3101
rect 6395 3045 6421 3101
rect 6477 3045 6503 3101
rect 6559 3045 6585 3101
rect 6641 3045 6666 3101
rect 6722 3045 6747 3101
rect 6803 3045 6828 3101
rect 6884 3045 6909 3101
rect 6965 3045 6990 3101
rect 7046 3045 7071 3101
rect 7127 3045 7152 3101
rect 7208 3045 7233 3101
rect 7289 3045 7314 3101
rect 7370 3045 7379 3101
rect 5179 3021 7379 3045
rect 5179 2965 5191 3021
rect 5247 2965 5273 3021
rect 5329 2965 5355 3021
rect 5411 2965 5437 3021
rect 5493 2965 5519 3021
rect 5575 2965 5601 3021
rect 5657 2965 5683 3021
rect 5739 2965 5765 3021
rect 5821 2965 5847 3021
rect 5903 2965 5929 3021
rect 5985 2965 6011 3021
rect 6067 2965 6093 3021
rect 6149 2965 6175 3021
rect 6231 2965 6257 3021
rect 6313 2965 6339 3021
rect 6395 2965 6421 3021
rect 6477 2965 6503 3021
rect 6559 2965 6585 3021
rect 6641 2965 6666 3021
rect 6722 2965 6747 3021
rect 6803 2965 6828 3021
rect 6884 2965 6909 3021
rect 6965 2965 6990 3021
rect 7046 2965 7071 3021
rect 7127 2965 7152 3021
rect 7208 2965 7233 3021
rect 7289 2965 7314 3021
rect 7370 2965 7379 3021
rect 5179 2941 7379 2965
rect 5179 2885 5191 2941
rect 5247 2885 5273 2941
rect 5329 2885 5355 2941
rect 5411 2885 5437 2941
rect 5493 2885 5519 2941
rect 5575 2885 5601 2941
rect 5657 2885 5683 2941
rect 5739 2885 5765 2941
rect 5821 2885 5847 2941
rect 5903 2885 5929 2941
rect 5985 2885 6011 2941
rect 6067 2885 6093 2941
rect 6149 2885 6175 2941
rect 6231 2885 6257 2941
rect 6313 2885 6339 2941
rect 6395 2885 6421 2941
rect 6477 2885 6503 2941
rect 6559 2885 6585 2941
rect 6641 2885 6666 2941
rect 6722 2885 6747 2941
rect 6803 2885 6828 2941
rect 6884 2885 6909 2941
rect 6965 2885 6990 2941
rect 7046 2885 7071 2941
rect 7127 2885 7152 2941
rect 7208 2885 7233 2941
rect 7289 2885 7314 2941
rect 7370 2885 7379 2941
rect 5179 2861 7379 2885
rect 5179 2805 5191 2861
rect 5247 2805 5273 2861
rect 5329 2805 5355 2861
rect 5411 2805 5437 2861
rect 5493 2805 5519 2861
rect 5575 2805 5601 2861
rect 5657 2805 5683 2861
rect 5739 2805 5765 2861
rect 5821 2805 5847 2861
rect 5903 2805 5929 2861
rect 5985 2805 6011 2861
rect 6067 2805 6093 2861
rect 6149 2805 6175 2861
rect 6231 2805 6257 2861
rect 6313 2805 6339 2861
rect 6395 2805 6421 2861
rect 6477 2805 6503 2861
rect 6559 2805 6585 2861
rect 6641 2805 6666 2861
rect 6722 2805 6747 2861
rect 6803 2805 6828 2861
rect 6884 2805 6909 2861
rect 6965 2805 6990 2861
rect 7046 2805 7071 2861
rect 7127 2805 7152 2861
rect 7208 2805 7233 2861
rect 7289 2805 7314 2861
rect 7370 2805 7379 2861
rect 5179 2781 7379 2805
rect 5179 2725 5191 2781
rect 5247 2725 5273 2781
rect 5329 2725 5355 2781
rect 5411 2725 5437 2781
rect 5493 2725 5519 2781
rect 5575 2725 5601 2781
rect 5657 2725 5683 2781
rect 5739 2725 5765 2781
rect 5821 2725 5847 2781
rect 5903 2725 5929 2781
rect 5985 2725 6011 2781
rect 6067 2725 6093 2781
rect 6149 2725 6175 2781
rect 6231 2725 6257 2781
rect 6313 2725 6339 2781
rect 6395 2725 6421 2781
rect 6477 2725 6503 2781
rect 6559 2725 6585 2781
rect 6641 2725 6666 2781
rect 6722 2725 6747 2781
rect 6803 2725 6828 2781
rect 6884 2725 6909 2781
rect 6965 2725 6990 2781
rect 7046 2725 7071 2781
rect 7127 2725 7152 2781
rect 7208 2725 7233 2781
rect 7289 2725 7314 2781
rect 7370 2725 7379 2781
rect 5179 2701 7379 2725
rect 5179 2645 5191 2701
rect 5247 2645 5273 2701
rect 5329 2645 5355 2701
rect 5411 2645 5437 2701
rect 5493 2645 5519 2701
rect 5575 2645 5601 2701
rect 5657 2645 5683 2701
rect 5739 2645 5765 2701
rect 5821 2645 5847 2701
rect 5903 2645 5929 2701
rect 5985 2645 6011 2701
rect 6067 2645 6093 2701
rect 6149 2645 6175 2701
rect 6231 2645 6257 2701
rect 6313 2645 6339 2701
rect 6395 2645 6421 2701
rect 6477 2645 6503 2701
rect 6559 2645 6585 2701
rect 6641 2645 6666 2701
rect 6722 2645 6747 2701
rect 6803 2645 6828 2701
rect 6884 2645 6909 2701
rect 6965 2645 6990 2701
rect 7046 2645 7071 2701
rect 7127 2645 7152 2701
rect 7208 2645 7233 2701
rect 7289 2645 7314 2701
rect 7370 2645 7379 2701
rect 5179 2621 7379 2645
rect 5179 2565 5191 2621
rect 5247 2565 5273 2621
rect 5329 2565 5355 2621
rect 5411 2565 5437 2621
rect 5493 2565 5519 2621
rect 5575 2565 5601 2621
rect 5657 2565 5683 2621
rect 5739 2565 5765 2621
rect 5821 2565 5847 2621
rect 5903 2565 5929 2621
rect 5985 2565 6011 2621
rect 6067 2565 6093 2621
rect 6149 2565 6175 2621
rect 6231 2565 6257 2621
rect 6313 2565 6339 2621
rect 6395 2565 6421 2621
rect 6477 2565 6503 2621
rect 6559 2565 6585 2621
rect 6641 2565 6666 2621
rect 6722 2565 6747 2621
rect 6803 2565 6828 2621
rect 6884 2565 6909 2621
rect 6965 2565 6990 2621
rect 7046 2565 7071 2621
rect 7127 2565 7152 2621
rect 7208 2565 7233 2621
rect 7289 2565 7314 2621
rect 7370 2565 7379 2621
rect 5179 2541 7379 2565
rect 5179 2485 5191 2541
rect 5247 2485 5273 2541
rect 5329 2485 5355 2541
rect 5411 2485 5437 2541
rect 5493 2485 5519 2541
rect 5575 2485 5601 2541
rect 5657 2485 5683 2541
rect 5739 2485 5765 2541
rect 5821 2485 5847 2541
rect 5903 2485 5929 2541
rect 5985 2485 6011 2541
rect 6067 2485 6093 2541
rect 6149 2485 6175 2541
rect 6231 2485 6257 2541
rect 6313 2485 6339 2541
rect 6395 2485 6421 2541
rect 6477 2485 6503 2541
rect 6559 2485 6585 2541
rect 6641 2485 6666 2541
rect 6722 2485 6747 2541
rect 6803 2485 6828 2541
rect 6884 2485 6909 2541
rect 6965 2485 6990 2541
rect 7046 2485 7071 2541
rect 7127 2485 7152 2541
rect 7208 2485 7233 2541
rect 7289 2485 7314 2541
rect 7370 2485 7379 2541
rect 5179 0 7379 2485
rect 7578 19973 7640 20029
rect 7696 19973 7726 20029
rect 7782 19973 7812 20029
rect 7868 19973 7898 20029
rect 7954 19973 7984 20029
rect 8040 19973 8070 20029
rect 8126 19973 8156 20029
rect 8212 19973 8242 20029
rect 8298 19973 8327 20029
rect 8383 19973 8412 20029
rect 8468 19973 8497 20029
rect 8553 19973 8596 20029
tri 8596 19973 8652 20029 sw
tri 8997 19973 9053 20029 se
rect 9053 19973 9079 20029
rect 9135 19973 9170 20029
rect 9226 19973 9260 20029
rect 9316 19973 9350 20029
rect 9406 19973 9440 20029
rect 9496 19973 9530 20029
rect 9586 19973 9620 20029
rect 9676 19973 9710 20029
rect 9766 19973 10208 20029
rect 7578 19949 8652 19973
tri 8652 19949 8676 19973 sw
tri 8973 19949 8997 19973 se
rect 8997 19949 10208 19973
rect 7578 19893 7640 19949
rect 7696 19893 7726 19949
rect 7782 19893 7812 19949
rect 7868 19893 7898 19949
rect 7954 19893 7984 19949
rect 8040 19893 8070 19949
rect 8126 19893 8156 19949
rect 8212 19893 8242 19949
rect 8298 19893 8327 19949
rect 8383 19893 8412 19949
rect 8468 19893 8497 19949
rect 8553 19901 8676 19949
tri 8676 19901 8724 19949 sw
tri 8925 19901 8973 19949 se
rect 8973 19901 9079 19949
rect 8553 19893 9079 19901
rect 9135 19893 9170 19949
rect 9226 19893 9260 19949
rect 9316 19893 9350 19949
rect 9406 19893 9440 19949
rect 9496 19893 9530 19949
rect 9586 19893 9620 19949
rect 9676 19893 9710 19949
rect 9766 19893 10208 19949
tri 10208 19943 10311 20046 nw
rect 7578 19869 10208 19893
rect 7578 19813 7640 19869
rect 7696 19813 7726 19869
rect 7782 19813 7812 19869
rect 7868 19813 7898 19869
rect 7954 19813 7984 19869
rect 8040 19813 8070 19869
rect 8126 19813 8156 19869
rect 8212 19813 8242 19869
rect 8298 19813 8327 19869
rect 8383 19813 8412 19869
rect 8468 19813 8497 19869
rect 8553 19813 9079 19869
rect 9135 19813 9170 19869
rect 9226 19813 9260 19869
rect 9316 19813 9350 19869
rect 9406 19813 9440 19869
rect 9496 19813 9530 19869
rect 9586 19813 9620 19869
rect 9676 19813 9710 19869
rect 9766 19813 10208 19869
rect 7578 19789 10208 19813
rect 7578 19733 7640 19789
rect 7696 19733 7726 19789
rect 7782 19733 7812 19789
rect 7868 19733 7898 19789
rect 7954 19733 7984 19789
rect 8040 19733 8070 19789
rect 8126 19733 8156 19789
rect 8212 19733 8242 19789
rect 8298 19733 8327 19789
rect 8383 19733 8412 19789
rect 8468 19733 8497 19789
rect 8553 19733 9079 19789
rect 9135 19733 9170 19789
rect 9226 19733 9260 19789
rect 9316 19733 9350 19789
rect 9406 19733 9440 19789
rect 9496 19733 9530 19789
rect 9586 19733 9620 19789
rect 9676 19733 9710 19789
rect 9766 19733 10208 19789
rect 7578 19709 10208 19733
rect 7578 19653 7640 19709
rect 7696 19653 7726 19709
rect 7782 19653 7812 19709
rect 7868 19653 7898 19709
rect 7954 19653 7984 19709
rect 8040 19653 8070 19709
rect 8126 19653 8156 19709
rect 8212 19653 8242 19709
rect 8298 19653 8327 19709
rect 8383 19653 8412 19709
rect 8468 19653 8497 19709
rect 8553 19653 9079 19709
rect 9135 19653 9170 19709
rect 9226 19653 9260 19709
rect 9316 19653 9350 19709
rect 9406 19653 9440 19709
rect 9496 19653 9530 19709
rect 9586 19653 9620 19709
rect 9676 19653 9710 19709
rect 9766 19660 10208 19709
rect 9766 19653 9778 19660
rect 7578 19629 9778 19653
rect 7578 19573 7640 19629
rect 7696 19573 7726 19629
rect 7782 19573 7812 19629
rect 7868 19573 7898 19629
rect 7954 19573 7984 19629
rect 8040 19573 8070 19629
rect 8126 19573 8156 19629
rect 8212 19573 8242 19629
rect 8298 19573 8327 19629
rect 8383 19573 8412 19629
rect 8468 19573 8497 19629
rect 8553 19573 9079 19629
rect 9135 19573 9170 19629
rect 9226 19573 9260 19629
rect 9316 19573 9350 19629
rect 9406 19573 9440 19629
rect 9496 19573 9530 19629
rect 9586 19573 9620 19629
rect 9676 19573 9710 19629
rect 9766 19573 9778 19629
rect 7578 19549 9778 19573
rect 7578 19493 7640 19549
rect 7696 19493 7726 19549
rect 7782 19493 7812 19549
rect 7868 19493 7898 19549
rect 7954 19493 7984 19549
rect 8040 19493 8070 19549
rect 8126 19493 8156 19549
rect 8212 19493 8242 19549
rect 8298 19493 8327 19549
rect 8383 19493 8412 19549
rect 8468 19493 8497 19549
rect 8553 19493 9079 19549
rect 9135 19493 9170 19549
rect 9226 19493 9260 19549
rect 9316 19493 9350 19549
rect 9406 19493 9440 19549
rect 9496 19493 9530 19549
rect 9586 19493 9620 19549
rect 9676 19493 9710 19549
rect 9766 19493 9778 19549
rect 7578 19469 9778 19493
rect 7578 19413 7640 19469
rect 7696 19413 7726 19469
rect 7782 19413 7812 19469
rect 7868 19413 7898 19469
rect 7954 19413 7984 19469
rect 8040 19413 8070 19469
rect 8126 19413 8156 19469
rect 8212 19413 8242 19469
rect 8298 19413 8327 19469
rect 8383 19413 8412 19469
rect 8468 19413 8497 19469
rect 8553 19413 9079 19469
rect 9135 19413 9170 19469
rect 9226 19413 9260 19469
rect 9316 19413 9350 19469
rect 9406 19413 9440 19469
rect 9496 19413 9530 19469
rect 9586 19413 9620 19469
rect 9676 19413 9710 19469
rect 9766 19413 9778 19469
rect 7578 19389 9778 19413
rect 7578 19333 7640 19389
rect 7696 19333 7726 19389
rect 7782 19333 7812 19389
rect 7868 19333 7898 19389
rect 7954 19333 7984 19389
rect 8040 19333 8070 19389
rect 8126 19333 8156 19389
rect 8212 19333 8242 19389
rect 8298 19333 8327 19389
rect 8383 19333 8412 19389
rect 8468 19333 8497 19389
rect 8553 19333 9079 19389
rect 9135 19333 9170 19389
rect 9226 19333 9260 19389
rect 9316 19333 9350 19389
rect 9406 19333 9440 19389
rect 9496 19333 9530 19389
rect 9586 19333 9620 19389
rect 9676 19333 9710 19389
rect 9766 19333 9778 19389
rect 7578 19309 9778 19333
rect 7578 19253 7640 19309
rect 7696 19253 7726 19309
rect 7782 19253 7812 19309
rect 7868 19253 7898 19309
rect 7954 19253 7984 19309
rect 8040 19253 8070 19309
rect 8126 19253 8156 19309
rect 8212 19253 8242 19309
rect 8298 19253 8327 19309
rect 8383 19253 8412 19309
rect 8468 19253 8497 19309
rect 8553 19253 9079 19309
rect 9135 19253 9170 19309
rect 9226 19253 9260 19309
rect 9316 19253 9350 19309
rect 9406 19253 9440 19309
rect 9496 19253 9530 19309
rect 9586 19253 9620 19309
rect 9676 19253 9710 19309
rect 9766 19253 9778 19309
rect 7578 19229 9778 19253
tri 9778 19230 10208 19660 nw
rect 7578 19173 7640 19229
rect 7696 19173 7726 19229
rect 7782 19173 7812 19229
rect 7868 19173 7898 19229
rect 7954 19173 7984 19229
rect 8040 19173 8070 19229
rect 8126 19173 8156 19229
rect 8212 19173 8242 19229
rect 8298 19173 8327 19229
rect 8383 19173 8412 19229
rect 8468 19173 8497 19229
rect 8553 19173 9079 19229
rect 9135 19173 9170 19229
rect 9226 19173 9260 19229
rect 9316 19173 9350 19229
rect 9406 19173 9440 19229
rect 9496 19173 9530 19229
rect 9586 19173 9620 19229
rect 9676 19173 9710 19229
rect 9766 19173 9778 19229
rect 7578 19149 9778 19173
rect 7578 19093 7640 19149
rect 7696 19093 7726 19149
rect 7782 19093 7812 19149
rect 7868 19093 7898 19149
rect 7954 19093 7984 19149
rect 8040 19093 8070 19149
rect 8126 19093 8156 19149
rect 8212 19093 8242 19149
rect 8298 19093 8327 19149
rect 8383 19093 8412 19149
rect 8468 19093 8497 19149
rect 8553 19093 9079 19149
rect 9135 19093 9170 19149
rect 9226 19093 9260 19149
rect 9316 19093 9350 19149
rect 9406 19093 9440 19149
rect 9496 19093 9530 19149
rect 9586 19093 9620 19149
rect 9676 19093 9710 19149
rect 9766 19093 9778 19149
rect 7578 19069 9778 19093
rect 7578 19013 7640 19069
rect 7696 19013 7726 19069
rect 7782 19013 7812 19069
rect 7868 19013 7898 19069
rect 7954 19013 7984 19069
rect 8040 19013 8070 19069
rect 8126 19013 8156 19069
rect 8212 19013 8242 19069
rect 8298 19013 8327 19069
rect 8383 19013 8412 19069
rect 8468 19013 8497 19069
rect 8553 19013 9079 19069
rect 9135 19013 9170 19069
rect 9226 19013 9260 19069
rect 9316 19013 9350 19069
rect 9406 19013 9440 19069
rect 9496 19013 9530 19069
rect 9586 19013 9620 19069
rect 9676 19013 9710 19069
rect 9766 19013 9778 19069
rect 7578 18989 9778 19013
rect 7578 18933 7640 18989
rect 7696 18933 7726 18989
rect 7782 18933 7812 18989
rect 7868 18933 7898 18989
rect 7954 18933 7984 18989
rect 8040 18933 8070 18989
rect 8126 18933 8156 18989
rect 8212 18933 8242 18989
rect 8298 18933 8327 18989
rect 8383 18933 8412 18989
rect 8468 18933 8497 18989
rect 8553 18933 9079 18989
rect 9135 18933 9170 18989
rect 9226 18933 9260 18989
rect 9316 18933 9350 18989
rect 9406 18933 9440 18989
rect 9496 18933 9530 18989
rect 9586 18933 9620 18989
rect 9676 18933 9710 18989
rect 9766 18933 9778 18989
rect 7578 18909 9778 18933
rect 7578 18853 7640 18909
rect 7696 18853 7726 18909
rect 7782 18853 7812 18909
rect 7868 18853 7898 18909
rect 7954 18853 7984 18909
rect 8040 18853 8070 18909
rect 8126 18853 8156 18909
rect 8212 18853 8242 18909
rect 8298 18853 8327 18909
rect 8383 18853 8412 18909
rect 8468 18853 8497 18909
rect 8553 18853 9079 18909
rect 9135 18853 9170 18909
rect 9226 18853 9260 18909
rect 9316 18853 9350 18909
rect 9406 18853 9440 18909
rect 9496 18853 9530 18909
rect 9586 18853 9620 18909
rect 9676 18853 9710 18909
rect 9766 18853 9778 18909
rect 7578 18829 9778 18853
rect 7578 18773 7640 18829
rect 7696 18773 7726 18829
rect 7782 18773 7812 18829
rect 7868 18773 7898 18829
rect 7954 18773 7984 18829
rect 8040 18773 8070 18829
rect 8126 18773 8156 18829
rect 8212 18773 8242 18829
rect 8298 18773 8327 18829
rect 8383 18773 8412 18829
rect 8468 18773 8497 18829
rect 8553 18773 9079 18829
rect 9135 18773 9170 18829
rect 9226 18773 9260 18829
rect 9316 18773 9350 18829
rect 9406 18773 9440 18829
rect 9496 18773 9530 18829
rect 9586 18773 9620 18829
rect 9676 18773 9710 18829
rect 9766 18773 9778 18829
rect 7578 18749 9778 18773
rect 7578 18693 7640 18749
rect 7696 18693 7726 18749
rect 7782 18693 7812 18749
rect 7868 18693 7898 18749
rect 7954 18693 7984 18749
rect 8040 18693 8070 18749
rect 8126 18693 8156 18749
rect 8212 18693 8242 18749
rect 8298 18693 8327 18749
rect 8383 18693 8412 18749
rect 8468 18693 8497 18749
rect 8553 18693 9079 18749
rect 9135 18693 9170 18749
rect 9226 18693 9260 18749
rect 9316 18693 9350 18749
rect 9406 18693 9440 18749
rect 9496 18693 9530 18749
rect 9586 18693 9620 18749
rect 9676 18693 9710 18749
rect 9766 18693 9778 18749
rect 7578 15829 9778 18693
rect 7578 15773 7587 15829
rect 7643 15773 7669 15829
rect 7725 15773 7751 15829
rect 7807 15773 7833 15829
rect 7889 15773 7915 15829
rect 7971 15773 7997 15829
rect 8053 15773 8079 15829
rect 8135 15773 8161 15829
rect 8217 15773 8243 15829
rect 8299 15773 8325 15829
rect 8381 15773 8407 15829
rect 8463 15773 8489 15829
rect 8545 15773 8571 15829
rect 8627 15773 8653 15829
rect 8709 15773 8735 15829
rect 8791 15773 8817 15829
rect 8873 15773 8899 15829
rect 8955 15773 8981 15829
rect 9037 15773 9063 15829
rect 9119 15773 9145 15829
rect 9201 15773 9227 15829
rect 9283 15773 9308 15829
rect 9364 15773 9389 15829
rect 9445 15773 9470 15829
rect 9526 15773 9551 15829
rect 9607 15773 9632 15829
rect 9688 15773 9713 15829
rect 9769 15773 9778 15829
rect 7578 15749 9778 15773
rect 7578 15693 7587 15749
rect 7643 15693 7669 15749
rect 7725 15693 7751 15749
rect 7807 15693 7833 15749
rect 7889 15693 7915 15749
rect 7971 15693 7997 15749
rect 8053 15693 8079 15749
rect 8135 15693 8161 15749
rect 8217 15693 8243 15749
rect 8299 15693 8325 15749
rect 8381 15693 8407 15749
rect 8463 15693 8489 15749
rect 8545 15693 8571 15749
rect 8627 15693 8653 15749
rect 8709 15693 8735 15749
rect 8791 15693 8817 15749
rect 8873 15693 8899 15749
rect 8955 15693 8981 15749
rect 9037 15693 9063 15749
rect 9119 15693 9145 15749
rect 9201 15693 9227 15749
rect 9283 15693 9308 15749
rect 9364 15693 9389 15749
rect 9445 15693 9470 15749
rect 9526 15693 9551 15749
rect 9607 15693 9632 15749
rect 9688 15693 9713 15749
rect 9769 15693 9778 15749
rect 7578 15669 9778 15693
rect 7578 15613 7587 15669
rect 7643 15613 7669 15669
rect 7725 15613 7751 15669
rect 7807 15613 7833 15669
rect 7889 15613 7915 15669
rect 7971 15613 7997 15669
rect 8053 15613 8079 15669
rect 8135 15613 8161 15669
rect 8217 15613 8243 15669
rect 8299 15613 8325 15669
rect 8381 15613 8407 15669
rect 8463 15613 8489 15669
rect 8545 15613 8571 15669
rect 8627 15613 8653 15669
rect 8709 15613 8735 15669
rect 8791 15613 8817 15669
rect 8873 15613 8899 15669
rect 8955 15613 8981 15669
rect 9037 15613 9063 15669
rect 9119 15613 9145 15669
rect 9201 15613 9227 15669
rect 9283 15613 9308 15669
rect 9364 15613 9389 15669
rect 9445 15613 9470 15669
rect 9526 15613 9551 15669
rect 9607 15613 9632 15669
rect 9688 15613 9713 15669
rect 9769 15613 9778 15669
rect 7578 15589 9778 15613
rect 7578 15533 7587 15589
rect 7643 15533 7669 15589
rect 7725 15533 7751 15589
rect 7807 15533 7833 15589
rect 7889 15533 7915 15589
rect 7971 15533 7997 15589
rect 8053 15533 8079 15589
rect 8135 15533 8161 15589
rect 8217 15533 8243 15589
rect 8299 15533 8325 15589
rect 8381 15533 8407 15589
rect 8463 15533 8489 15589
rect 8545 15533 8571 15589
rect 8627 15533 8653 15589
rect 8709 15533 8735 15589
rect 8791 15533 8817 15589
rect 8873 15533 8899 15589
rect 8955 15533 8981 15589
rect 9037 15533 9063 15589
rect 9119 15533 9145 15589
rect 9201 15533 9227 15589
rect 9283 15533 9308 15589
rect 9364 15533 9389 15589
rect 9445 15533 9470 15589
rect 9526 15533 9551 15589
rect 9607 15533 9632 15589
rect 9688 15533 9713 15589
rect 9769 15533 9778 15589
rect 7578 15509 9778 15533
rect 7578 15453 7587 15509
rect 7643 15453 7669 15509
rect 7725 15453 7751 15509
rect 7807 15453 7833 15509
rect 7889 15453 7915 15509
rect 7971 15453 7997 15509
rect 8053 15453 8079 15509
rect 8135 15453 8161 15509
rect 8217 15453 8243 15509
rect 8299 15453 8325 15509
rect 8381 15453 8407 15509
rect 8463 15453 8489 15509
rect 8545 15453 8571 15509
rect 8627 15453 8653 15509
rect 8709 15453 8735 15509
rect 8791 15453 8817 15509
rect 8873 15453 8899 15509
rect 8955 15453 8981 15509
rect 9037 15453 9063 15509
rect 9119 15453 9145 15509
rect 9201 15453 9227 15509
rect 9283 15453 9308 15509
rect 9364 15453 9389 15509
rect 9445 15453 9470 15509
rect 9526 15453 9551 15509
rect 9607 15453 9632 15509
rect 9688 15453 9713 15509
rect 9769 15453 9778 15509
rect 7578 15429 9778 15453
rect 7578 15373 7587 15429
rect 7643 15373 7669 15429
rect 7725 15373 7751 15429
rect 7807 15373 7833 15429
rect 7889 15373 7915 15429
rect 7971 15373 7997 15429
rect 8053 15373 8079 15429
rect 8135 15373 8161 15429
rect 8217 15373 8243 15429
rect 8299 15373 8325 15429
rect 8381 15373 8407 15429
rect 8463 15373 8489 15429
rect 8545 15373 8571 15429
rect 8627 15373 8653 15429
rect 8709 15373 8735 15429
rect 8791 15373 8817 15429
rect 8873 15373 8899 15429
rect 8955 15373 8981 15429
rect 9037 15373 9063 15429
rect 9119 15373 9145 15429
rect 9201 15373 9227 15429
rect 9283 15373 9308 15429
rect 9364 15373 9389 15429
rect 9445 15373 9470 15429
rect 9526 15373 9551 15429
rect 9607 15373 9632 15429
rect 9688 15373 9713 15429
rect 9769 15373 9778 15429
rect 7578 15349 9778 15373
rect 7578 15293 7587 15349
rect 7643 15293 7669 15349
rect 7725 15293 7751 15349
rect 7807 15293 7833 15349
rect 7889 15293 7915 15349
rect 7971 15293 7997 15349
rect 8053 15293 8079 15349
rect 8135 15293 8161 15349
rect 8217 15293 8243 15349
rect 8299 15293 8325 15349
rect 8381 15293 8407 15349
rect 8463 15293 8489 15349
rect 8545 15293 8571 15349
rect 8627 15293 8653 15349
rect 8709 15293 8735 15349
rect 8791 15293 8817 15349
rect 8873 15293 8899 15349
rect 8955 15293 8981 15349
rect 9037 15293 9063 15349
rect 9119 15293 9145 15349
rect 9201 15293 9227 15349
rect 9283 15293 9308 15349
rect 9364 15293 9389 15349
rect 9445 15293 9470 15349
rect 9526 15293 9551 15349
rect 9607 15293 9632 15349
rect 9688 15293 9713 15349
rect 9769 15293 9778 15349
rect 7578 15269 9778 15293
rect 7578 15213 7587 15269
rect 7643 15213 7669 15269
rect 7725 15213 7751 15269
rect 7807 15213 7833 15269
rect 7889 15213 7915 15269
rect 7971 15213 7997 15269
rect 8053 15213 8079 15269
rect 8135 15213 8161 15269
rect 8217 15213 8243 15269
rect 8299 15213 8325 15269
rect 8381 15213 8407 15269
rect 8463 15213 8489 15269
rect 8545 15213 8571 15269
rect 8627 15213 8653 15269
rect 8709 15213 8735 15269
rect 8791 15213 8817 15269
rect 8873 15213 8899 15269
rect 8955 15213 8981 15269
rect 9037 15213 9063 15269
rect 9119 15213 9145 15269
rect 9201 15213 9227 15269
rect 9283 15213 9308 15269
rect 9364 15213 9389 15269
rect 9445 15213 9470 15269
rect 9526 15213 9551 15269
rect 9607 15213 9632 15269
rect 9688 15213 9713 15269
rect 9769 15213 9778 15269
rect 7578 15189 9778 15213
rect 7578 15133 7587 15189
rect 7643 15133 7669 15189
rect 7725 15133 7751 15189
rect 7807 15133 7833 15189
rect 7889 15133 7915 15189
rect 7971 15133 7997 15189
rect 8053 15133 8079 15189
rect 8135 15133 8161 15189
rect 8217 15133 8243 15189
rect 8299 15133 8325 15189
rect 8381 15133 8407 15189
rect 8463 15133 8489 15189
rect 8545 15133 8571 15189
rect 8627 15133 8653 15189
rect 8709 15133 8735 15189
rect 8791 15133 8817 15189
rect 8873 15133 8899 15189
rect 8955 15133 8981 15189
rect 9037 15133 9063 15189
rect 9119 15133 9145 15189
rect 9201 15133 9227 15189
rect 9283 15133 9308 15189
rect 9364 15133 9389 15189
rect 9445 15133 9470 15189
rect 9526 15133 9551 15189
rect 9607 15133 9632 15189
rect 9688 15133 9713 15189
rect 9769 15133 9778 15189
rect 7578 15109 9778 15133
rect 7578 15053 7587 15109
rect 7643 15053 7669 15109
rect 7725 15053 7751 15109
rect 7807 15053 7833 15109
rect 7889 15053 7915 15109
rect 7971 15053 7997 15109
rect 8053 15053 8079 15109
rect 8135 15053 8161 15109
rect 8217 15053 8243 15109
rect 8299 15053 8325 15109
rect 8381 15053 8407 15109
rect 8463 15053 8489 15109
rect 8545 15053 8571 15109
rect 8627 15053 8653 15109
rect 8709 15053 8735 15109
rect 8791 15053 8817 15109
rect 8873 15053 8899 15109
rect 8955 15053 8981 15109
rect 9037 15053 9063 15109
rect 9119 15053 9145 15109
rect 9201 15053 9227 15109
rect 9283 15053 9308 15109
rect 9364 15053 9389 15109
rect 9445 15053 9470 15109
rect 9526 15053 9551 15109
rect 9607 15053 9632 15109
rect 9688 15053 9713 15109
rect 9769 15053 9778 15109
rect 7578 15029 9778 15053
rect 7578 14973 7587 15029
rect 7643 14973 7669 15029
rect 7725 14973 7751 15029
rect 7807 14973 7833 15029
rect 7889 14973 7915 15029
rect 7971 14973 7997 15029
rect 8053 14973 8079 15029
rect 8135 14973 8161 15029
rect 8217 14973 8243 15029
rect 8299 14973 8325 15029
rect 8381 14973 8407 15029
rect 8463 14973 8489 15029
rect 8545 14973 8571 15029
rect 8627 14973 8653 15029
rect 8709 14973 8735 15029
rect 8791 14973 8817 15029
rect 8873 14973 8899 15029
rect 8955 14973 8981 15029
rect 9037 14973 9063 15029
rect 9119 14973 9145 15029
rect 9201 14973 9227 15029
rect 9283 14973 9308 15029
rect 9364 14973 9389 15029
rect 9445 14973 9470 15029
rect 9526 14973 9551 15029
rect 9607 14973 9632 15029
rect 9688 14973 9713 15029
rect 9769 14973 9778 15029
rect 7578 14949 9778 14973
rect 7578 14893 7587 14949
rect 7643 14893 7669 14949
rect 7725 14893 7751 14949
rect 7807 14893 7833 14949
rect 7889 14893 7915 14949
rect 7971 14893 7997 14949
rect 8053 14893 8079 14949
rect 8135 14893 8161 14949
rect 8217 14893 8243 14949
rect 8299 14893 8325 14949
rect 8381 14893 8407 14949
rect 8463 14893 8489 14949
rect 8545 14893 8571 14949
rect 8627 14893 8653 14949
rect 8709 14893 8735 14949
rect 8791 14893 8817 14949
rect 8873 14893 8899 14949
rect 8955 14893 8981 14949
rect 9037 14893 9063 14949
rect 9119 14893 9145 14949
rect 9201 14893 9227 14949
rect 9283 14893 9308 14949
rect 9364 14893 9389 14949
rect 9445 14893 9470 14949
rect 9526 14893 9551 14949
rect 9607 14893 9632 14949
rect 9688 14893 9713 14949
rect 9769 14893 9778 14949
rect 7578 14869 9778 14893
rect 7578 14813 7587 14869
rect 7643 14813 7669 14869
rect 7725 14813 7751 14869
rect 7807 14813 7833 14869
rect 7889 14813 7915 14869
rect 7971 14813 7997 14869
rect 8053 14813 8079 14869
rect 8135 14813 8161 14869
rect 8217 14813 8243 14869
rect 8299 14813 8325 14869
rect 8381 14813 8407 14869
rect 8463 14813 8489 14869
rect 8545 14813 8571 14869
rect 8627 14813 8653 14869
rect 8709 14813 8735 14869
rect 8791 14813 8817 14869
rect 8873 14813 8899 14869
rect 8955 14813 8981 14869
rect 9037 14813 9063 14869
rect 9119 14813 9145 14869
rect 9201 14813 9227 14869
rect 9283 14813 9308 14869
rect 9364 14813 9389 14869
rect 9445 14813 9470 14869
rect 9526 14813 9551 14869
rect 9607 14813 9632 14869
rect 9688 14813 9713 14869
rect 9769 14813 9778 14869
rect 7578 14789 9778 14813
rect 7578 14733 7587 14789
rect 7643 14733 7669 14789
rect 7725 14733 7751 14789
rect 7807 14733 7833 14789
rect 7889 14733 7915 14789
rect 7971 14733 7997 14789
rect 8053 14733 8079 14789
rect 8135 14733 8161 14789
rect 8217 14733 8243 14789
rect 8299 14733 8325 14789
rect 8381 14733 8407 14789
rect 8463 14733 8489 14789
rect 8545 14733 8571 14789
rect 8627 14733 8653 14789
rect 8709 14733 8735 14789
rect 8791 14733 8817 14789
rect 8873 14733 8899 14789
rect 8955 14733 8981 14789
rect 9037 14733 9063 14789
rect 9119 14733 9145 14789
rect 9201 14733 9227 14789
rect 9283 14733 9308 14789
rect 9364 14733 9389 14789
rect 9445 14733 9470 14789
rect 9526 14733 9551 14789
rect 9607 14733 9632 14789
rect 9688 14733 9713 14789
rect 9769 14733 9778 14789
rect 7578 14709 9778 14733
rect 7578 14653 7587 14709
rect 7643 14653 7669 14709
rect 7725 14653 7751 14709
rect 7807 14653 7833 14709
rect 7889 14653 7915 14709
rect 7971 14653 7997 14709
rect 8053 14653 8079 14709
rect 8135 14653 8161 14709
rect 8217 14653 8243 14709
rect 8299 14653 8325 14709
rect 8381 14653 8407 14709
rect 8463 14653 8489 14709
rect 8545 14653 8571 14709
rect 8627 14653 8653 14709
rect 8709 14653 8735 14709
rect 8791 14653 8817 14709
rect 8873 14653 8899 14709
rect 8955 14653 8981 14709
rect 9037 14653 9063 14709
rect 9119 14653 9145 14709
rect 9201 14653 9227 14709
rect 9283 14653 9308 14709
rect 9364 14653 9389 14709
rect 9445 14653 9470 14709
rect 9526 14653 9551 14709
rect 9607 14653 9632 14709
rect 9688 14653 9713 14709
rect 9769 14653 9778 14709
rect 7578 14629 9778 14653
rect 7578 14573 7587 14629
rect 7643 14573 7669 14629
rect 7725 14573 7751 14629
rect 7807 14573 7833 14629
rect 7889 14573 7915 14629
rect 7971 14573 7997 14629
rect 8053 14573 8079 14629
rect 8135 14573 8161 14629
rect 8217 14573 8243 14629
rect 8299 14573 8325 14629
rect 8381 14573 8407 14629
rect 8463 14573 8489 14629
rect 8545 14573 8571 14629
rect 8627 14573 8653 14629
rect 8709 14573 8735 14629
rect 8791 14573 8817 14629
rect 8873 14573 8899 14629
rect 8955 14573 8981 14629
rect 9037 14573 9063 14629
rect 9119 14573 9145 14629
rect 9201 14573 9227 14629
rect 9283 14573 9308 14629
rect 9364 14573 9389 14629
rect 9445 14573 9470 14629
rect 9526 14573 9551 14629
rect 9607 14573 9632 14629
rect 9688 14573 9713 14629
rect 9769 14573 9778 14629
rect 7578 14549 9778 14573
rect 7578 14493 7587 14549
rect 7643 14493 7669 14549
rect 7725 14493 7751 14549
rect 7807 14493 7833 14549
rect 7889 14493 7915 14549
rect 7971 14493 7997 14549
rect 8053 14493 8079 14549
rect 8135 14493 8161 14549
rect 8217 14493 8243 14549
rect 8299 14493 8325 14549
rect 8381 14493 8407 14549
rect 8463 14493 8489 14549
rect 8545 14493 8571 14549
rect 8627 14493 8653 14549
rect 8709 14493 8735 14549
rect 8791 14493 8817 14549
rect 8873 14493 8899 14549
rect 8955 14493 8981 14549
rect 9037 14493 9063 14549
rect 9119 14493 9145 14549
rect 9201 14493 9227 14549
rect 9283 14493 9308 14549
rect 9364 14493 9389 14549
rect 9445 14493 9470 14549
rect 9526 14493 9551 14549
rect 9607 14493 9632 14549
rect 9688 14493 9713 14549
rect 9769 14493 9778 14549
rect 7578 14469 9778 14493
rect 7578 14413 7587 14469
rect 7643 14413 7669 14469
rect 7725 14413 7751 14469
rect 7807 14413 7833 14469
rect 7889 14413 7915 14469
rect 7971 14413 7997 14469
rect 8053 14413 8079 14469
rect 8135 14413 8161 14469
rect 8217 14413 8243 14469
rect 8299 14413 8325 14469
rect 8381 14413 8407 14469
rect 8463 14413 8489 14469
rect 8545 14413 8571 14469
rect 8627 14413 8653 14469
rect 8709 14413 8735 14469
rect 8791 14413 8817 14469
rect 8873 14413 8899 14469
rect 8955 14413 8981 14469
rect 9037 14413 9063 14469
rect 9119 14413 9145 14469
rect 9201 14413 9227 14469
rect 9283 14413 9308 14469
rect 9364 14413 9389 14469
rect 9445 14413 9470 14469
rect 9526 14413 9551 14469
rect 9607 14413 9632 14469
rect 9688 14413 9713 14469
rect 9769 14413 9778 14469
rect 7578 14389 9778 14413
rect 7578 14333 7587 14389
rect 7643 14333 7669 14389
rect 7725 14333 7751 14389
rect 7807 14333 7833 14389
rect 7889 14333 7915 14389
rect 7971 14333 7997 14389
rect 8053 14333 8079 14389
rect 8135 14333 8161 14389
rect 8217 14333 8243 14389
rect 8299 14333 8325 14389
rect 8381 14333 8407 14389
rect 8463 14333 8489 14389
rect 8545 14333 8571 14389
rect 8627 14333 8653 14389
rect 8709 14333 8735 14389
rect 8791 14333 8817 14389
rect 8873 14333 8899 14389
rect 8955 14333 8981 14389
rect 9037 14333 9063 14389
rect 9119 14333 9145 14389
rect 9201 14333 9227 14389
rect 9283 14333 9308 14389
rect 9364 14333 9389 14389
rect 9445 14333 9470 14389
rect 9526 14333 9551 14389
rect 9607 14333 9632 14389
rect 9688 14333 9713 14389
rect 9769 14333 9778 14389
rect 7578 14309 9778 14333
rect 7578 14253 7587 14309
rect 7643 14253 7669 14309
rect 7725 14253 7751 14309
rect 7807 14253 7833 14309
rect 7889 14253 7915 14309
rect 7971 14253 7997 14309
rect 8053 14253 8079 14309
rect 8135 14253 8161 14309
rect 8217 14253 8243 14309
rect 8299 14253 8325 14309
rect 8381 14253 8407 14309
rect 8463 14253 8489 14309
rect 8545 14253 8571 14309
rect 8627 14253 8653 14309
rect 8709 14253 8735 14309
rect 8791 14253 8817 14309
rect 8873 14253 8899 14309
rect 8955 14253 8981 14309
rect 9037 14253 9063 14309
rect 9119 14253 9145 14309
rect 9201 14253 9227 14309
rect 9283 14253 9308 14309
rect 9364 14253 9389 14309
rect 9445 14253 9470 14309
rect 9526 14253 9551 14309
rect 9607 14253 9632 14309
rect 9688 14253 9713 14309
rect 9769 14253 9778 14309
rect 7578 14229 9778 14253
rect 7578 14173 7587 14229
rect 7643 14173 7669 14229
rect 7725 14173 7751 14229
rect 7807 14173 7833 14229
rect 7889 14173 7915 14229
rect 7971 14173 7997 14229
rect 8053 14173 8079 14229
rect 8135 14173 8161 14229
rect 8217 14173 8243 14229
rect 8299 14173 8325 14229
rect 8381 14173 8407 14229
rect 8463 14173 8489 14229
rect 8545 14173 8571 14229
rect 8627 14173 8653 14229
rect 8709 14173 8735 14229
rect 8791 14173 8817 14229
rect 8873 14173 8899 14229
rect 8955 14173 8981 14229
rect 9037 14173 9063 14229
rect 9119 14173 9145 14229
rect 9201 14173 9227 14229
rect 9283 14173 9308 14229
rect 9364 14173 9389 14229
rect 9445 14173 9470 14229
rect 9526 14173 9551 14229
rect 9607 14173 9632 14229
rect 9688 14173 9713 14229
rect 9769 14173 9778 14229
rect 7578 14149 9778 14173
rect 7578 14093 7587 14149
rect 7643 14093 7669 14149
rect 7725 14093 7751 14149
rect 7807 14093 7833 14149
rect 7889 14093 7915 14149
rect 7971 14093 7997 14149
rect 8053 14093 8079 14149
rect 8135 14093 8161 14149
rect 8217 14093 8243 14149
rect 8299 14093 8325 14149
rect 8381 14093 8407 14149
rect 8463 14093 8489 14149
rect 8545 14093 8571 14149
rect 8627 14093 8653 14149
rect 8709 14093 8735 14149
rect 8791 14093 8817 14149
rect 8873 14093 8899 14149
rect 8955 14093 8981 14149
rect 9037 14093 9063 14149
rect 9119 14093 9145 14149
rect 9201 14093 9227 14149
rect 9283 14093 9308 14149
rect 9364 14093 9389 14149
rect 9445 14093 9470 14149
rect 9526 14093 9551 14149
rect 9607 14093 9632 14149
rect 9688 14093 9713 14149
rect 9769 14093 9778 14149
rect 7578 11229 9778 14093
rect 7578 11173 7587 11229
rect 7643 11173 7669 11229
rect 7725 11173 7751 11229
rect 7807 11173 7833 11229
rect 7889 11173 7915 11229
rect 7971 11173 7997 11229
rect 8053 11173 8079 11229
rect 8135 11173 8161 11229
rect 8217 11173 8243 11229
rect 8299 11173 8325 11229
rect 8381 11173 8407 11229
rect 8463 11173 8489 11229
rect 8545 11173 8571 11229
rect 8627 11173 8653 11229
rect 8709 11173 8735 11229
rect 8791 11173 8817 11229
rect 8873 11173 8899 11229
rect 8955 11173 8981 11229
rect 9037 11173 9063 11229
rect 9119 11173 9145 11229
rect 9201 11173 9227 11229
rect 9283 11173 9308 11229
rect 9364 11173 9389 11229
rect 9445 11173 9470 11229
rect 9526 11173 9551 11229
rect 9607 11173 9632 11229
rect 9688 11173 9713 11229
rect 9769 11173 9778 11229
rect 7578 11149 9778 11173
rect 7578 11093 7587 11149
rect 7643 11093 7669 11149
rect 7725 11093 7751 11149
rect 7807 11093 7833 11149
rect 7889 11093 7915 11149
rect 7971 11093 7997 11149
rect 8053 11093 8079 11149
rect 8135 11093 8161 11149
rect 8217 11093 8243 11149
rect 8299 11093 8325 11149
rect 8381 11093 8407 11149
rect 8463 11093 8489 11149
rect 8545 11093 8571 11149
rect 8627 11093 8653 11149
rect 8709 11093 8735 11149
rect 8791 11093 8817 11149
rect 8873 11093 8899 11149
rect 8955 11093 8981 11149
rect 9037 11093 9063 11149
rect 9119 11093 9145 11149
rect 9201 11093 9227 11149
rect 9283 11093 9308 11149
rect 9364 11093 9389 11149
rect 9445 11093 9470 11149
rect 9526 11093 9551 11149
rect 9607 11093 9632 11149
rect 9688 11093 9713 11149
rect 9769 11093 9778 11149
rect 7578 11069 9778 11093
rect 7578 11013 7587 11069
rect 7643 11013 7669 11069
rect 7725 11013 7751 11069
rect 7807 11013 7833 11069
rect 7889 11013 7915 11069
rect 7971 11013 7997 11069
rect 8053 11013 8079 11069
rect 8135 11013 8161 11069
rect 8217 11013 8243 11069
rect 8299 11013 8325 11069
rect 8381 11013 8407 11069
rect 8463 11013 8489 11069
rect 8545 11013 8571 11069
rect 8627 11013 8653 11069
rect 8709 11013 8735 11069
rect 8791 11013 8817 11069
rect 8873 11013 8899 11069
rect 8955 11013 8981 11069
rect 9037 11013 9063 11069
rect 9119 11013 9145 11069
rect 9201 11013 9227 11069
rect 9283 11013 9308 11069
rect 9364 11013 9389 11069
rect 9445 11013 9470 11069
rect 9526 11013 9551 11069
rect 9607 11013 9632 11069
rect 9688 11013 9713 11069
rect 9769 11013 9778 11069
rect 7578 10989 9778 11013
rect 7578 10933 7587 10989
rect 7643 10933 7669 10989
rect 7725 10933 7751 10989
rect 7807 10933 7833 10989
rect 7889 10933 7915 10989
rect 7971 10933 7997 10989
rect 8053 10933 8079 10989
rect 8135 10933 8161 10989
rect 8217 10933 8243 10989
rect 8299 10933 8325 10989
rect 8381 10933 8407 10989
rect 8463 10933 8489 10989
rect 8545 10933 8571 10989
rect 8627 10933 8653 10989
rect 8709 10933 8735 10989
rect 8791 10933 8817 10989
rect 8873 10933 8899 10989
rect 8955 10933 8981 10989
rect 9037 10933 9063 10989
rect 9119 10933 9145 10989
rect 9201 10933 9227 10989
rect 9283 10933 9308 10989
rect 9364 10933 9389 10989
rect 9445 10933 9470 10989
rect 9526 10933 9551 10989
rect 9607 10933 9632 10989
rect 9688 10933 9713 10989
rect 9769 10933 9778 10989
rect 7578 10909 9778 10933
rect 7578 10853 7587 10909
rect 7643 10853 7669 10909
rect 7725 10853 7751 10909
rect 7807 10853 7833 10909
rect 7889 10853 7915 10909
rect 7971 10853 7997 10909
rect 8053 10853 8079 10909
rect 8135 10853 8161 10909
rect 8217 10853 8243 10909
rect 8299 10853 8325 10909
rect 8381 10853 8407 10909
rect 8463 10853 8489 10909
rect 8545 10853 8571 10909
rect 8627 10853 8653 10909
rect 8709 10853 8735 10909
rect 8791 10853 8817 10909
rect 8873 10853 8899 10909
rect 8955 10853 8981 10909
rect 9037 10853 9063 10909
rect 9119 10853 9145 10909
rect 9201 10853 9227 10909
rect 9283 10853 9308 10909
rect 9364 10853 9389 10909
rect 9445 10853 9470 10909
rect 9526 10853 9551 10909
rect 9607 10853 9632 10909
rect 9688 10853 9713 10909
rect 9769 10853 9778 10909
rect 7578 10829 9778 10853
rect 7578 10773 7587 10829
rect 7643 10773 7669 10829
rect 7725 10773 7751 10829
rect 7807 10773 7833 10829
rect 7889 10773 7915 10829
rect 7971 10773 7997 10829
rect 8053 10773 8079 10829
rect 8135 10773 8161 10829
rect 8217 10773 8243 10829
rect 8299 10773 8325 10829
rect 8381 10773 8407 10829
rect 8463 10773 8489 10829
rect 8545 10773 8571 10829
rect 8627 10773 8653 10829
rect 8709 10773 8735 10829
rect 8791 10773 8817 10829
rect 8873 10773 8899 10829
rect 8955 10773 8981 10829
rect 9037 10773 9063 10829
rect 9119 10773 9145 10829
rect 9201 10773 9227 10829
rect 9283 10773 9308 10829
rect 9364 10773 9389 10829
rect 9445 10773 9470 10829
rect 9526 10773 9551 10829
rect 9607 10773 9632 10829
rect 9688 10773 9713 10829
rect 9769 10773 9778 10829
rect 7578 10749 9778 10773
rect 7578 10693 7587 10749
rect 7643 10693 7669 10749
rect 7725 10693 7751 10749
rect 7807 10693 7833 10749
rect 7889 10693 7915 10749
rect 7971 10693 7997 10749
rect 8053 10693 8079 10749
rect 8135 10693 8161 10749
rect 8217 10693 8243 10749
rect 8299 10693 8325 10749
rect 8381 10693 8407 10749
rect 8463 10693 8489 10749
rect 8545 10693 8571 10749
rect 8627 10693 8653 10749
rect 8709 10693 8735 10749
rect 8791 10693 8817 10749
rect 8873 10693 8899 10749
rect 8955 10693 8981 10749
rect 9037 10693 9063 10749
rect 9119 10693 9145 10749
rect 9201 10693 9227 10749
rect 9283 10693 9308 10749
rect 9364 10693 9389 10749
rect 9445 10693 9470 10749
rect 9526 10693 9551 10749
rect 9607 10693 9632 10749
rect 9688 10693 9713 10749
rect 9769 10693 9778 10749
rect 7578 10669 9778 10693
rect 7578 10613 7587 10669
rect 7643 10613 7669 10669
rect 7725 10613 7751 10669
rect 7807 10613 7833 10669
rect 7889 10613 7915 10669
rect 7971 10613 7997 10669
rect 8053 10613 8079 10669
rect 8135 10613 8161 10669
rect 8217 10613 8243 10669
rect 8299 10613 8325 10669
rect 8381 10613 8407 10669
rect 8463 10613 8489 10669
rect 8545 10613 8571 10669
rect 8627 10613 8653 10669
rect 8709 10613 8735 10669
rect 8791 10613 8817 10669
rect 8873 10613 8899 10669
rect 8955 10613 8981 10669
rect 9037 10613 9063 10669
rect 9119 10613 9145 10669
rect 9201 10613 9227 10669
rect 9283 10613 9308 10669
rect 9364 10613 9389 10669
rect 9445 10613 9470 10669
rect 9526 10613 9551 10669
rect 9607 10613 9632 10669
rect 9688 10613 9713 10669
rect 9769 10613 9778 10669
rect 7578 10589 9778 10613
rect 7578 10533 7587 10589
rect 7643 10533 7669 10589
rect 7725 10533 7751 10589
rect 7807 10533 7833 10589
rect 7889 10533 7915 10589
rect 7971 10533 7997 10589
rect 8053 10533 8079 10589
rect 8135 10533 8161 10589
rect 8217 10533 8243 10589
rect 8299 10533 8325 10589
rect 8381 10533 8407 10589
rect 8463 10533 8489 10589
rect 8545 10533 8571 10589
rect 8627 10533 8653 10589
rect 8709 10533 8735 10589
rect 8791 10533 8817 10589
rect 8873 10533 8899 10589
rect 8955 10533 8981 10589
rect 9037 10533 9063 10589
rect 9119 10533 9145 10589
rect 9201 10533 9227 10589
rect 9283 10533 9308 10589
rect 9364 10533 9389 10589
rect 9445 10533 9470 10589
rect 9526 10533 9551 10589
rect 9607 10533 9632 10589
rect 9688 10533 9713 10589
rect 9769 10533 9778 10589
rect 7578 10509 9778 10533
rect 7578 10453 7587 10509
rect 7643 10453 7669 10509
rect 7725 10453 7751 10509
rect 7807 10453 7833 10509
rect 7889 10453 7915 10509
rect 7971 10453 7997 10509
rect 8053 10453 8079 10509
rect 8135 10453 8161 10509
rect 8217 10453 8243 10509
rect 8299 10453 8325 10509
rect 8381 10453 8407 10509
rect 8463 10453 8489 10509
rect 8545 10453 8571 10509
rect 8627 10453 8653 10509
rect 8709 10453 8735 10509
rect 8791 10453 8817 10509
rect 8873 10453 8899 10509
rect 8955 10453 8981 10509
rect 9037 10453 9063 10509
rect 9119 10453 9145 10509
rect 9201 10453 9227 10509
rect 9283 10453 9308 10509
rect 9364 10453 9389 10509
rect 9445 10453 9470 10509
rect 9526 10453 9551 10509
rect 9607 10453 9632 10509
rect 9688 10453 9713 10509
rect 9769 10453 9778 10509
rect 7578 10429 9778 10453
rect 7578 10373 7587 10429
rect 7643 10373 7669 10429
rect 7725 10373 7751 10429
rect 7807 10373 7833 10429
rect 7889 10373 7915 10429
rect 7971 10373 7997 10429
rect 8053 10373 8079 10429
rect 8135 10373 8161 10429
rect 8217 10373 8243 10429
rect 8299 10373 8325 10429
rect 8381 10373 8407 10429
rect 8463 10373 8489 10429
rect 8545 10373 8571 10429
rect 8627 10373 8653 10429
rect 8709 10373 8735 10429
rect 8791 10373 8817 10429
rect 8873 10373 8899 10429
rect 8955 10373 8981 10429
rect 9037 10373 9063 10429
rect 9119 10373 9145 10429
rect 9201 10373 9227 10429
rect 9283 10373 9308 10429
rect 9364 10373 9389 10429
rect 9445 10373 9470 10429
rect 9526 10373 9551 10429
rect 9607 10373 9632 10429
rect 9688 10373 9713 10429
rect 9769 10373 9778 10429
rect 7578 10349 9778 10373
rect 7578 10293 7587 10349
rect 7643 10293 7669 10349
rect 7725 10293 7751 10349
rect 7807 10293 7833 10349
rect 7889 10293 7915 10349
rect 7971 10293 7997 10349
rect 8053 10293 8079 10349
rect 8135 10293 8161 10349
rect 8217 10293 8243 10349
rect 8299 10293 8325 10349
rect 8381 10293 8407 10349
rect 8463 10293 8489 10349
rect 8545 10293 8571 10349
rect 8627 10293 8653 10349
rect 8709 10293 8735 10349
rect 8791 10293 8817 10349
rect 8873 10293 8899 10349
rect 8955 10293 8981 10349
rect 9037 10293 9063 10349
rect 9119 10293 9145 10349
rect 9201 10293 9227 10349
rect 9283 10293 9308 10349
rect 9364 10293 9389 10349
rect 9445 10293 9470 10349
rect 9526 10293 9551 10349
rect 9607 10293 9632 10349
rect 9688 10293 9713 10349
rect 9769 10293 9778 10349
rect 7578 10269 9778 10293
rect 7578 10213 7587 10269
rect 7643 10213 7669 10269
rect 7725 10213 7751 10269
rect 7807 10213 7833 10269
rect 7889 10213 7915 10269
rect 7971 10213 7997 10269
rect 8053 10213 8079 10269
rect 8135 10213 8161 10269
rect 8217 10213 8243 10269
rect 8299 10213 8325 10269
rect 8381 10213 8407 10269
rect 8463 10213 8489 10269
rect 8545 10213 8571 10269
rect 8627 10213 8653 10269
rect 8709 10213 8735 10269
rect 8791 10213 8817 10269
rect 8873 10213 8899 10269
rect 8955 10213 8981 10269
rect 9037 10213 9063 10269
rect 9119 10213 9145 10269
rect 9201 10213 9227 10269
rect 9283 10213 9308 10269
rect 9364 10213 9389 10269
rect 9445 10213 9470 10269
rect 9526 10213 9551 10269
rect 9607 10213 9632 10269
rect 9688 10213 9713 10269
rect 9769 10213 9778 10269
rect 7578 10189 9778 10213
rect 7578 10133 7587 10189
rect 7643 10133 7669 10189
rect 7725 10133 7751 10189
rect 7807 10133 7833 10189
rect 7889 10133 7915 10189
rect 7971 10133 7997 10189
rect 8053 10133 8079 10189
rect 8135 10133 8161 10189
rect 8217 10133 8243 10189
rect 8299 10133 8325 10189
rect 8381 10133 8407 10189
rect 8463 10133 8489 10189
rect 8545 10133 8571 10189
rect 8627 10133 8653 10189
rect 8709 10133 8735 10189
rect 8791 10133 8817 10189
rect 8873 10133 8899 10189
rect 8955 10133 8981 10189
rect 9037 10133 9063 10189
rect 9119 10133 9145 10189
rect 9201 10133 9227 10189
rect 9283 10133 9308 10189
rect 9364 10133 9389 10189
rect 9445 10133 9470 10189
rect 9526 10133 9551 10189
rect 9607 10133 9632 10189
rect 9688 10133 9713 10189
rect 9769 10133 9778 10189
rect 7578 10109 9778 10133
rect 7578 10053 7587 10109
rect 7643 10053 7669 10109
rect 7725 10053 7751 10109
rect 7807 10053 7833 10109
rect 7889 10053 7915 10109
rect 7971 10053 7997 10109
rect 8053 10053 8079 10109
rect 8135 10053 8161 10109
rect 8217 10053 8243 10109
rect 8299 10053 8325 10109
rect 8381 10053 8407 10109
rect 8463 10053 8489 10109
rect 8545 10053 8571 10109
rect 8627 10053 8653 10109
rect 8709 10053 8735 10109
rect 8791 10053 8817 10109
rect 8873 10053 8899 10109
rect 8955 10053 8981 10109
rect 9037 10053 9063 10109
rect 9119 10053 9145 10109
rect 9201 10053 9227 10109
rect 9283 10053 9308 10109
rect 9364 10053 9389 10109
rect 9445 10053 9470 10109
rect 9526 10053 9551 10109
rect 9607 10053 9632 10109
rect 9688 10053 9713 10109
rect 9769 10053 9778 10109
rect 7578 10029 9778 10053
rect 7578 9973 7587 10029
rect 7643 9973 7669 10029
rect 7725 9973 7751 10029
rect 7807 9973 7833 10029
rect 7889 9973 7915 10029
rect 7971 9973 7997 10029
rect 8053 9973 8079 10029
rect 8135 9973 8161 10029
rect 8217 9973 8243 10029
rect 8299 9973 8325 10029
rect 8381 9973 8407 10029
rect 8463 9973 8489 10029
rect 8545 9973 8571 10029
rect 8627 9973 8653 10029
rect 8709 9973 8735 10029
rect 8791 9973 8817 10029
rect 8873 9973 8899 10029
rect 8955 9973 8981 10029
rect 9037 9973 9063 10029
rect 9119 9973 9145 10029
rect 9201 9973 9227 10029
rect 9283 9973 9308 10029
rect 9364 9973 9389 10029
rect 9445 9973 9470 10029
rect 9526 9973 9551 10029
rect 9607 9973 9632 10029
rect 9688 9973 9713 10029
rect 9769 9973 9778 10029
rect 7578 9949 9778 9973
rect 7578 9893 7587 9949
rect 7643 9893 7669 9949
rect 7725 9893 7751 9949
rect 7807 9893 7833 9949
rect 7889 9893 7915 9949
rect 7971 9893 7997 9949
rect 8053 9893 8079 9949
rect 8135 9893 8161 9949
rect 8217 9893 8243 9949
rect 8299 9893 8325 9949
rect 8381 9893 8407 9949
rect 8463 9893 8489 9949
rect 8545 9893 8571 9949
rect 8627 9893 8653 9949
rect 8709 9893 8735 9949
rect 8791 9893 8817 9949
rect 8873 9893 8899 9949
rect 8955 9893 8981 9949
rect 9037 9893 9063 9949
rect 9119 9893 9145 9949
rect 9201 9893 9227 9949
rect 9283 9893 9308 9949
rect 9364 9893 9389 9949
rect 9445 9893 9470 9949
rect 9526 9893 9551 9949
rect 9607 9893 9632 9949
rect 9688 9893 9713 9949
rect 9769 9893 9778 9949
rect 7578 9869 9778 9893
rect 7578 9813 7587 9869
rect 7643 9813 7669 9869
rect 7725 9813 7751 9869
rect 7807 9813 7833 9869
rect 7889 9813 7915 9869
rect 7971 9813 7997 9869
rect 8053 9813 8079 9869
rect 8135 9813 8161 9869
rect 8217 9813 8243 9869
rect 8299 9813 8325 9869
rect 8381 9813 8407 9869
rect 8463 9813 8489 9869
rect 8545 9813 8571 9869
rect 8627 9813 8653 9869
rect 8709 9813 8735 9869
rect 8791 9813 8817 9869
rect 8873 9813 8899 9869
rect 8955 9813 8981 9869
rect 9037 9813 9063 9869
rect 9119 9813 9145 9869
rect 9201 9813 9227 9869
rect 9283 9813 9308 9869
rect 9364 9813 9389 9869
rect 9445 9813 9470 9869
rect 9526 9813 9551 9869
rect 9607 9813 9632 9869
rect 9688 9813 9713 9869
rect 9769 9813 9778 9869
rect 7578 9789 9778 9813
rect 7578 9733 7587 9789
rect 7643 9733 7669 9789
rect 7725 9733 7751 9789
rect 7807 9733 7833 9789
rect 7889 9733 7915 9789
rect 7971 9733 7997 9789
rect 8053 9733 8079 9789
rect 8135 9733 8161 9789
rect 8217 9733 8243 9789
rect 8299 9733 8325 9789
rect 8381 9733 8407 9789
rect 8463 9733 8489 9789
rect 8545 9733 8571 9789
rect 8627 9733 8653 9789
rect 8709 9733 8735 9789
rect 8791 9733 8817 9789
rect 8873 9733 8899 9789
rect 8955 9733 8981 9789
rect 9037 9733 9063 9789
rect 9119 9733 9145 9789
rect 9201 9733 9227 9789
rect 9283 9733 9308 9789
rect 9364 9733 9389 9789
rect 9445 9733 9470 9789
rect 9526 9733 9551 9789
rect 9607 9733 9632 9789
rect 9688 9733 9713 9789
rect 9769 9733 9778 9789
rect 7578 9709 9778 9733
rect 7578 9653 7587 9709
rect 7643 9653 7669 9709
rect 7725 9653 7751 9709
rect 7807 9653 7833 9709
rect 7889 9653 7915 9709
rect 7971 9653 7997 9709
rect 8053 9653 8079 9709
rect 8135 9653 8161 9709
rect 8217 9653 8243 9709
rect 8299 9653 8325 9709
rect 8381 9653 8407 9709
rect 8463 9653 8489 9709
rect 8545 9653 8571 9709
rect 8627 9653 8653 9709
rect 8709 9653 8735 9709
rect 8791 9653 8817 9709
rect 8873 9653 8899 9709
rect 8955 9653 8981 9709
rect 9037 9653 9063 9709
rect 9119 9653 9145 9709
rect 9201 9653 9227 9709
rect 9283 9653 9308 9709
rect 9364 9653 9389 9709
rect 9445 9653 9470 9709
rect 9526 9653 9551 9709
rect 9607 9653 9632 9709
rect 9688 9653 9713 9709
rect 9769 9653 9778 9709
rect 7578 9629 9778 9653
rect 7578 9573 7587 9629
rect 7643 9573 7669 9629
rect 7725 9573 7751 9629
rect 7807 9573 7833 9629
rect 7889 9573 7915 9629
rect 7971 9573 7997 9629
rect 8053 9573 8079 9629
rect 8135 9573 8161 9629
rect 8217 9573 8243 9629
rect 8299 9573 8325 9629
rect 8381 9573 8407 9629
rect 8463 9573 8489 9629
rect 8545 9573 8571 9629
rect 8627 9573 8653 9629
rect 8709 9573 8735 9629
rect 8791 9573 8817 9629
rect 8873 9573 8899 9629
rect 8955 9573 8981 9629
rect 9037 9573 9063 9629
rect 9119 9573 9145 9629
rect 9201 9573 9227 9629
rect 9283 9573 9308 9629
rect 9364 9573 9389 9629
rect 9445 9573 9470 9629
rect 9526 9573 9551 9629
rect 9607 9573 9632 9629
rect 9688 9573 9713 9629
rect 9769 9573 9778 9629
rect 7578 9549 9778 9573
rect 7578 9493 7587 9549
rect 7643 9493 7669 9549
rect 7725 9493 7751 9549
rect 7807 9493 7833 9549
rect 7889 9493 7915 9549
rect 7971 9493 7997 9549
rect 8053 9493 8079 9549
rect 8135 9493 8161 9549
rect 8217 9493 8243 9549
rect 8299 9493 8325 9549
rect 8381 9493 8407 9549
rect 8463 9493 8489 9549
rect 8545 9493 8571 9549
rect 8627 9493 8653 9549
rect 8709 9493 8735 9549
rect 8791 9493 8817 9549
rect 8873 9493 8899 9549
rect 8955 9493 8981 9549
rect 9037 9493 9063 9549
rect 9119 9493 9145 9549
rect 9201 9493 9227 9549
rect 9283 9493 9308 9549
rect 9364 9493 9389 9549
rect 9445 9493 9470 9549
rect 9526 9493 9551 9549
rect 9607 9493 9632 9549
rect 9688 9493 9713 9549
rect 9769 9493 9778 9549
rect 7578 7296 9778 9493
rect 7578 7240 7588 7296
rect 7644 7240 7670 7296
rect 7726 7240 7751 7296
rect 7807 7240 7832 7296
rect 7888 7240 7913 7296
rect 7969 7240 7994 7296
rect 8050 7240 8075 7296
rect 8131 7240 8156 7296
rect 8212 7240 8237 7296
rect 8293 7240 8318 7296
rect 8374 7240 8399 7296
rect 8455 7240 8480 7296
rect 8536 7240 8561 7296
rect 8617 7240 8642 7296
rect 8698 7240 8723 7296
rect 8779 7240 8804 7296
rect 8860 7240 8885 7296
rect 8941 7240 8966 7296
rect 9022 7240 9047 7296
rect 9103 7240 9778 7296
rect 7578 7214 9778 7240
rect 7578 7158 7588 7214
rect 7644 7158 7670 7214
rect 7726 7158 7751 7214
rect 7807 7158 7832 7214
rect 7888 7158 7913 7214
rect 7969 7158 7994 7214
rect 8050 7158 8075 7214
rect 8131 7158 8156 7214
rect 8212 7158 8237 7214
rect 8293 7158 8318 7214
rect 8374 7158 8399 7214
rect 8455 7158 8480 7214
rect 8536 7158 8561 7214
rect 8617 7158 8642 7214
rect 8698 7158 8723 7214
rect 8779 7158 8804 7214
rect 8860 7158 8885 7214
rect 8941 7158 8966 7214
rect 9022 7158 9047 7214
rect 9103 7158 9778 7214
rect 7578 7132 9778 7158
rect 7578 7076 7588 7132
rect 7644 7076 7670 7132
rect 7726 7076 7751 7132
rect 7807 7076 7832 7132
rect 7888 7076 7913 7132
rect 7969 7076 7994 7132
rect 8050 7076 8075 7132
rect 8131 7076 8156 7132
rect 8212 7076 8237 7132
rect 8293 7076 8318 7132
rect 8374 7076 8399 7132
rect 8455 7076 8480 7132
rect 8536 7076 8561 7132
rect 8617 7076 8642 7132
rect 8698 7076 8723 7132
rect 8779 7076 8804 7132
rect 8860 7076 8885 7132
rect 8941 7076 8966 7132
rect 9022 7076 9047 7132
rect 9103 7076 9778 7132
rect 7578 7050 9778 7076
rect 7578 6994 7588 7050
rect 7644 6994 7670 7050
rect 7726 6994 7751 7050
rect 7807 6994 7832 7050
rect 7888 6994 7913 7050
rect 7969 6994 7994 7050
rect 8050 6994 8075 7050
rect 8131 6994 8156 7050
rect 8212 6994 8237 7050
rect 8293 6994 8318 7050
rect 8374 6994 8399 7050
rect 8455 6994 8480 7050
rect 8536 6994 8561 7050
rect 8617 6994 8642 7050
rect 8698 6994 8723 7050
rect 8779 6994 8804 7050
rect 8860 6994 8885 7050
rect 8941 6994 8966 7050
rect 9022 6994 9047 7050
rect 9103 6994 9778 7050
rect 7578 6968 9778 6994
rect 7578 6912 7588 6968
rect 7644 6912 7670 6968
rect 7726 6912 7751 6968
rect 7807 6912 7832 6968
rect 7888 6912 7913 6968
rect 7969 6912 7994 6968
rect 8050 6912 8075 6968
rect 8131 6912 8156 6968
rect 8212 6912 8237 6968
rect 8293 6912 8318 6968
rect 8374 6912 8399 6968
rect 8455 6912 8480 6968
rect 8536 6912 8561 6968
rect 8617 6912 8642 6968
rect 8698 6912 8723 6968
rect 8779 6912 8804 6968
rect 8860 6912 8885 6968
rect 8941 6912 8966 6968
rect 9022 6912 9047 6968
rect 9103 6912 9778 6968
rect 7578 6886 9778 6912
rect 7578 6830 7588 6886
rect 7644 6830 7670 6886
rect 7726 6830 7751 6886
rect 7807 6830 7832 6886
rect 7888 6830 7913 6886
rect 7969 6830 7994 6886
rect 8050 6830 8075 6886
rect 8131 6830 8156 6886
rect 8212 6830 8237 6886
rect 8293 6830 8318 6886
rect 8374 6830 8399 6886
rect 8455 6830 8480 6886
rect 8536 6830 8561 6886
rect 8617 6830 8642 6886
rect 8698 6830 8723 6886
rect 8779 6830 8804 6886
rect 8860 6830 8885 6886
rect 8941 6830 8966 6886
rect 9022 6830 9047 6886
rect 9103 6830 9778 6886
rect 7578 6804 9778 6830
rect 7578 6748 7588 6804
rect 7644 6748 7670 6804
rect 7726 6748 7751 6804
rect 7807 6748 7832 6804
rect 7888 6748 7913 6804
rect 7969 6748 7994 6804
rect 8050 6748 8075 6804
rect 8131 6748 8156 6804
rect 8212 6748 8237 6804
rect 8293 6748 8318 6804
rect 8374 6748 8399 6804
rect 8455 6748 8480 6804
rect 8536 6748 8561 6804
rect 8617 6748 8642 6804
rect 8698 6748 8723 6804
rect 8779 6748 8804 6804
rect 8860 6748 8885 6804
rect 8941 6748 8966 6804
rect 9022 6748 9047 6804
rect 9103 6748 9778 6804
rect 7578 6722 9778 6748
rect 7578 6666 7588 6722
rect 7644 6666 7670 6722
rect 7726 6666 7751 6722
rect 7807 6666 7832 6722
rect 7888 6666 7913 6722
rect 7969 6666 7994 6722
rect 8050 6666 8075 6722
rect 8131 6666 8156 6722
rect 8212 6666 8237 6722
rect 8293 6666 8318 6722
rect 8374 6666 8399 6722
rect 8455 6666 8480 6722
rect 8536 6666 8561 6722
rect 8617 6666 8642 6722
rect 8698 6666 8723 6722
rect 8779 6666 8804 6722
rect 8860 6666 8885 6722
rect 8941 6666 8966 6722
rect 9022 6666 9047 6722
rect 9103 6666 9778 6722
rect 7578 5092 9778 6666
rect 7578 5036 7587 5092
rect 7643 5036 7669 5092
rect 7725 5036 7751 5092
rect 7807 5036 7833 5092
rect 7889 5036 7915 5092
rect 7971 5036 7997 5092
rect 8053 5036 8079 5092
rect 8135 5036 8161 5092
rect 8217 5036 8243 5092
rect 8299 5036 8325 5092
rect 8381 5036 8407 5092
rect 8463 5036 8489 5092
rect 8545 5036 8571 5092
rect 8627 5036 8653 5092
rect 8709 5036 8735 5092
rect 8791 5036 8817 5092
rect 8873 5036 8899 5092
rect 8955 5036 8981 5092
rect 9037 5036 9063 5092
rect 9119 5036 9145 5092
rect 9201 5036 9227 5092
rect 9283 5036 9308 5092
rect 9364 5036 9389 5092
rect 9445 5036 9470 5092
rect 9526 5036 9551 5092
rect 9607 5036 9632 5092
rect 9688 5036 9713 5092
rect 9769 5036 9778 5092
rect 7578 5012 9778 5036
rect 7578 4956 7587 5012
rect 7643 4956 7669 5012
rect 7725 4956 7751 5012
rect 7807 4956 7833 5012
rect 7889 4956 7915 5012
rect 7971 4956 7997 5012
rect 8053 4956 8079 5012
rect 8135 4956 8161 5012
rect 8217 4956 8243 5012
rect 8299 4956 8325 5012
rect 8381 4956 8407 5012
rect 8463 4956 8489 5012
rect 8545 4956 8571 5012
rect 8627 4956 8653 5012
rect 8709 4956 8735 5012
rect 8791 4956 8817 5012
rect 8873 4956 8899 5012
rect 8955 4956 8981 5012
rect 9037 4956 9063 5012
rect 9119 4956 9145 5012
rect 9201 4956 9227 5012
rect 9283 4956 9308 5012
rect 9364 4956 9389 5012
rect 9445 4956 9470 5012
rect 9526 4956 9551 5012
rect 9607 4956 9632 5012
rect 9688 4956 9713 5012
rect 9769 4956 9778 5012
rect 7578 4932 9778 4956
rect 7578 4876 7587 4932
rect 7643 4876 7669 4932
rect 7725 4876 7751 4932
rect 7807 4876 7833 4932
rect 7889 4876 7915 4932
rect 7971 4876 7997 4932
rect 8053 4876 8079 4932
rect 8135 4876 8161 4932
rect 8217 4876 8243 4932
rect 8299 4876 8325 4932
rect 8381 4876 8407 4932
rect 8463 4876 8489 4932
rect 8545 4876 8571 4932
rect 8627 4876 8653 4932
rect 8709 4876 8735 4932
rect 8791 4876 8817 4932
rect 8873 4876 8899 4932
rect 8955 4876 8981 4932
rect 9037 4876 9063 4932
rect 9119 4876 9145 4932
rect 9201 4876 9227 4932
rect 9283 4876 9308 4932
rect 9364 4876 9389 4932
rect 9445 4876 9470 4932
rect 9526 4876 9551 4932
rect 9607 4876 9632 4932
rect 9688 4876 9713 4932
rect 9769 4876 9778 4932
rect 7578 4852 9778 4876
rect 7578 4796 7587 4852
rect 7643 4796 7669 4852
rect 7725 4796 7751 4852
rect 7807 4796 7833 4852
rect 7889 4796 7915 4852
rect 7971 4796 7997 4852
rect 8053 4796 8079 4852
rect 8135 4796 8161 4852
rect 8217 4796 8243 4852
rect 8299 4796 8325 4852
rect 8381 4796 8407 4852
rect 8463 4796 8489 4852
rect 8545 4796 8571 4852
rect 8627 4796 8653 4852
rect 8709 4796 8735 4852
rect 8791 4796 8817 4852
rect 8873 4796 8899 4852
rect 8955 4796 8981 4852
rect 9037 4796 9063 4852
rect 9119 4796 9145 4852
rect 9201 4796 9227 4852
rect 9283 4796 9308 4852
rect 9364 4796 9389 4852
rect 9445 4796 9470 4852
rect 9526 4796 9551 4852
rect 9607 4796 9632 4852
rect 9688 4796 9713 4852
rect 9769 4796 9778 4852
rect 7578 4772 9778 4796
rect 7578 4716 7587 4772
rect 7643 4716 7669 4772
rect 7725 4716 7751 4772
rect 7807 4716 7833 4772
rect 7889 4716 7915 4772
rect 7971 4716 7997 4772
rect 8053 4716 8079 4772
rect 8135 4716 8161 4772
rect 8217 4716 8243 4772
rect 8299 4716 8325 4772
rect 8381 4716 8407 4772
rect 8463 4716 8489 4772
rect 8545 4716 8571 4772
rect 8627 4716 8653 4772
rect 8709 4716 8735 4772
rect 8791 4716 8817 4772
rect 8873 4716 8899 4772
rect 8955 4716 8981 4772
rect 9037 4716 9063 4772
rect 9119 4716 9145 4772
rect 9201 4716 9227 4772
rect 9283 4716 9308 4772
rect 9364 4716 9389 4772
rect 9445 4716 9470 4772
rect 9526 4716 9551 4772
rect 9607 4716 9632 4772
rect 9688 4716 9713 4772
rect 9769 4716 9778 4772
rect 7578 4692 9778 4716
rect 7578 4636 7587 4692
rect 7643 4636 7669 4692
rect 7725 4636 7751 4692
rect 7807 4636 7833 4692
rect 7889 4636 7915 4692
rect 7971 4636 7997 4692
rect 8053 4636 8079 4692
rect 8135 4636 8161 4692
rect 8217 4636 8243 4692
rect 8299 4636 8325 4692
rect 8381 4636 8407 4692
rect 8463 4636 8489 4692
rect 8545 4636 8571 4692
rect 8627 4636 8653 4692
rect 8709 4636 8735 4692
rect 8791 4636 8817 4692
rect 8873 4636 8899 4692
rect 8955 4636 8981 4692
rect 9037 4636 9063 4692
rect 9119 4636 9145 4692
rect 9201 4636 9227 4692
rect 9283 4636 9308 4692
rect 9364 4636 9389 4692
rect 9445 4636 9470 4692
rect 9526 4636 9551 4692
rect 9607 4636 9632 4692
rect 9688 4636 9713 4692
rect 9769 4636 9778 4692
rect 7578 4612 9778 4636
rect 7578 4556 7587 4612
rect 7643 4556 7669 4612
rect 7725 4556 7751 4612
rect 7807 4556 7833 4612
rect 7889 4556 7915 4612
rect 7971 4556 7997 4612
rect 8053 4556 8079 4612
rect 8135 4556 8161 4612
rect 8217 4556 8243 4612
rect 8299 4556 8325 4612
rect 8381 4556 8407 4612
rect 8463 4556 8489 4612
rect 8545 4556 8571 4612
rect 8627 4556 8653 4612
rect 8709 4556 8735 4612
rect 8791 4556 8817 4612
rect 8873 4556 8899 4612
rect 8955 4556 8981 4612
rect 9037 4556 9063 4612
rect 9119 4556 9145 4612
rect 9201 4556 9227 4612
rect 9283 4556 9308 4612
rect 9364 4556 9389 4612
rect 9445 4556 9470 4612
rect 9526 4556 9551 4612
rect 9607 4556 9632 4612
rect 9688 4556 9713 4612
rect 9769 4556 9778 4612
rect 7578 4532 9778 4556
rect 7578 4476 7587 4532
rect 7643 4476 7669 4532
rect 7725 4476 7751 4532
rect 7807 4476 7833 4532
rect 7889 4476 7915 4532
rect 7971 4476 7997 4532
rect 8053 4476 8079 4532
rect 8135 4476 8161 4532
rect 8217 4476 8243 4532
rect 8299 4476 8325 4532
rect 8381 4476 8407 4532
rect 8463 4476 8489 4532
rect 8545 4476 8571 4532
rect 8627 4476 8653 4532
rect 8709 4476 8735 4532
rect 8791 4476 8817 4532
rect 8873 4476 8899 4532
rect 8955 4476 8981 4532
rect 9037 4476 9063 4532
rect 9119 4476 9145 4532
rect 9201 4476 9227 4532
rect 9283 4476 9308 4532
rect 9364 4476 9389 4532
rect 9445 4476 9470 4532
rect 9526 4476 9551 4532
rect 9607 4476 9632 4532
rect 9688 4476 9713 4532
rect 9769 4476 9778 4532
rect 7578 4452 9778 4476
rect 7578 4396 7587 4452
rect 7643 4396 7669 4452
rect 7725 4396 7751 4452
rect 7807 4396 7833 4452
rect 7889 4396 7915 4452
rect 7971 4396 7997 4452
rect 8053 4396 8079 4452
rect 8135 4396 8161 4452
rect 8217 4396 8243 4452
rect 8299 4396 8325 4452
rect 8381 4396 8407 4452
rect 8463 4396 8489 4452
rect 8545 4396 8571 4452
rect 8627 4396 8653 4452
rect 8709 4396 8735 4452
rect 8791 4396 8817 4452
rect 8873 4396 8899 4452
rect 8955 4396 8981 4452
rect 9037 4396 9063 4452
rect 9119 4396 9145 4452
rect 9201 4396 9227 4452
rect 9283 4396 9308 4452
rect 9364 4396 9389 4452
rect 9445 4396 9470 4452
rect 9526 4396 9551 4452
rect 9607 4396 9632 4452
rect 9688 4396 9713 4452
rect 9769 4396 9778 4452
rect 7578 4372 9778 4396
rect 7578 4316 7587 4372
rect 7643 4316 7669 4372
rect 7725 4316 7751 4372
rect 7807 4316 7833 4372
rect 7889 4316 7915 4372
rect 7971 4316 7997 4372
rect 8053 4316 8079 4372
rect 8135 4316 8161 4372
rect 8217 4316 8243 4372
rect 8299 4316 8325 4372
rect 8381 4316 8407 4372
rect 8463 4316 8489 4372
rect 8545 4316 8571 4372
rect 8627 4316 8653 4372
rect 8709 4316 8735 4372
rect 8791 4316 8817 4372
rect 8873 4316 8899 4372
rect 8955 4316 8981 4372
rect 9037 4316 9063 4372
rect 9119 4316 9145 4372
rect 9201 4316 9227 4372
rect 9283 4316 9308 4372
rect 9364 4316 9389 4372
rect 9445 4316 9470 4372
rect 9526 4316 9551 4372
rect 9607 4316 9632 4372
rect 9688 4316 9713 4372
rect 9769 4316 9778 4372
rect 7578 4292 9778 4316
rect 7578 4236 7587 4292
rect 7643 4236 7669 4292
rect 7725 4236 7751 4292
rect 7807 4236 7833 4292
rect 7889 4236 7915 4292
rect 7971 4236 7997 4292
rect 8053 4236 8079 4292
rect 8135 4236 8161 4292
rect 8217 4236 8243 4292
rect 8299 4236 8325 4292
rect 8381 4236 8407 4292
rect 8463 4236 8489 4292
rect 8545 4236 8571 4292
rect 8627 4236 8653 4292
rect 8709 4236 8735 4292
rect 8791 4236 8817 4292
rect 8873 4236 8899 4292
rect 8955 4236 8981 4292
rect 9037 4236 9063 4292
rect 9119 4236 9145 4292
rect 9201 4236 9227 4292
rect 9283 4236 9308 4292
rect 9364 4236 9389 4292
rect 9445 4236 9470 4292
rect 9526 4236 9551 4292
rect 9607 4236 9632 4292
rect 9688 4236 9713 4292
rect 9769 4236 9778 4292
rect 7578 4212 9778 4236
rect 7578 4156 7587 4212
rect 7643 4156 7669 4212
rect 7725 4156 7751 4212
rect 7807 4156 7833 4212
rect 7889 4156 7915 4212
rect 7971 4156 7997 4212
rect 8053 4156 8079 4212
rect 8135 4156 8161 4212
rect 8217 4156 8243 4212
rect 8299 4156 8325 4212
rect 8381 4156 8407 4212
rect 8463 4156 8489 4212
rect 8545 4156 8571 4212
rect 8627 4156 8653 4212
rect 8709 4156 8735 4212
rect 8791 4156 8817 4212
rect 8873 4156 8899 4212
rect 8955 4156 8981 4212
rect 9037 4156 9063 4212
rect 9119 4156 9145 4212
rect 9201 4156 9227 4212
rect 9283 4156 9308 4212
rect 9364 4156 9389 4212
rect 9445 4156 9470 4212
rect 9526 4156 9551 4212
rect 9607 4156 9632 4212
rect 9688 4156 9713 4212
rect 9769 4156 9778 4212
rect 7578 4132 9778 4156
rect 7578 4076 7587 4132
rect 7643 4076 7669 4132
rect 7725 4076 7751 4132
rect 7807 4076 7833 4132
rect 7889 4076 7915 4132
rect 7971 4076 7997 4132
rect 8053 4076 8079 4132
rect 8135 4076 8161 4132
rect 8217 4076 8243 4132
rect 8299 4076 8325 4132
rect 8381 4076 8407 4132
rect 8463 4076 8489 4132
rect 8545 4076 8571 4132
rect 8627 4076 8653 4132
rect 8709 4076 8735 4132
rect 8791 4076 8817 4132
rect 8873 4076 8899 4132
rect 8955 4076 8981 4132
rect 9037 4076 9063 4132
rect 9119 4076 9145 4132
rect 9201 4076 9227 4132
rect 9283 4076 9308 4132
rect 9364 4076 9389 4132
rect 9445 4076 9470 4132
rect 9526 4076 9551 4132
rect 9607 4076 9632 4132
rect 9688 4076 9713 4132
rect 9769 4076 9778 4132
rect 7578 4052 9778 4076
rect 7578 3996 7587 4052
rect 7643 3996 7669 4052
rect 7725 3996 7751 4052
rect 7807 3996 7833 4052
rect 7889 3996 7915 4052
rect 7971 3996 7997 4052
rect 8053 3996 8079 4052
rect 8135 3996 8161 4052
rect 8217 3996 8243 4052
rect 8299 3996 8325 4052
rect 8381 3996 8407 4052
rect 8463 3996 8489 4052
rect 8545 3996 8571 4052
rect 8627 3996 8653 4052
rect 8709 3996 8735 4052
rect 8791 3996 8817 4052
rect 8873 3996 8899 4052
rect 8955 3996 8981 4052
rect 9037 3996 9063 4052
rect 9119 3996 9145 4052
rect 9201 3996 9227 4052
rect 9283 3996 9308 4052
rect 9364 3996 9389 4052
rect 9445 3996 9470 4052
rect 9526 3996 9551 4052
rect 9607 3996 9632 4052
rect 9688 3996 9713 4052
rect 9769 3996 9778 4052
rect 7578 3972 9778 3996
rect 7578 3916 7587 3972
rect 7643 3916 7669 3972
rect 7725 3916 7751 3972
rect 7807 3916 7833 3972
rect 7889 3916 7915 3972
rect 7971 3916 7997 3972
rect 8053 3916 8079 3972
rect 8135 3916 8161 3972
rect 8217 3916 8243 3972
rect 8299 3916 8325 3972
rect 8381 3916 8407 3972
rect 8463 3916 8489 3972
rect 8545 3916 8571 3972
rect 8627 3916 8653 3972
rect 8709 3916 8735 3972
rect 8791 3916 8817 3972
rect 8873 3916 8899 3972
rect 8955 3916 8981 3972
rect 9037 3916 9063 3972
rect 9119 3916 9145 3972
rect 9201 3916 9227 3972
rect 9283 3916 9308 3972
rect 9364 3916 9389 3972
rect 9445 3916 9470 3972
rect 9526 3916 9551 3972
rect 9607 3916 9632 3972
rect 9688 3916 9713 3972
rect 9769 3916 9778 3972
rect 7578 3892 9778 3916
rect 7578 3836 7587 3892
rect 7643 3836 7669 3892
rect 7725 3836 7751 3892
rect 7807 3836 7833 3892
rect 7889 3836 7915 3892
rect 7971 3836 7997 3892
rect 8053 3836 8079 3892
rect 8135 3836 8161 3892
rect 8217 3836 8243 3892
rect 8299 3836 8325 3892
rect 8381 3836 8407 3892
rect 8463 3836 8489 3892
rect 8545 3836 8571 3892
rect 8627 3836 8653 3892
rect 8709 3836 8735 3892
rect 8791 3836 8817 3892
rect 8873 3836 8899 3892
rect 8955 3836 8981 3892
rect 9037 3836 9063 3892
rect 9119 3836 9145 3892
rect 9201 3836 9227 3892
rect 9283 3836 9308 3892
rect 9364 3836 9389 3892
rect 9445 3836 9470 3892
rect 9526 3836 9551 3892
rect 9607 3836 9632 3892
rect 9688 3836 9713 3892
rect 9769 3836 9778 3892
rect 7578 3812 9778 3836
rect 7578 3756 7587 3812
rect 7643 3756 7669 3812
rect 7725 3756 7751 3812
rect 7807 3756 7833 3812
rect 7889 3756 7915 3812
rect 7971 3756 7997 3812
rect 8053 3756 8079 3812
rect 8135 3756 8161 3812
rect 8217 3756 8243 3812
rect 8299 3756 8325 3812
rect 8381 3756 8407 3812
rect 8463 3756 8489 3812
rect 8545 3756 8571 3812
rect 8627 3756 8653 3812
rect 8709 3756 8735 3812
rect 8791 3756 8817 3812
rect 8873 3756 8899 3812
rect 8955 3756 8981 3812
rect 9037 3756 9063 3812
rect 9119 3756 9145 3812
rect 9201 3756 9227 3812
rect 9283 3756 9308 3812
rect 9364 3756 9389 3812
rect 9445 3756 9470 3812
rect 9526 3756 9551 3812
rect 9607 3756 9632 3812
rect 9688 3756 9713 3812
rect 9769 3756 9778 3812
rect 7578 3732 9778 3756
rect 7578 3676 7587 3732
rect 7643 3676 7669 3732
rect 7725 3676 7751 3732
rect 7807 3676 7833 3732
rect 7889 3676 7915 3732
rect 7971 3676 7997 3732
rect 8053 3676 8079 3732
rect 8135 3676 8161 3732
rect 8217 3676 8243 3732
rect 8299 3676 8325 3732
rect 8381 3676 8407 3732
rect 8463 3676 8489 3732
rect 8545 3676 8571 3732
rect 8627 3676 8653 3732
rect 8709 3676 8735 3732
rect 8791 3676 8817 3732
rect 8873 3676 8899 3732
rect 8955 3676 8981 3732
rect 9037 3676 9063 3732
rect 9119 3676 9145 3732
rect 9201 3676 9227 3732
rect 9283 3676 9308 3732
rect 9364 3676 9389 3732
rect 9445 3676 9470 3732
rect 9526 3676 9551 3732
rect 9607 3676 9632 3732
rect 9688 3676 9713 3732
rect 9769 3676 9778 3732
rect 7578 3652 9778 3676
rect 7578 3596 7587 3652
rect 7643 3596 7669 3652
rect 7725 3596 7751 3652
rect 7807 3596 7833 3652
rect 7889 3596 7915 3652
rect 7971 3596 7997 3652
rect 8053 3596 8079 3652
rect 8135 3596 8161 3652
rect 8217 3596 8243 3652
rect 8299 3596 8325 3652
rect 8381 3596 8407 3652
rect 8463 3596 8489 3652
rect 8545 3596 8571 3652
rect 8627 3596 8653 3652
rect 8709 3596 8735 3652
rect 8791 3596 8817 3652
rect 8873 3596 8899 3652
rect 8955 3596 8981 3652
rect 9037 3596 9063 3652
rect 9119 3596 9145 3652
rect 9201 3596 9227 3652
rect 9283 3596 9308 3652
rect 9364 3596 9389 3652
rect 9445 3596 9470 3652
rect 9526 3596 9551 3652
rect 9607 3596 9632 3652
rect 9688 3596 9713 3652
rect 9769 3596 9778 3652
rect 7578 3572 9778 3596
rect 7578 3516 7587 3572
rect 7643 3516 7669 3572
rect 7725 3516 7751 3572
rect 7807 3516 7833 3572
rect 7889 3516 7915 3572
rect 7971 3516 7997 3572
rect 8053 3516 8079 3572
rect 8135 3516 8161 3572
rect 8217 3516 8243 3572
rect 8299 3516 8325 3572
rect 8381 3516 8407 3572
rect 8463 3516 8489 3572
rect 8545 3516 8571 3572
rect 8627 3516 8653 3572
rect 8709 3516 8735 3572
rect 8791 3516 8817 3572
rect 8873 3516 8899 3572
rect 8955 3516 8981 3572
rect 9037 3516 9063 3572
rect 9119 3516 9145 3572
rect 9201 3516 9227 3572
rect 9283 3516 9308 3572
rect 9364 3516 9389 3572
rect 9445 3516 9470 3572
rect 9526 3516 9551 3572
rect 9607 3516 9632 3572
rect 9688 3516 9713 3572
rect 9769 3516 9778 3572
rect 7578 3492 9778 3516
rect 7578 3436 7587 3492
rect 7643 3436 7669 3492
rect 7725 3436 7751 3492
rect 7807 3436 7833 3492
rect 7889 3436 7915 3492
rect 7971 3436 7997 3492
rect 8053 3436 8079 3492
rect 8135 3436 8161 3492
rect 8217 3436 8243 3492
rect 8299 3436 8325 3492
rect 8381 3436 8407 3492
rect 8463 3436 8489 3492
rect 8545 3436 8571 3492
rect 8627 3436 8653 3492
rect 8709 3436 8735 3492
rect 8791 3436 8817 3492
rect 8873 3436 8899 3492
rect 8955 3436 8981 3492
rect 9037 3436 9063 3492
rect 9119 3436 9145 3492
rect 9201 3436 9227 3492
rect 9283 3436 9308 3492
rect 9364 3436 9389 3492
rect 9445 3436 9470 3492
rect 9526 3436 9551 3492
rect 9607 3436 9632 3492
rect 9688 3436 9713 3492
rect 9769 3436 9778 3492
rect 7578 3412 9778 3436
rect 7578 3356 7587 3412
rect 7643 3356 7669 3412
rect 7725 3356 7751 3412
rect 7807 3356 7833 3412
rect 7889 3356 7915 3412
rect 7971 3356 7997 3412
rect 8053 3356 8079 3412
rect 8135 3356 8161 3412
rect 8217 3356 8243 3412
rect 8299 3356 8325 3412
rect 8381 3356 8407 3412
rect 8463 3356 8489 3412
rect 8545 3356 8571 3412
rect 8627 3356 8653 3412
rect 8709 3356 8735 3412
rect 8791 3356 8817 3412
rect 8873 3356 8899 3412
rect 8955 3356 8981 3412
rect 9037 3356 9063 3412
rect 9119 3356 9145 3412
rect 9201 3356 9227 3412
rect 9283 3356 9308 3412
rect 9364 3356 9389 3412
rect 9445 3356 9470 3412
rect 9526 3356 9551 3412
rect 9607 3356 9632 3412
rect 9688 3356 9713 3412
rect 9769 3356 9778 3412
rect 7578 3332 9778 3356
rect 7578 3276 7587 3332
rect 7643 3276 7669 3332
rect 7725 3276 7751 3332
rect 7807 3276 7833 3332
rect 7889 3276 7915 3332
rect 7971 3276 7997 3332
rect 8053 3276 8079 3332
rect 8135 3276 8161 3332
rect 8217 3276 8243 3332
rect 8299 3276 8325 3332
rect 8381 3276 8407 3332
rect 8463 3276 8489 3332
rect 8545 3276 8571 3332
rect 8627 3276 8653 3332
rect 8709 3276 8735 3332
rect 8791 3276 8817 3332
rect 8873 3276 8899 3332
rect 8955 3276 8981 3332
rect 9037 3276 9063 3332
rect 9119 3276 9145 3332
rect 9201 3276 9227 3332
rect 9283 3276 9308 3332
rect 9364 3276 9389 3332
rect 9445 3276 9470 3332
rect 9526 3276 9551 3332
rect 9607 3276 9632 3332
rect 9688 3276 9713 3332
rect 9769 3276 9778 3332
rect 7578 3252 9778 3276
rect 7578 3196 7587 3252
rect 7643 3196 7669 3252
rect 7725 3196 7751 3252
rect 7807 3196 7833 3252
rect 7889 3196 7915 3252
rect 7971 3196 7997 3252
rect 8053 3196 8079 3252
rect 8135 3196 8161 3252
rect 8217 3196 8243 3252
rect 8299 3196 8325 3252
rect 8381 3196 8407 3252
rect 8463 3196 8489 3252
rect 8545 3196 8571 3252
rect 8627 3196 8653 3252
rect 8709 3196 8735 3252
rect 8791 3196 8817 3252
rect 8873 3196 8899 3252
rect 8955 3196 8981 3252
rect 9037 3196 9063 3252
rect 9119 3196 9145 3252
rect 9201 3196 9227 3252
rect 9283 3196 9308 3252
rect 9364 3196 9389 3252
rect 9445 3196 9470 3252
rect 9526 3196 9551 3252
rect 9607 3196 9632 3252
rect 9688 3196 9713 3252
rect 9769 3196 9778 3252
rect 7578 3172 9778 3196
rect 7578 3116 7587 3172
rect 7643 3116 7669 3172
rect 7725 3116 7751 3172
rect 7807 3116 7833 3172
rect 7889 3116 7915 3172
rect 7971 3116 7997 3172
rect 8053 3116 8079 3172
rect 8135 3116 8161 3172
rect 8217 3116 8243 3172
rect 8299 3116 8325 3172
rect 8381 3116 8407 3172
rect 8463 3116 8489 3172
rect 8545 3116 8571 3172
rect 8627 3116 8653 3172
rect 8709 3116 8735 3172
rect 8791 3116 8817 3172
rect 8873 3116 8899 3172
rect 8955 3116 8981 3172
rect 9037 3116 9063 3172
rect 9119 3116 9145 3172
rect 9201 3116 9227 3172
rect 9283 3116 9308 3172
rect 9364 3116 9389 3172
rect 9445 3116 9470 3172
rect 9526 3116 9551 3172
rect 9607 3116 9632 3172
rect 9688 3116 9713 3172
rect 9769 3116 9778 3172
rect 7578 3092 9778 3116
rect 7578 3036 7587 3092
rect 7643 3036 7669 3092
rect 7725 3036 7751 3092
rect 7807 3036 7833 3092
rect 7889 3036 7915 3092
rect 7971 3036 7997 3092
rect 8053 3036 8079 3092
rect 8135 3036 8161 3092
rect 8217 3036 8243 3092
rect 8299 3036 8325 3092
rect 8381 3036 8407 3092
rect 8463 3036 8489 3092
rect 8545 3036 8571 3092
rect 8627 3036 8653 3092
rect 8709 3036 8735 3092
rect 8791 3036 8817 3092
rect 8873 3036 8899 3092
rect 8955 3036 8981 3092
rect 9037 3036 9063 3092
rect 9119 3036 9145 3092
rect 9201 3036 9227 3092
rect 9283 3036 9308 3092
rect 9364 3036 9389 3092
rect 9445 3036 9470 3092
rect 9526 3036 9551 3092
rect 9607 3036 9632 3092
rect 9688 3036 9713 3092
rect 9769 3036 9778 3092
rect 7578 3012 9778 3036
rect 7578 2956 7587 3012
rect 7643 2956 7669 3012
rect 7725 2956 7751 3012
rect 7807 2956 7833 3012
rect 7889 2956 7915 3012
rect 7971 2956 7997 3012
rect 8053 2956 8079 3012
rect 8135 2956 8161 3012
rect 8217 2956 8243 3012
rect 8299 2956 8325 3012
rect 8381 2956 8407 3012
rect 8463 2956 8489 3012
rect 8545 2956 8571 3012
rect 8627 2956 8653 3012
rect 8709 2956 8735 3012
rect 8791 2956 8817 3012
rect 8873 2956 8899 3012
rect 8955 2956 8981 3012
rect 9037 2956 9063 3012
rect 9119 2956 9145 3012
rect 9201 2956 9227 3012
rect 9283 2956 9308 3012
rect 9364 2956 9389 3012
rect 9445 2956 9470 3012
rect 9526 2956 9551 3012
rect 9607 2956 9632 3012
rect 9688 2956 9713 3012
rect 9769 2956 9778 3012
rect 7578 2932 9778 2956
rect 7578 2876 7587 2932
rect 7643 2876 7669 2932
rect 7725 2876 7751 2932
rect 7807 2876 7833 2932
rect 7889 2876 7915 2932
rect 7971 2876 7997 2932
rect 8053 2876 8079 2932
rect 8135 2876 8161 2932
rect 8217 2876 8243 2932
rect 8299 2876 8325 2932
rect 8381 2876 8407 2932
rect 8463 2876 8489 2932
rect 8545 2876 8571 2932
rect 8627 2876 8653 2932
rect 8709 2876 8735 2932
rect 8791 2876 8817 2932
rect 8873 2876 8899 2932
rect 8955 2876 8981 2932
rect 9037 2876 9063 2932
rect 9119 2876 9145 2932
rect 9201 2876 9227 2932
rect 9283 2876 9308 2932
rect 9364 2876 9389 2932
rect 9445 2876 9470 2932
rect 9526 2876 9551 2932
rect 9607 2876 9632 2932
rect 9688 2876 9713 2932
rect 9769 2876 9778 2932
rect 7578 2852 9778 2876
rect 7578 2796 7587 2852
rect 7643 2796 7669 2852
rect 7725 2796 7751 2852
rect 7807 2796 7833 2852
rect 7889 2796 7915 2852
rect 7971 2796 7997 2852
rect 8053 2796 8079 2852
rect 8135 2796 8161 2852
rect 8217 2796 8243 2852
rect 8299 2796 8325 2852
rect 8381 2796 8407 2852
rect 8463 2796 8489 2852
rect 8545 2796 8571 2852
rect 8627 2796 8653 2852
rect 8709 2796 8735 2852
rect 8791 2796 8817 2852
rect 8873 2796 8899 2852
rect 8955 2796 8981 2852
rect 9037 2796 9063 2852
rect 9119 2796 9145 2852
rect 9201 2796 9227 2852
rect 9283 2796 9308 2852
rect 9364 2796 9389 2852
rect 9445 2796 9470 2852
rect 9526 2796 9551 2852
rect 9607 2796 9632 2852
rect 9688 2796 9713 2852
rect 9769 2796 9778 2852
rect 7578 2772 9778 2796
rect 7578 2716 7587 2772
rect 7643 2716 7669 2772
rect 7725 2716 7751 2772
rect 7807 2716 7833 2772
rect 7889 2716 7915 2772
rect 7971 2716 7997 2772
rect 8053 2716 8079 2772
rect 8135 2716 8161 2772
rect 8217 2716 8243 2772
rect 8299 2716 8325 2772
rect 8381 2716 8407 2772
rect 8463 2716 8489 2772
rect 8545 2716 8571 2772
rect 8627 2716 8653 2772
rect 8709 2716 8735 2772
rect 8791 2716 8817 2772
rect 8873 2716 8899 2772
rect 8955 2716 8981 2772
rect 9037 2716 9063 2772
rect 9119 2716 9145 2772
rect 9201 2716 9227 2772
rect 9283 2716 9308 2772
rect 9364 2716 9389 2772
rect 9445 2716 9470 2772
rect 9526 2716 9551 2772
rect 9607 2716 9632 2772
rect 9688 2716 9713 2772
rect 9769 2716 9778 2772
rect 7578 2692 9778 2716
rect 7578 2636 7587 2692
rect 7643 2636 7669 2692
rect 7725 2636 7751 2692
rect 7807 2636 7833 2692
rect 7889 2636 7915 2692
rect 7971 2636 7997 2692
rect 8053 2636 8079 2692
rect 8135 2636 8161 2692
rect 8217 2636 8243 2692
rect 8299 2636 8325 2692
rect 8381 2636 8407 2692
rect 8463 2636 8489 2692
rect 8545 2636 8571 2692
rect 8627 2636 8653 2692
rect 8709 2636 8735 2692
rect 8791 2636 8817 2692
rect 8873 2636 8899 2692
rect 8955 2636 8981 2692
rect 9037 2636 9063 2692
rect 9119 2636 9145 2692
rect 9201 2636 9227 2692
rect 9283 2636 9308 2692
rect 9364 2636 9389 2692
rect 9445 2636 9470 2692
rect 9526 2636 9551 2692
rect 9607 2636 9632 2692
rect 9688 2636 9713 2692
rect 9769 2636 9778 2692
rect 7578 2612 9778 2636
rect 7578 2556 7587 2612
rect 7643 2556 7669 2612
rect 7725 2556 7751 2612
rect 7807 2556 7833 2612
rect 7889 2556 7915 2612
rect 7971 2556 7997 2612
rect 8053 2556 8079 2612
rect 8135 2556 8161 2612
rect 8217 2556 8243 2612
rect 8299 2556 8325 2612
rect 8381 2556 8407 2612
rect 8463 2556 8489 2612
rect 8545 2556 8571 2612
rect 8627 2556 8653 2612
rect 8709 2556 8735 2612
rect 8791 2556 8817 2612
rect 8873 2556 8899 2612
rect 8955 2556 8981 2612
rect 9037 2556 9063 2612
rect 9119 2556 9145 2612
rect 9201 2556 9227 2612
rect 9283 2556 9308 2612
rect 9364 2556 9389 2612
rect 9445 2556 9470 2612
rect 9526 2556 9551 2612
rect 9607 2556 9632 2612
rect 9688 2556 9713 2612
rect 9769 2556 9778 2612
rect 7578 2532 9778 2556
rect 7578 2476 7587 2532
rect 7643 2476 7669 2532
rect 7725 2476 7751 2532
rect 7807 2476 7833 2532
rect 7889 2476 7915 2532
rect 7971 2476 7997 2532
rect 8053 2476 8079 2532
rect 8135 2476 8161 2532
rect 8217 2476 8243 2532
rect 8299 2476 8325 2532
rect 8381 2476 8407 2532
rect 8463 2476 8489 2532
rect 8545 2476 8571 2532
rect 8627 2476 8653 2532
rect 8709 2476 8735 2532
rect 8791 2476 8817 2532
rect 8873 2476 8899 2532
rect 8955 2476 8981 2532
rect 9037 2476 9063 2532
rect 9119 2476 9145 2532
rect 9201 2476 9227 2532
rect 9283 2476 9308 2532
rect 9364 2476 9389 2532
rect 9445 2476 9470 2532
rect 9526 2476 9551 2532
rect 9607 2476 9632 2532
rect 9688 2476 9713 2532
rect 9769 2476 9778 2532
rect 7578 0 9778 2476
<< comment >>
rect 2898 37036 13268 39036
rect 2898 34080 13268 36436
tri 1500 33090 2490 34080 se
rect 2490 33090 13268 34080
tri 13268 33090 13500 33322 sw
rect 1500 21070 13500 33090
tri 1500 20080 2490 21070 ne
rect 2490 20080 12510 21070
tri 12510 20080 13500 21070 nw
rect 2898 9436 13268 13436
use DFL1_CDNS_52468879185823  DFL1_CDNS_52468879185823_0
timestamp 1707688321
transform 1 0 12569 0 1 37069
box -26 -26 144 1920
use DFL1_CDNS_52468879185823  DFL1_CDNS_52468879185823_1
timestamp 1707688321
transform 1 0 11649 0 1 37069
box -26 -26 144 1920
use DFL1_CDNS_52468879185823  DFL1_CDNS_52468879185823_2
timestamp 1707688321
transform 1 0 10729 0 1 37069
box -26 -26 144 1920
use DFL1_CDNS_52468879185823  DFL1_CDNS_52468879185823_3
timestamp 1707688321
transform 1 0 9809 0 1 37069
box -26 -26 144 1920
use DFL1_CDNS_52468879185823  DFL1_CDNS_52468879185823_4
timestamp 1707688321
transform 1 0 8889 0 1 37069
box -26 -26 144 1920
use DFL1_CDNS_52468879185823  DFL1_CDNS_52468879185823_5
timestamp 1707688321
transform 1 0 7969 0 1 37069
box -26 -26 144 1920
use DFL1_CDNS_52468879185823  DFL1_CDNS_52468879185823_6
timestamp 1707688321
transform 1 0 7049 0 1 37069
box -26 -26 144 1920
use DFL1_CDNS_52468879185823  DFL1_CDNS_52468879185823_7
timestamp 1707688321
transform 1 0 6129 0 1 37069
box -26 -26 144 1920
use DFL1_CDNS_52468879185823  DFL1_CDNS_52468879185823_8
timestamp 1707688321
transform 1 0 5209 0 1 37069
box -26 -26 144 1920
use DFL1_CDNS_52468879185823  DFL1_CDNS_52468879185823_9
timestamp 1707688321
transform 1 0 4289 0 1 37069
box -26 -26 144 1920
use DFL1_CDNS_52468879185823  DFL1_CDNS_52468879185823_10
timestamp 1707688321
transform 1 0 3369 0 1 37069
box -26 -26 144 1920
use DFL1_CDNS_52468879185824  DFL1_CDNS_52468879185824_0
timestamp 1707688321
transform 1 0 6129 0 1 18669
box -26 -26 144 3960
use DFL1_CDNS_52468879185824  DFL1_CDNS_52468879185824_1
timestamp 1707688321
transform 1 0 12569 0 1 18669
box -26 -26 144 3960
use DFL1_CDNS_52468879185824  DFL1_CDNS_52468879185824_2
timestamp 1707688321
transform 1 0 11649 0 1 18669
box -26 -26 144 3960
use DFL1_CDNS_52468879185824  DFL1_CDNS_52468879185824_3
timestamp 1707688321
transform 1 0 10729 0 1 18669
box -26 -26 144 3960
use DFL1_CDNS_52468879185824  DFL1_CDNS_52468879185824_4
timestamp 1707688321
transform 1 0 9809 0 1 18669
box -26 -26 144 3960
use DFL1_CDNS_52468879185824  DFL1_CDNS_52468879185824_5
timestamp 1707688321
transform 1 0 8889 0 1 18669
box -26 -26 144 3960
use DFL1_CDNS_52468879185824  DFL1_CDNS_52468879185824_6
timestamp 1707688321
transform 1 0 7969 0 1 18669
box -26 -26 144 3960
use DFL1_CDNS_52468879185824  DFL1_CDNS_52468879185824_7
timestamp 1707688321
transform 1 0 7049 0 1 18669
box -26 -26 144 3960
use DFL1_CDNS_52468879185824  DFL1_CDNS_52468879185824_8
timestamp 1707688321
transform 1 0 5209 0 1 18669
box -26 -26 144 3960
use DFL1_CDNS_52468879185824  DFL1_CDNS_52468879185824_9
timestamp 1707688321
transform 1 0 3369 0 1 27869
box -26 -26 144 3960
use DFL1_CDNS_52468879185824  DFL1_CDNS_52468879185824_10
timestamp 1707688321
transform 1 0 5209 0 1 27869
box -26 -26 144 3960
use DFL1_CDNS_52468879185824  DFL1_CDNS_52468879185824_11
timestamp 1707688321
transform 1 0 6129 0 1 27869
box -26 -26 144 3960
use DFL1_CDNS_52468879185824  DFL1_CDNS_52468879185824_12
timestamp 1707688321
transform 1 0 7049 0 1 27869
box -26 -26 144 3960
use DFL1_CDNS_52468879185824  DFL1_CDNS_52468879185824_13
timestamp 1707688321
transform 1 0 7969 0 1 27869
box -26 -26 144 3960
use DFL1_CDNS_52468879185824  DFL1_CDNS_52468879185824_14
timestamp 1707688321
transform 1 0 8889 0 1 27869
box -26 -26 144 3960
use DFL1_CDNS_52468879185824  DFL1_CDNS_52468879185824_15
timestamp 1707688321
transform 1 0 9809 0 1 27869
box -26 -26 144 3960
use DFL1_CDNS_52468879185824  DFL1_CDNS_52468879185824_16
timestamp 1707688321
transform 1 0 10729 0 1 27869
box -26 -26 144 3960
use DFL1_CDNS_52468879185824  DFL1_CDNS_52468879185824_17
timestamp 1707688321
transform 1 0 11649 0 1 27869
box -26 -26 144 3960
use DFL1_CDNS_52468879185824  DFL1_CDNS_52468879185824_18
timestamp 1707688321
transform 1 0 12569 0 1 27869
box -26 -26 144 3960
use DFL1_CDNS_52468879185824  DFL1_CDNS_52468879185824_19
timestamp 1707688321
transform 1 0 4289 0 1 27869
box -26 -26 144 3960
use DFL1_CDNS_52468879185824  DFL1_CDNS_52468879185824_20
timestamp 1707688321
transform 1 0 3369 0 1 32469
box -26 -26 144 3960
use DFL1_CDNS_52468879185824  DFL1_CDNS_52468879185824_21
timestamp 1707688321
transform 1 0 5209 0 1 32469
box -26 -26 144 3960
use DFL1_CDNS_52468879185824  DFL1_CDNS_52468879185824_22
timestamp 1707688321
transform 1 0 6129 0 1 32469
box -26 -26 144 3960
use DFL1_CDNS_52468879185824  DFL1_CDNS_52468879185824_23
timestamp 1707688321
transform 1 0 7049 0 1 32469
box -26 -26 144 3960
use DFL1_CDNS_52468879185824  DFL1_CDNS_52468879185824_24
timestamp 1707688321
transform 1 0 7969 0 1 32469
box -26 -26 144 3960
use DFL1_CDNS_52468879185824  DFL1_CDNS_52468879185824_25
timestamp 1707688321
transform 1 0 8889 0 1 32469
box -26 -26 144 3960
use DFL1_CDNS_52468879185824  DFL1_CDNS_52468879185824_26
timestamp 1707688321
transform 1 0 9809 0 1 32469
box -26 -26 144 3960
use DFL1_CDNS_52468879185824  DFL1_CDNS_52468879185824_27
timestamp 1707688321
transform 1 0 10729 0 1 32469
box -26 -26 144 3960
use DFL1_CDNS_52468879185824  DFL1_CDNS_52468879185824_28
timestamp 1707688321
transform 1 0 11649 0 1 32469
box -26 -26 144 3960
use DFL1_CDNS_52468879185824  DFL1_CDNS_52468879185824_29
timestamp 1707688321
transform 1 0 12569 0 1 32469
box -26 -26 144 3960
use DFL1_CDNS_52468879185824  DFL1_CDNS_52468879185824_30
timestamp 1707688321
transform 1 0 4289 0 1 32469
box -26 -26 144 3960
use DFL1_CDNS_52468879185824  DFL1_CDNS_52468879185824_31
timestamp 1707688321
transform 1 0 6129 0 1 23269
box -26 -26 144 3960
use DFL1_CDNS_52468879185824  DFL1_CDNS_52468879185824_32
timestamp 1707688321
transform 1 0 12569 0 1 23269
box -26 -26 144 3960
use DFL1_CDNS_52468879185824  DFL1_CDNS_52468879185824_33
timestamp 1707688321
transform 1 0 11649 0 1 23269
box -26 -26 144 3960
use DFL1_CDNS_52468879185824  DFL1_CDNS_52468879185824_34
timestamp 1707688321
transform 1 0 10729 0 1 23269
box -26 -26 144 3960
use DFL1_CDNS_52468879185824  DFL1_CDNS_52468879185824_35
timestamp 1707688321
transform 1 0 9809 0 1 23269
box -26 -26 144 3960
use DFL1_CDNS_52468879185824  DFL1_CDNS_52468879185824_36
timestamp 1707688321
transform 1 0 8889 0 1 23269
box -26 -26 144 3960
use DFL1_CDNS_52468879185824  DFL1_CDNS_52468879185824_37
timestamp 1707688321
transform 1 0 7969 0 1 23269
box -26 -26 144 3960
use DFL1_CDNS_52468879185824  DFL1_CDNS_52468879185824_38
timestamp 1707688321
transform 1 0 7049 0 1 23269
box -26 -26 144 3960
use DFL1_CDNS_52468879185824  DFL1_CDNS_52468879185824_39
timestamp 1707688321
transform 1 0 5209 0 1 23269
box -26 -26 144 3960
use DFL1_CDNS_52468879185824  DFL1_CDNS_52468879185824_40
timestamp 1707688321
transform 1 0 5209 0 1 14069
box -26 -26 144 3960
use DFL1_CDNS_52468879185824  DFL1_CDNS_52468879185824_41
timestamp 1707688321
transform 1 0 7049 0 1 14069
box -26 -26 144 3960
use DFL1_CDNS_52468879185824  DFL1_CDNS_52468879185824_42
timestamp 1707688321
transform 1 0 7969 0 1 14069
box -26 -26 144 3960
use DFL1_CDNS_52468879185824  DFL1_CDNS_52468879185824_43
timestamp 1707688321
transform 1 0 8889 0 1 14069
box -26 -26 144 3960
use DFL1_CDNS_52468879185824  DFL1_CDNS_52468879185824_44
timestamp 1707688321
transform 1 0 9809 0 1 14069
box -26 -26 144 3960
use DFL1_CDNS_52468879185824  DFL1_CDNS_52468879185824_45
timestamp 1707688321
transform 1 0 10729 0 1 14069
box -26 -26 144 3960
use DFL1_CDNS_52468879185824  DFL1_CDNS_52468879185824_46
timestamp 1707688321
transform 1 0 11649 0 1 14069
box -26 -26 144 3960
use DFL1_CDNS_52468879185824  DFL1_CDNS_52468879185824_47
timestamp 1707688321
transform 1 0 12569 0 1 14069
box -26 -26 144 3960
use DFL1_CDNS_52468879185824  DFL1_CDNS_52468879185824_48
timestamp 1707688321
transform 1 0 6129 0 1 14069
box -26 -26 144 3960
use DFL1_CDNS_52468879185824  DFL1_CDNS_52468879185824_49
timestamp 1707688321
transform 1 0 4289 0 1 9469
box -26 -26 144 3960
use DFL1_CDNS_52468879185824  DFL1_CDNS_52468879185824_50
timestamp 1707688321
transform 1 0 12569 0 1 9469
box -26 -26 144 3960
use DFL1_CDNS_52468879185824  DFL1_CDNS_52468879185824_51
timestamp 1707688321
transform 1 0 11649 0 1 9469
box -26 -26 144 3960
use DFL1_CDNS_52468879185824  DFL1_CDNS_52468879185824_52
timestamp 1707688321
transform 1 0 10729 0 1 9469
box -26 -26 144 3960
use DFL1_CDNS_52468879185824  DFL1_CDNS_52468879185824_53
timestamp 1707688321
transform 1 0 9809 0 1 9469
box -26 -26 144 3960
use DFL1_CDNS_52468879185824  DFL1_CDNS_52468879185824_54
timestamp 1707688321
transform 1 0 8889 0 1 9469
box -26 -26 144 3960
use DFL1_CDNS_52468879185824  DFL1_CDNS_52468879185824_55
timestamp 1707688321
transform 1 0 7969 0 1 9469
box -26 -26 144 3960
use DFL1_CDNS_52468879185824  DFL1_CDNS_52468879185824_56
timestamp 1707688321
transform 1 0 7049 0 1 9469
box -26 -26 144 3960
use DFL1_CDNS_52468879185824  DFL1_CDNS_52468879185824_57
timestamp 1707688321
transform 1 0 6129 0 1 9469
box -26 -26 144 3960
use DFL1_CDNS_52468879185824  DFL1_CDNS_52468879185824_58
timestamp 1707688321
transform 1 0 5209 0 1 9469
box -26 -26 144 3960
use DFL1_CDNS_52468879185824  DFL1_CDNS_52468879185824_59
timestamp 1707688321
transform 1 0 3369 0 1 9469
box -26 -26 144 3960
use hvnTran_CDNS_52468879185825  hvnTran_CDNS_52468879185825_0
timestamp 1707688321
transform -1 0 12363 0 -1 5429
box -79 -26 879 1026
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_0
timestamp 1707688321
transform 1 0 4096 0 1 39074
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_1
timestamp 1707688321
transform 1 0 5016 0 1 39074
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_2
timestamp 1707688321
transform 1 0 5936 0 1 39074
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_3
timestamp 1707688321
transform 1 0 6856 0 1 39074
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_4
timestamp 1707688321
transform 1 0 7776 0 1 39074
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_5
timestamp 1707688321
transform 1 0 8696 0 1 39074
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_6
timestamp 1707688321
transform 1 0 9616 0 1 39074
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_7
timestamp 1707688321
transform 1 0 10536 0 1 39074
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_8
timestamp 1707688321
transform 1 0 11456 0 1 39074
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_9
timestamp 1707688321
transform 1 0 12376 0 1 39074
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_10
timestamp 1707688321
transform 1 0 3176 0 1 39074
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_11
timestamp 1707688321
transform 1 0 12778 0 1 39074
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_12
timestamp 1707688321
transform 1 0 11858 0 1 39074
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_13
timestamp 1707688321
transform 1 0 10938 0 1 39074
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_14
timestamp 1707688321
transform 1 0 10018 0 1 39074
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_15
timestamp 1707688321
transform 1 0 9098 0 1 39074
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_16
timestamp 1707688321
transform 1 0 8178 0 1 39074
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_17
timestamp 1707688321
transform 1 0 7258 0 1 39074
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_18
timestamp 1707688321
transform 1 0 6338 0 1 39074
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_19
timestamp 1707688321
transform 1 0 5418 0 1 39074
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_20
timestamp 1707688321
transform 1 0 4498 0 1 39074
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_21
timestamp 1707688321
transform 1 0 3578 0 1 39074
box 0 0 1 1
use L1M1_CDNS_52468879185821  L1M1_CDNS_52468879185821_0
timestamp 1707688321
transform 1 0 5213 0 1 18705
box -12 -6 118 3640
use L1M1_CDNS_52468879185821  L1M1_CDNS_52468879185821_1
timestamp 1707688321
transform 1 0 6133 0 1 18705
box -12 -6 118 3640
use L1M1_CDNS_52468879185821  L1M1_CDNS_52468879185821_2
timestamp 1707688321
transform 1 0 7053 0 1 18705
box -12 -6 118 3640
use L1M1_CDNS_52468879185821  L1M1_CDNS_52468879185821_3
timestamp 1707688321
transform 1 0 7973 0 1 18705
box -12 -6 118 3640
use L1M1_CDNS_52468879185821  L1M1_CDNS_52468879185821_4
timestamp 1707688321
transform 1 0 8893 0 1 18705
box -12 -6 118 3640
use L1M1_CDNS_52468879185821  L1M1_CDNS_52468879185821_5
timestamp 1707688321
transform 1 0 9813 0 1 18705
box -12 -6 118 3640
use L1M1_CDNS_52468879185821  L1M1_CDNS_52468879185821_6
timestamp 1707688321
transform 1 0 10733 0 1 18705
box -12 -6 118 3640
use L1M1_CDNS_52468879185821  L1M1_CDNS_52468879185821_7
timestamp 1707688321
transform 1 0 11653 0 1 18705
box -12 -6 118 3640
use L1M1_CDNS_52468879185821  L1M1_CDNS_52468879185821_8
timestamp 1707688321
transform 1 0 12573 0 1 18705
box -12 -6 118 3640
use L1M1_CDNS_52468879185821  L1M1_CDNS_52468879185821_9
timestamp 1707688321
transform 1 0 12573 0 1 27905
box -12 -6 118 3640
use L1M1_CDNS_52468879185821  L1M1_CDNS_52468879185821_10
timestamp 1707688321
transform 1 0 11653 0 1 27905
box -12 -6 118 3640
use L1M1_CDNS_52468879185821  L1M1_CDNS_52468879185821_11
timestamp 1707688321
transform 1 0 10733 0 1 27905
box -12 -6 118 3640
use L1M1_CDNS_52468879185821  L1M1_CDNS_52468879185821_12
timestamp 1707688321
transform 1 0 9813 0 1 27905
box -12 -6 118 3640
use L1M1_CDNS_52468879185821  L1M1_CDNS_52468879185821_13
timestamp 1707688321
transform 1 0 8893 0 1 27905
box -12 -6 118 3640
use L1M1_CDNS_52468879185821  L1M1_CDNS_52468879185821_14
timestamp 1707688321
transform 1 0 7973 0 1 27905
box -12 -6 118 3640
use L1M1_CDNS_52468879185821  L1M1_CDNS_52468879185821_15
timestamp 1707688321
transform 1 0 7053 0 1 27905
box -12 -6 118 3640
use L1M1_CDNS_52468879185821  L1M1_CDNS_52468879185821_16
timestamp 1707688321
transform 1 0 6133 0 1 27905
box -12 -6 118 3640
use L1M1_CDNS_52468879185821  L1M1_CDNS_52468879185821_17
timestamp 1707688321
transform 1 0 5213 0 1 27905
box -12 -6 118 3640
use L1M1_CDNS_52468879185821  L1M1_CDNS_52468879185821_18
timestamp 1707688321
transform 1 0 4293 0 1 27905
box -12 -6 118 3640
use L1M1_CDNS_52468879185821  L1M1_CDNS_52468879185821_19
timestamp 1707688321
transform 1 0 3373 0 1 27905
box -12 -6 118 3640
use L1M1_CDNS_52468879185821  L1M1_CDNS_52468879185821_20
timestamp 1707688321
transform 1 0 12573 0 1 32505
box -12 -6 118 3640
use L1M1_CDNS_52468879185821  L1M1_CDNS_52468879185821_21
timestamp 1707688321
transform 1 0 11653 0 1 32505
box -12 -6 118 3640
use L1M1_CDNS_52468879185821  L1M1_CDNS_52468879185821_22
timestamp 1707688321
transform 1 0 10733 0 1 32505
box -12 -6 118 3640
use L1M1_CDNS_52468879185821  L1M1_CDNS_52468879185821_23
timestamp 1707688321
transform 1 0 9813 0 1 32505
box -12 -6 118 3640
use L1M1_CDNS_52468879185821  L1M1_CDNS_52468879185821_24
timestamp 1707688321
transform 1 0 8893 0 1 32505
box -12 -6 118 3640
use L1M1_CDNS_52468879185821  L1M1_CDNS_52468879185821_25
timestamp 1707688321
transform 1 0 7973 0 1 32505
box -12 -6 118 3640
use L1M1_CDNS_52468879185821  L1M1_CDNS_52468879185821_26
timestamp 1707688321
transform 1 0 7053 0 1 32505
box -12 -6 118 3640
use L1M1_CDNS_52468879185821  L1M1_CDNS_52468879185821_27
timestamp 1707688321
transform 1 0 6133 0 1 32505
box -12 -6 118 3640
use L1M1_CDNS_52468879185821  L1M1_CDNS_52468879185821_28
timestamp 1707688321
transform 1 0 5213 0 1 32505
box -12 -6 118 3640
use L1M1_CDNS_52468879185821  L1M1_CDNS_52468879185821_29
timestamp 1707688321
transform 1 0 4293 0 1 32505
box -12 -6 118 3640
use L1M1_CDNS_52468879185821  L1M1_CDNS_52468879185821_30
timestamp 1707688321
transform 1 0 3373 0 1 32505
box -12 -6 118 3640
use L1M1_CDNS_52468879185821  L1M1_CDNS_52468879185821_31
timestamp 1707688321
transform 1 0 5213 0 1 23305
box -12 -6 118 3640
use L1M1_CDNS_52468879185821  L1M1_CDNS_52468879185821_32
timestamp 1707688321
transform 1 0 6133 0 1 23305
box -12 -6 118 3640
use L1M1_CDNS_52468879185821  L1M1_CDNS_52468879185821_33
timestamp 1707688321
transform 1 0 7053 0 1 23305
box -12 -6 118 3640
use L1M1_CDNS_52468879185821  L1M1_CDNS_52468879185821_34
timestamp 1707688321
transform 1 0 7973 0 1 23305
box -12 -6 118 3640
use L1M1_CDNS_52468879185821  L1M1_CDNS_52468879185821_35
timestamp 1707688321
transform 1 0 8893 0 1 23305
box -12 -6 118 3640
use L1M1_CDNS_52468879185821  L1M1_CDNS_52468879185821_36
timestamp 1707688321
transform 1 0 9813 0 1 23305
box -12 -6 118 3640
use L1M1_CDNS_52468879185821  L1M1_CDNS_52468879185821_37
timestamp 1707688321
transform 1 0 10733 0 1 23305
box -12 -6 118 3640
use L1M1_CDNS_52468879185821  L1M1_CDNS_52468879185821_38
timestamp 1707688321
transform 1 0 11653 0 1 23305
box -12 -6 118 3640
use L1M1_CDNS_52468879185821  L1M1_CDNS_52468879185821_39
timestamp 1707688321
transform 1 0 12573 0 1 23305
box -12 -6 118 3640
use L1M1_CDNS_52468879185821  L1M1_CDNS_52468879185821_40
timestamp 1707688321
transform 1 0 12573 0 1 14105
box -12 -6 118 3640
use L1M1_CDNS_52468879185821  L1M1_CDNS_52468879185821_41
timestamp 1707688321
transform 1 0 11653 0 1 14105
box -12 -6 118 3640
use L1M1_CDNS_52468879185821  L1M1_CDNS_52468879185821_42
timestamp 1707688321
transform 1 0 10733 0 1 14105
box -12 -6 118 3640
use L1M1_CDNS_52468879185821  L1M1_CDNS_52468879185821_43
timestamp 1707688321
transform 1 0 9813 0 1 14105
box -12 -6 118 3640
use L1M1_CDNS_52468879185821  L1M1_CDNS_52468879185821_44
timestamp 1707688321
transform 1 0 8893 0 1 14105
box -12 -6 118 3640
use L1M1_CDNS_52468879185821  L1M1_CDNS_52468879185821_45
timestamp 1707688321
transform 1 0 7973 0 1 14105
box -12 -6 118 3640
use L1M1_CDNS_52468879185821  L1M1_CDNS_52468879185821_46
timestamp 1707688321
transform 1 0 7053 0 1 14105
box -12 -6 118 3640
use L1M1_CDNS_52468879185821  L1M1_CDNS_52468879185821_47
timestamp 1707688321
transform 1 0 6133 0 1 14105
box -12 -6 118 3640
use L1M1_CDNS_52468879185821  L1M1_CDNS_52468879185821_48
timestamp 1707688321
transform 1 0 5213 0 1 14105
box -12 -6 118 3640
use L1M1_CDNS_52468879185821  L1M1_CDNS_52468879185821_49
timestamp 1707688321
transform 1 0 3373 0 1 9505
box -12 -6 118 3640
use L1M1_CDNS_52468879185821  L1M1_CDNS_52468879185821_50
timestamp 1707688321
transform 1 0 4293 0 1 9505
box -12 -6 118 3640
use L1M1_CDNS_52468879185821  L1M1_CDNS_52468879185821_51
timestamp 1707688321
transform 1 0 5213 0 1 9505
box -12 -6 118 3640
use L1M1_CDNS_52468879185821  L1M1_CDNS_52468879185821_52
timestamp 1707688321
transform 1 0 6133 0 1 9505
box -12 -6 118 3640
use L1M1_CDNS_52468879185821  L1M1_CDNS_52468879185821_53
timestamp 1707688321
transform 1 0 7053 0 1 9505
box -12 -6 118 3640
use L1M1_CDNS_52468879185821  L1M1_CDNS_52468879185821_54
timestamp 1707688321
transform 1 0 7973 0 1 9505
box -12 -6 118 3640
use L1M1_CDNS_52468879185821  L1M1_CDNS_52468879185821_55
timestamp 1707688321
transform 1 0 8893 0 1 9505
box -12 -6 118 3640
use L1M1_CDNS_52468879185821  L1M1_CDNS_52468879185821_56
timestamp 1707688321
transform 1 0 9813 0 1 9505
box -12 -6 118 3640
use L1M1_CDNS_52468879185821  L1M1_CDNS_52468879185821_57
timestamp 1707688321
transform 1 0 10733 0 1 9505
box -12 -6 118 3640
use L1M1_CDNS_52468879185821  L1M1_CDNS_52468879185821_58
timestamp 1707688321
transform 1 0 11653 0 1 9505
box -12 -6 118 3640
use L1M1_CDNS_52468879185821  L1M1_CDNS_52468879185821_59
timestamp 1707688321
transform 1 0 12573 0 1 9505
box -12 -6 118 3640
use L1M1_CDNS_52468879185822  L1M1_CDNS_52468879185822_0
timestamp 1707688321
transform 1 0 12573 0 1 37105
box -12 -6 118 1912
use L1M1_CDNS_52468879185822  L1M1_CDNS_52468879185822_1
timestamp 1707688321
transform 1 0 11653 0 1 37105
box -12 -6 118 1912
use L1M1_CDNS_52468879185822  L1M1_CDNS_52468879185822_2
timestamp 1707688321
transform 1 0 10733 0 1 37105
box -12 -6 118 1912
use L1M1_CDNS_52468879185822  L1M1_CDNS_52468879185822_3
timestamp 1707688321
transform 1 0 9813 0 1 37105
box -12 -6 118 1912
use L1M1_CDNS_52468879185822  L1M1_CDNS_52468879185822_4
timestamp 1707688321
transform 1 0 8893 0 1 37105
box -12 -6 118 1912
use L1M1_CDNS_52468879185822  L1M1_CDNS_52468879185822_5
timestamp 1707688321
transform 1 0 7973 0 1 37105
box -12 -6 118 1912
use L1M1_CDNS_52468879185822  L1M1_CDNS_52468879185822_6
timestamp 1707688321
transform 1 0 7053 0 1 37105
box -12 -6 118 1912
use L1M1_CDNS_52468879185822  L1M1_CDNS_52468879185822_7
timestamp 1707688321
transform 1 0 6133 0 1 37105
box -12 -6 118 1912
use L1M1_CDNS_52468879185822  L1M1_CDNS_52468879185822_8
timestamp 1707688321
transform 1 0 5213 0 1 37105
box -12 -6 118 1912
use L1M1_CDNS_52468879185822  L1M1_CDNS_52468879185822_9
timestamp 1707688321
transform 1 0 4293 0 1 37105
box -12 -6 118 1912
use L1M1_CDNS_52468879185822  L1M1_CDNS_52468879185822_10
timestamp 1707688321
transform 1 0 3373 0 1 37105
box -12 -6 118 1912
use M2M3_C_CDNS_524688791859  M2M3_C_CDNS_524688791859_0
timestamp 1707688321
transform 1 0 8683 0 1 37536
box -1077 -437 1077 437
use M2M3_C_CDNS_5246887918510  M2M3_C_CDNS_5246887918510_0
timestamp 1707688321
transform 1 0 11112 0 1 37536
box -1157 -437 1157 437
use M2M3_C_CDNS_5246887918511  M2M3_C_CDNS_5246887918511_0
timestamp 1707688321
transform 1 0 9978 0 1 20026
box -197 -397 197 397
use M2M3_C_CDNS_5246887918512  M2M3_C_CDNS_5246887918512_0
timestamp 1707688321
transform 1 0 8805 0 1 19288
box -237 -597 237 597
use nfet_CDNS_52468879185830  nfet_CDNS_52468879185830_0
timestamp 1707688321
transform 1 0 5017 0 1 18636
box -305 -32 8167 4032
use nfet_CDNS_52468879185830  nfet_CDNS_52468879185830_1
timestamp 1707688321
transform 1 0 5017 0 1 23236
box -305 -32 8167 4032
use nfet_CDNS_52468879185830  nfet_CDNS_52468879185830_2
timestamp 1707688321
transform 1 0 5017 0 1 14036
box -305 -32 8167 4032
use nfet_CDNS_52468879185833  nfet_CDNS_52468879185833_0
timestamp 1707688321
transform 1 0 3177 0 1 27836
box -305 -32 10007 4032
use nfet_CDNS_52468879185833  nfet_CDNS_52468879185833_1
timestamp 1707688321
transform 1 0 3177 0 1 32436
box -305 -32 10007 4032
use nfet_CDNS_52468879185833  nfet_CDNS_52468879185833_2
timestamp 1707688321
transform 1 0 3177 0 1 9436
box -305 -32 10007 4032
use nfet_CDNS_52468879185834  nfet_CDNS_52468879185834_0
timestamp 1707688321
transform 1 0 3177 0 1 37036
box -305 -32 10007 2032
use nfet_CDNS_52468879185837  nfet_CDNS_52468879185837_0
timestamp 1707688321
transform 1 0 10983 0 1 6516
box -79 -26 2363 1426
use pfet_CDNS_52468879185826  pfet_CDNS_52468879185826_0
timestamp 1707688321
transform 1 0 1268 0 1 5960
box -119 -66 7863 1466
use PYbentRes_CDNS_52468879185827  PYbentRes_CDNS_52468879185827_0
timestamp 1707688321
transform 0 1 1672 1 0 8688
box -50 -1458 30933 66
use PYbentRes_CDNS_52468879185828  PYbentRes_CDNS_52468879185828_0
timestamp 1707688321
transform 0 -1 1966 1 0 14871
box -50 -1782 11598 66
use PYbentRes_CDNS_52468879185829  PYbentRes_CDNS_52468879185829_0
timestamp 1707688321
transform 0 -1 14211 1 0 8603
box -50 -324 31297 66
use sky130_fd_io__esd_rcclamp_nfetcap  sky130_fd_io__esd_rcclamp_nfetcap_0
array 0 4 1952 0 2 1244
timestamp 1707688321
transform -1 0 13694 0 -1 4311
box -40 -8 1998 1322
use sky130_fd_io__sio_clamp_Pcap_4x5  sky130_fd_io__sio_clamp_Pcap_4x5_0
timestamp 1707688321
transform -1 0 13744 0 -1 5573
box 10 10 1248 1340
use sky130_fd_io__sio_clamp_Pcap_4x5  sky130_fd_io__sio_clamp_Pcap_4x5_1
array 0 0 0 0 2 1244
timestamp 1707688321
transform -1 0 3984 0 -1 4329
box 10 10 1248 1340
<< labels >>
flabel comment s 10245 4347 10245 4347 0 FreeSans 400 0 0 0 condiode
flabel comment s 13675 39535 13675 39535 0 FreeSans 400 0 0 0 condiode
flabel comment s 12954 8167 12954 8167 0 FreeSans 400 0 0 0 condiode
flabel comment s 10245 9062 10245 9062 0 FreeSans 400 0 0 0 condiode
flabel metal3 s 5179 0 7379 148 2 FreeSans 96 90 0 0 src_bdy_hvc
port 2 nsew ground bidirectional
flabel metal3 s 7578 0 9778 318 0 FreeSans 96 0 0 0 drn_hvc
port 3 nsew power bidirectional
flabel metal2 s 5179 0 5579 107 2 FreeSans 1000 90 0 0 ogc_hvc
port 4 nsew power bidirectional
flabel metal2 s 99 0 4879 148 2 FreeSans 44 90 0 0 src_bdy_hvc
port 2 nsew ground bidirectional
flabel metal2 s 10078 0 14858 148 2 FreeSans 44 90 0 0 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 99 0 4879 411 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 495 4879 499 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 183 481 4879 495 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 169 467 4879 481 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 155 453 4879 467 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 141 439 4879 453 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 127 425 4879 439 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 113 411 4879 425 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 499 4879 1719 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 2475 5635 2480 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 2461 5621 2475 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 2447 5607 2461 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 2433 5593 2447 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 2419 5579 2433 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 2405 5565 2419 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 2391 5551 2405 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 2377 5537 2391 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 2363 5523 2377 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 2349 5509 2363 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 2335 5495 2349 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 2321 5481 2335 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 2307 5467 2321 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 2293 5453 2307 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 2279 5439 2293 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 2265 5425 2279 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 2251 5411 2265 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 2237 5397 2251 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 2223 5383 2237 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 2209 5369 2223 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 2195 5355 2209 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 2181 5341 2195 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 2167 5327 2181 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 2153 5313 2167 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 2139 5299 2153 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 2125 5285 2139 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 2111 5271 2125 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 2097 5257 2111 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 2083 5243 2097 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 2069 5229 2083 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 2055 5215 2069 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 2041 5201 2055 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 2027 5187 2041 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 2013 5173 2027 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 1999 5159 2013 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 1985 5145 1999 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 1971 5131 1985 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 1957 5117 1971 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 1943 5103 1957 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 1929 5089 1943 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 1915 5075 1929 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 1901 5061 1915 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 1887 5047 1901 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 1873 5033 1887 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 1859 5019 1873 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 1845 5005 1859 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 1831 4991 1845 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 1817 4977 1831 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 1803 4963 1817 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 1789 4949 1803 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 1775 4935 1789 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 1761 4921 1775 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 1747 4907 1761 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 1733 4893 1747 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 1719 4879 1733 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 2480 7379 5140 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 5854 3041 5863 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 5840 3050 5854 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 5826 3064 5840 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 5812 3078 5826 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 5798 3092 5812 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 5784 3106 5798 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 5770 3120 5784 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 5756 3134 5770 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 5742 3148 5756 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 5728 3162 5742 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 5714 3176 5728 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 5700 3190 5714 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 5686 3204 5700 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 5672 3218 5686 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 5658 3232 5672 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 5644 3246 5658 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 5630 3260 5644 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 5616 3274 5630 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 5602 3288 5616 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 5588 3302 5602 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 5574 3316 5588 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 5560 3330 5574 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 5546 3344 5560 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 5532 3358 5546 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 5518 3372 5532 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 5504 3386 5518 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 5490 3400 5504 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 5476 3414 5490 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 5462 3428 5476 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 5448 3442 5462 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 5434 3456 5448 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 5420 3470 5434 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 5406 3484 5420 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 5392 3498 5406 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 5378 3512 5392 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 5364 3526 5378 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 5350 3540 5364 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 5336 3554 5350 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 5322 3568 5336 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 5308 3582 5322 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 5294 3596 5308 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 5280 3610 5294 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 5266 3624 5280 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 5252 3638 5266 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 5238 3652 5252 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 5224 3666 5238 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 5210 3680 5224 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 5196 3694 5210 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 5182 3708 5196 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 5168 3722 5182 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 5154 3736 5168 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 5140 3750 5154 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 5863 3041 7133 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 7133 3041 7147 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 7147 3055 7161 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 7161 3069 7175 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 7175 3083 7189 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 7189 3097 7203 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 7203 3111 7217 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 7217 3125 7231 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 7231 3139 7245 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 7245 3153 7259 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 7259 3167 7273 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 7273 3181 7287 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 7287 3195 7301 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 7301 3209 7315 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 7315 3223 7329 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 7329 3237 7343 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 7343 3251 7357 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 7357 3265 7371 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 7371 3279 7385 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 7385 3293 7399 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 7399 3307 7413 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 7413 3321 7427 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 7427 3335 7441 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 7441 3349 7455 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 7455 3363 7469 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 7469 3377 7483 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 7483 3391 7497 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 7497 3405 7511 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 7511 3419 7525 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 7525 3433 7539 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 7539 3447 7553 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 7553 3461 7567 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 7567 3475 7581 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 7581 3489 7595 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 7595 3503 7609 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 7609 3517 7623 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 7623 3531 7637 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 7637 3545 7651 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 7651 3559 7665 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 7665 3573 7679 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 7679 3587 7693 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 7693 3601 7707 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 7707 3615 7721 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 7721 3629 7735 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 7735 3643 7749 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 7749 3657 7763 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 7763 3671 7777 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 7777 3685 7791 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 7791 3699 7805 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 7805 3713 7819 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 7819 3727 7833 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 7833 3741 7847 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 7847 3755 7861 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 7861 3769 7875 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 7875 3783 7889 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 7889 3797 7903 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 7903 3811 7917 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 7917 3825 7931 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 7931 3839 7945 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 7945 3853 7959 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 7959 3867 7973 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 7973 3881 7987 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 7987 3895 8001 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 8001 3909 8015 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 8015 3923 8029 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 8029 3937 8043 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 8043 3951 8057 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 8057 3965 8070 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 10934 7223 11383 7651 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 10654 7931 11383 7933 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 10668 7917 11383 7931 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 10682 7903 11383 7917 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 10696 7889 11383 7903 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 10710 7875 11383 7889 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 10724 7861 11383 7875 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 10738 7847 11383 7861 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 10752 7833 11383 7847 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 10766 7819 11383 7833 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 10780 7805 11383 7819 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 10794 7791 11383 7805 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 10808 7777 11383 7791 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 10822 7763 11383 7777 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 10836 7749 11383 7763 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 10850 7735 11383 7749 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 10864 7721 11383 7735 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 10878 7707 11383 7721 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 10892 7693 11383 7707 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 10906 7679 11383 7693 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 10920 7665 11383 7679 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 10934 7651 11383 7665 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 10526 8059 11246 8070 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 10540 8045 11257 8059 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 10554 8031 11271 8045 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 10568 8017 11285 8031 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 10582 8003 11299 8017 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 10596 7989 11313 8003 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 10610 7975 11327 7989 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 10624 7961 11341 7975 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 10638 7947 11355 7961 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 10652 7933 11369 7947 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 8462 10840 8476 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 8448 10854 8462 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 8434 10868 8448 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 8420 10882 8434 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 8406 10896 8420 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 8392 10910 8406 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 8378 10924 8392 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 8364 10938 8378 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 8350 10952 8364 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 8336 10966 8350 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 8322 10980 8336 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 8308 10994 8322 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 8294 11008 8308 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 8280 11022 8294 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 8266 11036 8280 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 8252 11050 8266 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 8238 11064 8252 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 8224 11078 8238 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 8210 11092 8224 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 8196 11106 8210 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 8182 11120 8196 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 8168 11134 8182 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 8154 11148 8168 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 8140 11162 8154 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 8126 11176 8140 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 8112 11190 8126 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 8098 11204 8112 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 8084 11218 8098 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 8070 11232 8084 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 9050 2824 9063 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 9036 2837 9050 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 9022 2851 9036 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 9008 2865 9022 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 8994 2879 9008 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 8980 2893 8994 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 8966 2907 8980 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 8952 2921 8966 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 8938 2935 8952 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 8924 2949 8938 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 8910 2963 8924 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 8896 2977 8910 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 8882 2991 8896 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 8868 3005 8882 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 8854 3019 8868 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 8840 3033 8854 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 8826 3047 8840 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 8812 3061 8826 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 8798 3075 8812 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 8784 3089 8798 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 8770 3103 8784 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 8756 3117 8770 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 8742 3131 8756 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 8728 3145 8742 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 8714 3159 8728 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 8700 3173 8714 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 8686 3187 8700 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 8672 3201 8686 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 8658 3215 8672 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 8644 3229 8658 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 8630 3243 8644 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 8616 3257 8630 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 8602 3271 8616 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 8588 3285 8602 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 8574 3299 8588 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 8560 3313 8574 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 8546 3327 8560 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 8532 3341 8546 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 8518 3355 8532 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 8504 3369 8518 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 8490 3383 8504 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 8476 3397 8490 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 9063 2824 10843 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 11543 3524 11556 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 11529 3510 11543 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 11515 3496 11529 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 11501 3482 11515 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 11487 3468 11501 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 11473 3454 11487 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 11459 3440 11473 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 11445 3426 11459 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 11431 3412 11445 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 11417 3398 11431 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 11403 3384 11417 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 11389 3370 11403 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 11375 3356 11389 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 11361 3342 11375 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 11347 3328 11361 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 11333 3314 11347 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 11319 3300 11333 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 11305 3286 11319 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 11291 3272 11305 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 11277 3258 11291 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 11263 3244 11277 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 11249 3230 11263 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 11235 3216 11249 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 11221 3202 11235 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 11207 3188 11221 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 11193 3174 11207 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 11179 3160 11193 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 11165 3146 11179 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 11151 3132 11165 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 11137 3118 11151 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 11123 3104 11137 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 11109 3090 11123 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 11095 3076 11109 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 11081 3062 11095 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 11067 3048 11081 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 11053 3034 11067 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 11039 3020 11053 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 11025 3006 11039 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 11011 2992 11025 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 10997 2978 11011 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 10983 2964 10997 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 10969 2950 10983 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 10955 2936 10969 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 10941 2922 10955 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 10927 2908 10941 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 10913 2894 10927 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 10899 2880 10913 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 10885 2866 10899 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 10871 2852 10885 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 10857 2838 10871 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 10843 2824 10857 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 11556 11342 13296 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 13996 2824 14005 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 13982 2833 13996 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 13968 2847 13982 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 13954 2861 13968 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 13940 2875 13954 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 13926 2889 13940 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 13912 2903 13926 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 13898 2917 13912 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 13884 2931 13898 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 13870 2945 13884 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 13856 2959 13870 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 13842 2973 13856 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 13828 2987 13842 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 13814 3001 13828 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 13800 3015 13814 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 13786 3029 13800 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 13772 3043 13786 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 13758 3057 13772 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 13744 3071 13758 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 13730 3085 13744 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 13716 3099 13730 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 13702 3113 13716 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 13688 3127 13702 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 13674 3141 13688 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 13660 3155 13674 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 13646 3169 13660 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 13632 3183 13646 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 13618 3197 13632 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 13604 3211 13618 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 13590 3225 13604 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 13576 3239 13590 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 13562 3253 13576 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 13548 3267 13562 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 13534 3281 13548 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 13520 3295 13534 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 13506 3309 13520 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 13492 3323 13506 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 13478 3337 13492 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 13464 3351 13478 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 13450 3365 13464 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 13436 3379 13450 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 13422 3393 13436 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 13408 3407 13422 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 13394 3421 13408 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 13380 3435 13394 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 13366 3449 13380 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 13352 3463 13366 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 13338 3477 13352 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 13324 3491 13338 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 13310 3505 13324 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 13296 3519 13310 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 14005 2824 15448 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 16148 3524 16156 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 16134 3510 16148 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 16120 3496 16134 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 16106 3482 16120 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 16092 3468 16106 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 16078 3454 16092 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 16064 3440 16078 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 16050 3426 16064 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 16036 3412 16050 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 16022 3398 16036 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 16008 3384 16022 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 15994 3370 16008 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 15980 3356 15994 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 15966 3342 15980 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 15952 3328 15966 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 15938 3314 15952 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 15924 3300 15938 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 15910 3286 15924 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 15896 3272 15910 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 15882 3258 15896 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 15868 3244 15882 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 15854 3230 15868 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 15840 3216 15854 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 15826 3202 15840 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 15812 3188 15826 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 15798 3174 15812 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 15784 3160 15798 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 15770 3146 15784 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 15756 3132 15770 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 15742 3118 15756 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 15728 3104 15742 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 15714 3090 15728 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 15700 3076 15714 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 15686 3062 15700 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 15672 3048 15686 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 15658 3034 15672 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 15644 3020 15658 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 15630 3006 15644 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 15616 2992 15630 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 15602 2978 15616 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 15588 2964 15602 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 15574 2950 15588 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 15560 2936 15574 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 15546 2922 15560 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 15532 2908 15546 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 15518 2894 15532 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 15504 2880 15518 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 15490 2866 15504 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 15476 2852 15490 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 15462 2838 15476 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 15448 2824 15462 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 16156 11341 17896 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 18596 2824 18605 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 18582 2833 18596 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 18568 2847 18582 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 18554 2861 18568 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 18540 2875 18554 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 18526 2889 18540 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 18512 2903 18526 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 18498 2917 18512 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 18484 2931 18498 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 18470 2945 18484 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 18456 2959 18470 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 18442 2973 18456 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 18428 2987 18442 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 18414 3001 18428 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 18400 3015 18414 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 18386 3029 18400 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 18372 3043 18386 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 18358 3057 18372 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 18344 3071 18358 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 18330 3085 18344 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 18316 3099 18330 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 18302 3113 18316 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 18288 3127 18302 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 18274 3141 18288 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 18260 3155 18274 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 18246 3169 18260 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 18232 3183 18246 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 18218 3197 18232 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 18204 3211 18218 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 18190 3225 18204 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 18176 3239 18190 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 18162 3253 18176 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 18148 3267 18162 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 18134 3281 18148 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 18120 3295 18134 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 18106 3309 18120 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 18092 3323 18106 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 18078 3337 18092 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 18064 3351 18078 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 18050 3365 18064 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 18036 3379 18050 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 18022 3393 18036 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 18008 3407 18022 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 17994 3421 18008 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 17980 3435 17994 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 17966 3449 17980 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 17952 3463 17966 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 17938 3477 17952 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 17924 3491 17938 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 17910 3505 17924 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 17896 3519 17910 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 18605 2824 20048 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 20748 3524 20756 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 20734 3510 20748 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 20720 3496 20734 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 20706 3482 20720 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 20692 3468 20706 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 20678 3454 20692 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 20664 3440 20678 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 20650 3426 20664 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 20636 3412 20650 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 20622 3398 20636 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 20608 3384 20622 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 20594 3370 20608 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 20580 3356 20594 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 20566 3342 20580 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 20552 3328 20566 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 20538 3314 20552 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 20524 3300 20538 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 20510 3286 20524 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 20496 3272 20510 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 20482 3258 20496 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 20468 3244 20482 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 20454 3230 20468 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 20440 3216 20454 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 20426 3202 20440 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 20412 3188 20426 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 20398 3174 20412 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 20384 3160 20398 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 20370 3146 20384 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 20356 3132 20370 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 20342 3118 20356 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 20328 3104 20342 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 20314 3090 20328 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 20300 3076 20314 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 20286 3062 20300 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 20272 3048 20286 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 20258 3034 20272 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 20244 3020 20258 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 20230 3006 20244 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 20216 2992 20230 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 20202 2978 20216 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 20188 2964 20202 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 20174 2950 20188 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 20160 2936 20174 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 20146 2922 20160 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 20132 2908 20146 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 20118 2894 20132 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 20104 2880 20118 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 20090 2866 20104 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 20076 2852 20090 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 20062 2838 20076 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 20048 2824 20062 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 20756 11341 22496 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 23210 2824 23213 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 23196 2827 23210 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 23182 2841 23196 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 23168 2855 23182 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 23154 2869 23168 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 23140 2883 23154 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 23126 2897 23140 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 23112 2911 23126 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 23098 2925 23112 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 23084 2939 23098 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 23070 2953 23084 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 23056 2967 23070 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 23042 2981 23056 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 23028 2995 23042 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 23014 3009 23028 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 23000 3023 23014 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 22986 3037 23000 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 22972 3051 22986 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 22958 3065 22972 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 22944 3079 22958 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 22930 3093 22944 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 22916 3107 22930 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 22902 3121 22916 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 22888 3135 22902 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 22874 3149 22888 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 22860 3163 22874 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 22846 3177 22860 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 22832 3191 22846 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 22818 3205 22832 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 22804 3219 22818 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 22790 3233 22804 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 22776 3247 22790 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 22762 3261 22776 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 22748 3275 22762 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 22734 3289 22748 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 22720 3303 22734 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 22706 3317 22720 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 22692 3331 22706 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 22678 3345 22692 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 22664 3359 22678 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 22650 3373 22664 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 22636 3387 22650 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 22622 3401 22636 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 22608 3415 22622 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 22594 3429 22608 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 22580 3443 22594 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 22566 3457 22580 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 22552 3471 22566 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 22538 3485 22552 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 22524 3499 22538 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 22510 3513 22524 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 22496 3527 22510 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 23213 2824 24629 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 25343 3538 25356 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 25329 3524 25343 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 25315 3510 25329 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 25301 3496 25315 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 25287 3482 25301 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 25273 3468 25287 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 25259 3454 25273 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 25245 3440 25259 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 25231 3426 25245 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 25217 3412 25231 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 25203 3398 25217 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 25189 3384 25203 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 25175 3370 25189 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 25161 3356 25175 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 25147 3342 25161 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 25133 3328 25147 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 25119 3314 25133 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 25105 3300 25119 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 25091 3286 25105 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 25077 3272 25091 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 25063 3258 25077 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 25049 3244 25063 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 25035 3230 25049 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 25021 3216 25035 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 25007 3202 25021 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 24993 3188 25007 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 24979 3174 24993 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 24965 3160 24979 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 24951 3146 24965 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 24937 3132 24951 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 24923 3118 24937 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 24909 3104 24923 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 24895 3090 24909 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 24881 3076 24895 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 24867 3062 24881 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 24853 3048 24867 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 24839 3034 24853 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 24825 3020 24839 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 24811 3006 24825 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 24797 2992 24811 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 24783 2978 24797 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 24769 2964 24783 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 24755 2950 24769 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 24741 2936 24755 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 24727 2922 24741 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 24713 2908 24727 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 24699 2894 24713 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 24685 2880 24699 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 24671 2866 24685 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 24657 2852 24671 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 24643 2838 24657 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 24629 2824 24643 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 25356 11341 27096 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 27824 2824 27834 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 27810 2834 27824 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 27796 2848 27810 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 27782 2862 27796 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 27768 2876 27782 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 27754 2890 27768 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 27740 2904 27754 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 27726 2918 27740 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 27712 2932 27726 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 27698 2946 27712 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 27684 2960 27698 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 27670 2974 27684 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 27656 2988 27670 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 27642 3002 27656 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 27628 3016 27642 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 27614 3030 27628 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 27600 3044 27614 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 27586 3058 27600 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 27572 3072 27586 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 27558 3086 27572 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 27544 3100 27558 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 27530 3114 27544 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 27516 3128 27530 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 27502 3142 27516 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 27488 3156 27502 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 27474 3170 27488 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 27460 3184 27474 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 27446 3198 27460 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 27432 3212 27446 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 27418 3226 27432 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 27404 3240 27418 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 27390 3254 27404 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 27376 3268 27390 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 27362 3282 27376 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 27348 3296 27362 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 27334 3310 27348 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 27320 3324 27334 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 27306 3338 27320 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 27292 3352 27306 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 27278 3366 27292 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 27264 3380 27278 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 27250 3394 27264 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 27236 3408 27250 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 27222 3422 27236 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 27208 3436 27222 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 27194 3450 27208 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 27180 3464 27194 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 27166 3478 27180 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 27152 3492 27166 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 27138 3506 27152 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 27124 3520 27138 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 27110 3534 27124 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 27096 3548 27110 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 27834 2824 29243 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 29943 3524 29956 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 29929 3510 29943 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 29915 3496 29929 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 29901 3482 29915 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 29887 3468 29901 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 29873 3454 29887 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 29859 3440 29873 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 29845 3426 29859 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 29831 3412 29845 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 29817 3398 29831 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 29803 3384 29817 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 29789 3370 29803 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 29775 3356 29789 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 29761 3342 29775 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 29747 3328 29761 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 29733 3314 29747 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 29719 3300 29733 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 29705 3286 29719 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 29691 3272 29705 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 29677 3258 29691 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 29663 3244 29677 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 29649 3230 29663 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 29635 3216 29649 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 29621 3202 29635 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 29607 3188 29621 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 29593 3174 29607 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 29579 3160 29593 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 29565 3146 29579 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 29551 3132 29565 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 29537 3118 29551 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 29523 3104 29537 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 29509 3090 29523 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 29495 3076 29509 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 29481 3062 29495 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 29467 3048 29481 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 29453 3034 29467 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 29439 3020 29453 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 29425 3006 29439 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 29411 2992 29425 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 29397 2978 29411 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 29383 2964 29397 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 29369 2950 29383 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 29355 2936 29369 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 29341 2922 29355 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 29327 2908 29341 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 29313 2894 29327 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 29299 2880 29313 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 29285 2866 29299 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 29271 2852 29285 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 29257 2838 29271 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 29243 2824 29257 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 29956 11341 31696 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 32410 2824 32416 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 32396 2830 32410 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 32382 2844 32396 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 32368 2858 32382 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 32354 2872 32368 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 32340 2886 32354 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 32326 2900 32340 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 32312 2914 32326 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 32298 2928 32312 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 32284 2942 32298 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 32270 2956 32284 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 32256 2970 32270 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 32242 2984 32256 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 32228 2998 32242 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 32214 3012 32228 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 32200 3026 32214 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 32186 3040 32200 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 32172 3054 32186 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 32158 3068 32172 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 32144 3082 32158 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 32130 3096 32144 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 32116 3110 32130 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 32102 3124 32116 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 32088 3138 32102 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 32074 3152 32088 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 32060 3166 32074 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 32046 3180 32060 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 32032 3194 32046 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 32018 3208 32032 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 32004 3222 32018 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 31990 3236 32004 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 31976 3250 31990 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 31962 3264 31976 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 31948 3278 31962 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 31934 3292 31948 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 31920 3306 31934 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 31906 3320 31920 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 31892 3334 31906 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 31878 3348 31892 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 31864 3362 31878 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 31850 3376 31864 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 31836 3390 31850 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 31822 3404 31836 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 31808 3418 31822 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 31794 3432 31808 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 31780 3446 31794 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 31766 3460 31780 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 31752 3474 31766 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 31738 3488 31752 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 31724 3502 31738 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 31710 3516 31724 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 31696 3530 31710 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 32416 2824 33844 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 34544 3524 34556 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 34530 3510 34544 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 34516 3496 34530 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 34502 3482 34516 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 34488 3468 34502 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 34474 3454 34488 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 34460 3440 34474 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 34446 3426 34460 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 34432 3412 34446 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 34418 3398 34432 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 34404 3384 34418 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 34390 3370 34404 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 34376 3356 34390 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 34362 3342 34376 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 34348 3328 34362 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 34334 3314 34348 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 34320 3300 34334 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 34306 3286 34320 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 34292 3272 34306 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 34278 3258 34292 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 34264 3244 34278 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 34250 3230 34264 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 34236 3216 34250 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 34222 3202 34236 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 34208 3188 34222 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 34194 3174 34208 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 34180 3160 34194 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 34166 3146 34180 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 34152 3132 34166 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 34138 3118 34152 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 34124 3104 34138 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 34110 3090 34124 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 34096 3076 34110 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 34082 3062 34096 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 34068 3048 34082 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 34054 3034 34068 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 34040 3020 34054 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 34026 3006 34040 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 34012 2992 34026 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 33998 2978 34012 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 33984 2964 33998 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 33970 2950 33984 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 33956 2936 33970 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 33942 2922 33956 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 33928 2908 33942 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 33914 2894 33928 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 33900 2880 33914 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 33886 2866 33900 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 33872 2852 33886 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 33858 2838 33872 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 33844 2824 33858 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 34556 11592 36296 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 36758 3064 36771 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 36744 3077 36758 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 36730 3091 36744 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 36716 3105 36730 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 36702 3119 36716 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 36688 3133 36702 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 36674 3147 36688 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 36660 3161 36674 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 36646 3175 36660 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 36632 3189 36646 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 36618 3203 36632 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 36604 3217 36618 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 36590 3231 36604 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 36576 3245 36590 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 36562 3259 36576 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 36548 3273 36562 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 36534 3287 36548 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 36520 3301 36534 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 36506 3315 36520 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 36492 3329 36506 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 36478 3343 36492 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 36464 3357 36478 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 36450 3371 36464 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 36436 3385 36450 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 36422 3399 36436 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 36408 3413 36422 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 36394 3427 36408 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 36380 3441 36394 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 36366 3455 36380 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 36352 3469 36366 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 36338 3483 36352 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 36324 3497 36338 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 36310 3511 36324 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 36296 3525 36310 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 36771 3064 36781 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 37005 2824 37011 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 36991 2830 37005 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 36977 2844 36991 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 36963 2858 36977 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 36949 2872 36963 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 36935 2886 36949 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 36921 2900 36935 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 36907 2914 36921 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 36893 2928 36907 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 36879 2942 36893 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 36865 2956 36879 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 36851 2970 36865 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 36837 2984 36851 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 36823 2998 36837 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 36809 3012 36823 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 36795 3026 36809 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 36781 3040 36795 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 37011 2824 37917 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 38099 3006 38112 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 38085 2992 38099 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 38071 2978 38085 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 38057 2964 38071 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 38043 2950 38057 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 38029 2936 38043 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 38015 2922 38029 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 38001 2908 38015 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 37987 2894 38001 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 37973 2880 37987 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 37959 2866 37973 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 37945 2852 37959 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 37931 2838 37945 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 37917 2824 37931 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 187 38112 13440 39015 1 src_bdy_hvc
port 2 nsew ground bidirectional
rlabel metal2 s 10078 0 14858 1725 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 9350 2453 14858 2459 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 9364 2439 14858 2453 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 9378 2425 14858 2439 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 9392 2411 14858 2425 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 9406 2397 14858 2411 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 9420 2383 14858 2397 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 9434 2369 14858 2383 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 9448 2355 14858 2369 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 9462 2341 14858 2355 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 9476 2327 14858 2341 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 9490 2313 14858 2327 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 9504 2299 14858 2313 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 9518 2285 14858 2299 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 9532 2271 14858 2285 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 9546 2257 14858 2271 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 9560 2243 14858 2257 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 9574 2229 14858 2243 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 9588 2215 14858 2229 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 9602 2201 14858 2215 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 9616 2187 14858 2201 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 9630 2173 14858 2187 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 9644 2159 14858 2173 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 9658 2145 14858 2159 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 9672 2131 14858 2145 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 9686 2117 14858 2131 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 9700 2103 14858 2117 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 9714 2089 14858 2103 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 9728 2075 14858 2089 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 9742 2061 14858 2075 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 9756 2047 14858 2061 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 9770 2033 14858 2047 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 9784 2019 14858 2033 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 9798 2005 14858 2019 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 9812 1991 14858 2005 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 9826 1977 14858 1991 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 9840 1963 14858 1977 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 9854 1949 14858 1963 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 9868 1935 14858 1949 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 9882 1921 14858 1935 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 9896 1907 14858 1921 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 9910 1893 14858 1907 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 9924 1879 14858 1893 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 9938 1865 14858 1879 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 9952 1851 14858 1865 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 9966 1837 14858 1851 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 9980 1823 14858 1837 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 9994 1809 14858 1823 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 10008 1795 14858 1809 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 10022 1781 14858 1795 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 10036 1767 14858 1781 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 10050 1753 14858 1767 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 10064 1739 14858 1753 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 10078 1725 14858 1739 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 7578 2459 14858 5132 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11177 5132 14858 5146 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11191 5146 14858 5160 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11205 5160 14858 5174 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11219 5174 14858 5188 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11233 5188 14858 5202 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11247 5202 14858 5216 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11261 5216 14858 5230 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11275 5230 14858 5244 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11289 5244 14858 5258 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11303 5258 14858 5272 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11317 5272 14858 5286 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11331 5286 14858 5300 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11345 5300 14858 5314 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11359 5314 14858 5328 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11373 5328 14858 5342 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11387 5342 14858 5356 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11401 5356 14858 5370 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11415 5370 14858 5384 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11429 5384 14858 5398 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11443 5398 14858 5412 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11457 5412 14858 5426 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11471 5426 14858 5440 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11485 5440 14858 5454 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11499 5454 14858 5468 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11513 5468 14858 5482 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11527 5482 14858 5496 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11541 5496 14858 5510 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11555 5510 14858 5524 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11569 5524 14858 5538 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11583 5538 14858 5552 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11597 5552 14858 5566 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11611 5566 14858 5580 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11625 5580 14858 5594 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11639 5594 14858 5608 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11653 5608 14858 5622 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11667 5622 14858 5636 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11681 5636 14858 5650 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11695 5650 14858 5664 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11709 5664 14858 5678 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11723 5678 14858 5692 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11737 5692 14858 5706 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11751 5706 14858 5720 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11765 5720 14858 5734 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11779 5734 14858 5748 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11793 5748 14858 5762 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11807 5762 14858 5776 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11821 5776 14858 5790 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11835 5790 14858 5804 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11849 5804 14858 5818 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11863 5818 14858 5832 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11877 5832 14858 5846 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11891 5846 14858 5860 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11905 5860 14858 5874 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11919 5874 14858 5888 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11933 5888 14858 5902 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11947 5902 14858 5916 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11961 5916 14858 5930 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11975 5930 14858 5944 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11989 5944 14858 5958 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 12003 5958 14858 5972 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 12017 5972 14858 5986 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 12031 5986 14858 6000 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 12045 6000 14858 6014 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 12059 6014 14858 6028 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 12073 6028 14858 6042 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 12087 6042 14858 6056 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 12101 6056 14858 6070 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 12115 6070 14858 6084 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 12129 6084 14858 6098 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 12143 6098 14858 6112 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 12157 6112 14858 6126 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 12171 6126 14858 6140 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 12185 6140 14858 6154 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 12199 6154 14858 6168 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 12213 6168 14858 6182 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 12222 6182 14858 6191 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 12222 6191 14858 8764 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11508 9478 14858 9491 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11522 9464 14858 9478 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11536 9450 14858 9464 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11550 9436 14858 9450 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11564 9422 14858 9436 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11578 9408 14858 9422 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11592 9394 14858 9408 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11606 9380 14858 9394 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11620 9366 14858 9380 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11634 9352 14858 9366 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11648 9338 14858 9352 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11662 9324 14858 9338 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11676 9310 14858 9324 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11690 9296 14858 9310 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11704 9282 14858 9296 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11718 9268 14858 9282 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11732 9254 14858 9268 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11746 9240 14858 9254 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11760 9226 14858 9240 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11774 9212 14858 9226 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11788 9198 14858 9212 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11802 9184 14858 9198 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11816 9170 14858 9184 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11830 9156 14858 9170 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11844 9142 14858 9156 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11858 9128 14858 9142 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11872 9114 14858 9128 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11886 9100 14858 9114 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11900 9086 14858 9100 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11914 9072 14858 9086 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11928 9058 14858 9072 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11942 9044 14858 9058 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11956 9030 14858 9044 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11970 9016 14858 9030 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11984 9002 14858 9016 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11998 8988 14858 9002 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 12012 8974 14858 8988 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 12026 8960 14858 8974 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 12040 8946 14858 8960 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 12054 8932 14858 8946 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 12068 8918 14858 8932 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 12082 8904 14858 8918 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 12096 8890 14858 8904 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 12110 8876 14858 8890 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 12124 8862 14858 8876 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 12138 8848 14858 8862 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 12152 8834 14858 8848 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 12166 8820 14858 8834 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 12180 8806 14858 8820 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 12194 8792 14858 8806 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 12208 8778 14858 8792 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 12222 8764 14858 8778 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 3361 9491 14858 10953 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 3770 11219 14858 11231 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 3758 11205 14858 11219 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 3744 11191 14858 11205 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 3730 11177 14858 11191 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 3716 11163 14858 11177 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 3702 11149 14858 11163 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 3688 11135 14858 11149 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 3674 11121 14858 11135 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 3660 11107 14858 11121 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 3646 11093 14858 11107 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 3632 11079 14858 11093 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 3618 11065 14858 11079 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 3604 11051 14858 11065 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 3590 11037 14858 11051 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 3576 11023 14858 11037 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 3562 11009 14858 11023 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 3548 10995 14858 11009 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 3534 10981 14858 10995 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 3520 10967 14858 10981 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 3506 10953 14858 10967 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 12222 11945 14858 11948 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 12219 11931 14858 11945 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 12205 11917 14858 11931 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 12191 11903 14858 11917 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 12177 11889 14858 11903 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 12163 11875 14858 11889 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 12149 11861 14858 11875 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 12135 11847 14858 11861 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 12121 11833 14858 11847 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 12107 11819 14858 11833 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 12093 11805 14858 11819 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 12079 11791 14858 11805 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 12065 11777 14858 11791 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 12051 11763 14858 11777 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 12037 11749 14858 11763 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 12023 11735 14858 11749 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 12009 11721 14858 11735 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11995 11707 14858 11721 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11981 11693 14858 11707 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11967 11679 14858 11693 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11953 11665 14858 11679 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11939 11651 14858 11665 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11925 11637 14858 11651 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11911 11623 14858 11637 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11897 11609 14858 11623 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11883 11595 14858 11609 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11869 11581 14858 11595 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11855 11567 14858 11581 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11841 11553 14858 11567 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11827 11539 14858 11553 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11813 11525 14858 11539 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11799 11511 14858 11525 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11785 11497 14858 11511 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11771 11483 14858 11497 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11757 11469 14858 11483 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11743 11455 14858 11469 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11729 11441 14858 11455 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11715 11427 14858 11441 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11701 11413 14858 11427 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11687 11399 14858 11413 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11673 11385 14858 11399 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11659 11371 14858 11385 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11645 11357 14858 11371 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11631 11343 14858 11357 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11617 11329 14858 11343 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11603 11315 14858 11329 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11589 11301 14858 11315 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11575 11287 14858 11301 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11561 11273 14858 11287 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11547 11259 14858 11273 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11533 11245 14858 11259 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11519 11231 14858 11245 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 12222 11948 14858 13370 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11508 14084 14858 14091 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11522 14070 14858 14084 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11536 14056 14858 14070 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11550 14042 14858 14056 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11564 14028 14858 14042 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11578 14014 14858 14028 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11592 14000 14858 14014 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11606 13986 14858 14000 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11620 13972 14858 13986 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11634 13958 14858 13972 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11648 13944 14858 13958 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11662 13930 14858 13944 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11676 13916 14858 13930 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11690 13902 14858 13916 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11704 13888 14858 13902 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11718 13874 14858 13888 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11732 13860 14858 13874 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11746 13846 14858 13860 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11760 13832 14858 13846 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11774 13818 14858 13832 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11788 13804 14858 13818 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11802 13790 14858 13804 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11816 13776 14858 13790 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11830 13762 14858 13776 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11844 13748 14858 13762 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11858 13734 14858 13748 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11872 13720 14858 13734 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11886 13706 14858 13720 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11900 13692 14858 13706 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11914 13678 14858 13692 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11928 13664 14858 13678 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11942 13650 14858 13664 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11956 13636 14858 13650 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11970 13622 14858 13636 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11984 13608 14858 13622 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11998 13594 14858 13608 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 12012 13580 14858 13594 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 12026 13566 14858 13580 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 12040 13552 14858 13566 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 12054 13538 14858 13552 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 12068 13524 14858 13538 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 12082 13510 14858 13524 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 12096 13496 14858 13510 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 12110 13482 14858 13496 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 12124 13468 14858 13482 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 12138 13454 14858 13468 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 12152 13440 14858 13454 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 12166 13426 14858 13440 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 12180 13412 14858 13426 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 12194 13398 14858 13412 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 12208 13384 14858 13398 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 12222 13370 14858 13384 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 4964 14091 14858 14597 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 4740 14821 14858 14831 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 4754 14807 14858 14821 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 4768 14793 14858 14807 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 4782 14779 14858 14793 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 4796 14765 14858 14779 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 4810 14751 14858 14765 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 4824 14737 14858 14751 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 4838 14723 14858 14737 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 4852 14709 14858 14723 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 4866 14695 14858 14709 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 4880 14681 14858 14695 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 4894 14667 14858 14681 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 4908 14653 14858 14667 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 4922 14639 14858 14653 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 4936 14625 14858 14639 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 4950 14611 14858 14625 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 4964 14597 14858 14611 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 3682 14831 14858 14883 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 4964 15121 14858 15123 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 4962 15107 14858 15121 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 4948 15093 14858 15107 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 4934 15079 14858 15093 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 4920 15065 14858 15079 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 4906 15051 14858 15065 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 4892 15037 14858 15051 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 4878 15023 14858 15037 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 4864 15009 14858 15023 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 4850 14995 14858 15009 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 4836 14981 14858 14995 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 4822 14967 14858 14981 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 4808 14953 14858 14967 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 4794 14939 14858 14953 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 4780 14925 14858 14939 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 4766 14911 14858 14925 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 4752 14897 14858 14911 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 4738 14883 14858 14897 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 4964 15123 14858 15831 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 12222 16531 14858 16542 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 12211 16517 14858 16531 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 12197 16503 14858 16517 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 12183 16489 14858 16503 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 12169 16475 14858 16489 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 12155 16461 14858 16475 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 12141 16447 14858 16461 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 12127 16433 14858 16447 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 12113 16419 14858 16433 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 12099 16405 14858 16419 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 12085 16391 14858 16405 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 12071 16377 14858 16391 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 12057 16363 14858 16377 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 12043 16349 14858 16363 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 12029 16335 14858 16349 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 12015 16321 14858 16335 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 12001 16307 14858 16321 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11987 16293 14858 16307 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11973 16279 14858 16293 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11959 16265 14858 16279 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11945 16251 14858 16265 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11931 16237 14858 16251 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11917 16223 14858 16237 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11903 16209 14858 16223 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11889 16195 14858 16209 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11875 16181 14858 16195 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11861 16167 14858 16181 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11847 16153 14858 16167 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11833 16139 14858 16153 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11819 16125 14858 16139 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11805 16111 14858 16125 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11791 16097 14858 16111 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11777 16083 14858 16097 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11763 16069 14858 16083 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11749 16055 14858 16069 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11735 16041 14858 16055 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11721 16027 14858 16041 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11707 16013 14858 16027 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11693 15999 14858 16013 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11679 15985 14858 15999 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11665 15971 14858 15985 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11651 15957 14858 15971 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11637 15943 14858 15957 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11623 15929 14858 15943 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11609 15915 14858 15929 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11595 15901 14858 15915 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11581 15887 14858 15901 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11567 15873 14858 15887 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11553 15859 14858 15873 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11539 15845 14858 15859 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11525 15831 14858 15845 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 12222 16542 14858 17982 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11522 18682 14858 18691 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11536 18668 14858 18682 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11550 18654 14858 18668 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11564 18640 14858 18654 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11578 18626 14858 18640 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11592 18612 14858 18626 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11606 18598 14858 18612 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11620 18584 14858 18598 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11634 18570 14858 18584 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11648 18556 14858 18570 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11662 18542 14858 18556 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11676 18528 14858 18542 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11690 18514 14858 18528 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11704 18500 14858 18514 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11718 18486 14858 18500 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11732 18472 14858 18486 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11746 18458 14858 18472 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11760 18444 14858 18458 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11774 18430 14858 18444 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11788 18416 14858 18430 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11802 18402 14858 18416 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11816 18388 14858 18402 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11830 18374 14858 18388 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11844 18360 14858 18374 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11858 18346 14858 18360 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11872 18332 14858 18346 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11886 18318 14858 18332 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11900 18304 14858 18318 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11914 18290 14858 18304 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11928 18276 14858 18290 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11942 18262 14858 18276 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11956 18248 14858 18262 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11970 18234 14858 18248 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11984 18220 14858 18234 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11998 18206 14858 18220 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 12012 18192 14858 18206 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 12026 18178 14858 18192 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 12040 18164 14858 18178 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 12054 18150 14858 18164 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 12068 18136 14858 18150 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 12082 18122 14858 18136 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 12096 18108 14858 18122 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 12110 18094 14858 18108 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 12124 18080 14858 18094 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 12138 18066 14858 18080 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 12152 18052 14858 18066 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 12166 18038 14858 18052 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 12180 18024 14858 18038 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 12194 18010 14858 18024 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 12208 17996 14858 18010 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 12222 17982 14858 17996 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 4964 18691 14858 20431 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 12222 21131 14858 21142 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 12211 21117 14858 21131 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 12197 21103 14858 21117 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 12183 21089 14858 21103 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 12169 21075 14858 21089 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 12155 21061 14858 21075 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 12141 21047 14858 21061 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 12127 21033 14858 21047 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 12113 21019 14858 21033 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 12099 21005 14858 21019 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 12085 20991 14858 21005 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 12071 20977 14858 20991 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 12057 20963 14858 20977 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 12043 20949 14858 20963 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 12029 20935 14858 20949 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 12015 20921 14858 20935 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 12001 20907 14858 20921 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11987 20893 14858 20907 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11973 20879 14858 20893 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11959 20865 14858 20879 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11945 20851 14858 20865 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11931 20837 14858 20851 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11917 20823 14858 20837 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11903 20809 14858 20823 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11889 20795 14858 20809 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11875 20781 14858 20795 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11861 20767 14858 20781 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11847 20753 14858 20767 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11833 20739 14858 20753 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11819 20725 14858 20739 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11805 20711 14858 20725 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11791 20697 14858 20711 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11777 20683 14858 20697 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11763 20669 14858 20683 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11749 20655 14858 20669 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11735 20641 14858 20655 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11721 20627 14858 20641 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11707 20613 14858 20627 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11693 20599 14858 20613 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11679 20585 14858 20599 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11665 20571 14858 20585 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11651 20557 14858 20571 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11637 20543 14858 20557 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11623 20529 14858 20543 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11609 20515 14858 20529 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11595 20501 14858 20515 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11581 20487 14858 20501 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11567 20473 14858 20487 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11553 20459 14858 20473 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11539 20445 14858 20459 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11525 20431 14858 20445 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 12222 21142 14858 22564 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11508 23278 14858 23291 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11522 23264 14858 23278 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11536 23250 14858 23264 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11550 23236 14858 23250 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11564 23222 14858 23236 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11578 23208 14858 23222 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11592 23194 14858 23208 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11606 23180 14858 23194 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11620 23166 14858 23180 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11634 23152 14858 23166 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11648 23138 14858 23152 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11662 23124 14858 23138 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11676 23110 14858 23124 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11690 23096 14858 23110 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11704 23082 14858 23096 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11718 23068 14858 23082 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11732 23054 14858 23068 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11746 23040 14858 23054 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11760 23026 14858 23040 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11774 23012 14858 23026 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11788 22998 14858 23012 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11802 22984 14858 22998 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11816 22970 14858 22984 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11830 22956 14858 22970 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11844 22942 14858 22956 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11858 22928 14858 22942 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11872 22914 14858 22928 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11886 22900 14858 22914 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11900 22886 14858 22900 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11914 22872 14858 22886 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11928 22858 14858 22872 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11942 22844 14858 22858 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11956 22830 14858 22844 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11970 22816 14858 22830 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11984 22802 14858 22816 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11998 22788 14858 22802 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 12012 22774 14858 22788 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 12026 22760 14858 22774 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 12040 22746 14858 22760 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 12054 22732 14858 22746 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 12068 22718 14858 22732 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 12082 22704 14858 22718 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 12096 22690 14858 22704 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 12110 22676 14858 22690 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 12124 22662 14858 22676 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 12138 22648 14858 22662 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 12152 22634 14858 22648 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 12166 22620 14858 22634 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 12180 22606 14858 22620 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 12194 22592 14858 22606 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 12208 22578 14858 22592 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 12222 22564 14858 22578 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 4964 23291 14858 25031 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 12222 25731 14858 25742 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 12211 25717 14858 25731 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 12197 25703 14858 25717 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 12183 25689 14858 25703 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 12169 25675 14858 25689 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 12155 25661 14858 25675 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 12141 25647 14858 25661 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 12127 25633 14858 25647 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 12113 25619 14858 25633 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 12099 25605 14858 25619 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 12085 25591 14858 25605 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 12071 25577 14858 25591 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 12057 25563 14858 25577 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 12043 25549 14858 25563 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 12029 25535 14858 25549 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 12015 25521 14858 25535 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 12001 25507 14858 25521 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11987 25493 14858 25507 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11973 25479 14858 25493 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11959 25465 14858 25479 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11945 25451 14858 25465 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11931 25437 14858 25451 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11917 25423 14858 25437 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11903 25409 14858 25423 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11889 25395 14858 25409 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11875 25381 14858 25395 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11861 25367 14858 25381 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11847 25353 14858 25367 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11833 25339 14858 25353 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11819 25325 14858 25339 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11805 25311 14858 25325 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11791 25297 14858 25311 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11777 25283 14858 25297 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11763 25269 14858 25283 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11749 25255 14858 25269 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11735 25241 14858 25255 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11721 25227 14858 25241 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11707 25213 14858 25227 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11693 25199 14858 25213 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11679 25185 14858 25199 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11665 25171 14858 25185 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11651 25157 14858 25171 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11637 25143 14858 25157 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11623 25129 14858 25143 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11609 25115 14858 25129 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11595 25101 14858 25115 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11581 25087 14858 25101 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11567 25073 14858 25087 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11553 25059 14858 25073 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11539 25045 14858 25059 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11525 25031 14858 25045 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 12222 25742 14858 27171 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11508 27885 14858 27891 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11522 27871 14858 27885 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11536 27857 14858 27871 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11550 27843 14858 27857 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11564 27829 14858 27843 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11578 27815 14858 27829 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11592 27801 14858 27815 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11606 27787 14858 27801 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11620 27773 14858 27787 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11634 27759 14858 27773 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11648 27745 14858 27759 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11662 27731 14858 27745 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11676 27717 14858 27731 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11690 27703 14858 27717 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11704 27689 14858 27703 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11718 27675 14858 27689 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11732 27661 14858 27675 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11746 27647 14858 27661 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11760 27633 14858 27647 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11774 27619 14858 27633 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11788 27605 14858 27619 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11802 27591 14858 27605 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11816 27577 14858 27591 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11830 27563 14858 27577 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11844 27549 14858 27563 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11858 27535 14858 27549 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11872 27521 14858 27535 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11886 27507 14858 27521 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11900 27493 14858 27507 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11914 27479 14858 27493 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11928 27465 14858 27479 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11942 27451 14858 27465 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11956 27437 14858 27451 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11970 27423 14858 27437 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11984 27409 14858 27423 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11998 27395 14858 27409 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 12012 27381 14858 27395 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 12026 27367 14858 27381 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 12040 27353 14858 27367 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 12054 27339 14858 27353 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 12068 27325 14858 27339 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 12082 27311 14858 27325 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 12096 27297 14858 27311 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 12110 27283 14858 27297 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 12124 27269 14858 27283 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 12138 27255 14858 27269 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 12152 27241 14858 27255 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 12166 27227 14858 27241 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 12180 27213 14858 27227 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 12194 27199 14858 27213 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 12208 27185 14858 27199 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 12222 27171 14858 27185 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 3361 27891 14858 29342 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 3650 29622 14858 29631 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 3641 29608 14858 29622 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 3627 29594 14858 29608 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 3613 29580 14858 29594 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 3599 29566 14858 29580 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 3585 29552 14858 29566 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 3571 29538 14858 29552 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 3557 29524 14858 29538 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 3543 29510 14858 29524 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 3529 29496 14858 29510 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 3515 29482 14858 29496 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 3501 29468 14858 29482 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 3487 29454 14858 29468 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 3473 29440 14858 29454 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 3459 29426 14858 29440 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 3445 29412 14858 29426 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 3431 29398 14858 29412 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 3417 29384 14858 29398 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 3403 29370 14858 29384 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 3389 29356 14858 29370 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 3375 29342 14858 29356 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 12222 30345 14858 30356 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 12211 30331 14858 30345 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 12197 30317 14858 30331 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 12183 30303 14858 30317 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 12169 30289 14858 30303 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 12155 30275 14858 30289 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 12141 30261 14858 30275 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 12127 30247 14858 30261 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 12113 30233 14858 30247 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 12099 30219 14858 30233 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 12085 30205 14858 30219 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 12071 30191 14858 30205 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 12057 30177 14858 30191 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 12043 30163 14858 30177 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 12029 30149 14858 30163 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 12015 30135 14858 30149 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 12001 30121 14858 30135 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11987 30107 14858 30121 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11973 30093 14858 30107 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11959 30079 14858 30093 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11945 30065 14858 30079 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11931 30051 14858 30065 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11917 30037 14858 30051 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11903 30023 14858 30037 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11889 30009 14858 30023 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11875 29995 14858 30009 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11861 29981 14858 29995 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11847 29967 14858 29981 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11833 29953 14858 29967 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11819 29939 14858 29953 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11805 29925 14858 29939 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11791 29911 14858 29925 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11777 29897 14858 29911 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11763 29883 14858 29897 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11749 29869 14858 29883 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11735 29855 14858 29869 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11721 29841 14858 29855 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11707 29827 14858 29841 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11693 29813 14858 29827 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11679 29799 14858 29813 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11665 29785 14858 29799 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11651 29771 14858 29785 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11637 29757 14858 29771 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11623 29743 14858 29757 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11609 29729 14858 29743 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11595 29715 14858 29729 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11581 29701 14858 29715 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11567 29687 14858 29701 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11553 29673 14858 29687 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11539 29659 14858 29673 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11525 29645 14858 29659 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11511 29631 14858 29645 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 12222 30356 14858 31774 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11508 32488 14858 32491 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11522 32474 14858 32488 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11536 32460 14858 32474 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11550 32446 14858 32460 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11564 32432 14858 32446 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11578 32418 14858 32432 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11592 32404 14858 32418 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11606 32390 14858 32404 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11620 32376 14858 32390 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11634 32362 14858 32376 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11648 32348 14858 32362 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11662 32334 14858 32348 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11676 32320 14858 32334 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11690 32306 14858 32320 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11704 32292 14858 32306 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11718 32278 14858 32292 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11732 32264 14858 32278 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11746 32250 14858 32264 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11760 32236 14858 32250 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11774 32222 14858 32236 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11788 32208 14858 32222 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11802 32194 14858 32208 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11816 32180 14858 32194 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11830 32166 14858 32180 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11844 32152 14858 32166 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11858 32138 14858 32152 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11872 32124 14858 32138 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11886 32110 14858 32124 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11900 32096 14858 32110 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11914 32082 14858 32096 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11928 32068 14858 32082 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11942 32054 14858 32068 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11956 32040 14858 32054 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11970 32026 14858 32040 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11984 32012 14858 32026 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11998 31998 14858 32012 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 12012 31984 14858 31998 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 12026 31970 14858 31984 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 12040 31956 14858 31970 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 12054 31942 14858 31956 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 12068 31928 14858 31942 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 12082 31914 14858 31928 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 12096 31900 14858 31914 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 12110 31886 14858 31900 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 12124 31872 14858 31886 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 12138 31858 14858 31872 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 12152 31844 14858 31858 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 12166 31830 14858 31844 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 12180 31816 14858 31830 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 12194 31802 14858 31816 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 12208 31788 14858 31802 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 12222 31774 14858 31788 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 3361 32491 14858 34231 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 12222 34931 14858 34940 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 12213 34917 14858 34931 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 12199 34903 14858 34917 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 12185 34889 14858 34903 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 12171 34875 14858 34889 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 12157 34861 14858 34875 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 12143 34847 14858 34861 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 12129 34833 14858 34847 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 12115 34819 14858 34833 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 12101 34805 14858 34819 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 12087 34791 14858 34805 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 12073 34777 14858 34791 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 12059 34763 14858 34777 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 12045 34749 14858 34763 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 12031 34735 14858 34749 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 12017 34721 14858 34735 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 12003 34707 14858 34721 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11989 34693 14858 34707 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11975 34679 14858 34693 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11961 34665 14858 34679 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11947 34651 14858 34665 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11933 34637 14858 34651 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11919 34623 14858 34637 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11905 34609 14858 34623 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11891 34595 14858 34609 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11877 34581 14858 34595 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11863 34567 14858 34581 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11849 34553 14858 34567 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11835 34539 14858 34553 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11821 34525 14858 34539 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11807 34511 14858 34525 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11793 34497 14858 34511 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11779 34483 14858 34497 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11765 34469 14858 34483 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11751 34455 14858 34469 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11737 34441 14858 34455 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11723 34427 14858 34441 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11709 34413 14858 34427 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11695 34399 14858 34413 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11681 34385 14858 34399 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11667 34371 14858 34385 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11653 34357 14858 34371 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11639 34343 14858 34357 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11625 34329 14858 34343 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11611 34315 14858 34329 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11597 34301 14858 34315 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11583 34287 14858 34301 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11569 34273 14858 34287 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11555 34259 14858 34273 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11541 34245 14858 34259 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11527 34231 14858 34245 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 12222 34940 14858 36576 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11746 37052 14858 37059 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11760 37038 14858 37052 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11774 37024 14858 37038 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11788 37010 14858 37024 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11802 36996 14858 37010 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11816 36982 14858 36996 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11830 36968 14858 36982 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11844 36954 14858 36968 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11858 36940 14858 36954 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11872 36926 14858 36940 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11886 36912 14858 36926 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11900 36898 14858 36912 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11914 36884 14858 36898 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11928 36870 14858 36884 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11942 36856 14858 36870 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11956 36842 14858 36856 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11970 36828 14858 36842 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11984 36814 14858 36828 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 11998 36800 14858 36814 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 12012 36786 14858 36800 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 12026 36772 14858 36786 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 12040 36758 14858 36772 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 12054 36744 14858 36758 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 12068 36730 14858 36744 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 12082 36716 14858 36730 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 12096 36702 14858 36716 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 12110 36688 14858 36702 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 12124 36674 14858 36688 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 12138 36660 14858 36674 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 12152 36646 14858 36660 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 12166 36632 14858 36646 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 12180 36618 14858 36632 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 12194 36604 14858 36618 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 12208 36590 14858 36604 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 12222 36576 14858 36590 1 drn_hvc
port 3 nsew power bidirectional
rlabel metal2 s 3124 37059 14858 38003 1 drn_hvc
port 3 nsew power bidirectional
<< properties >>
string FIXED_BBOX 0 0 15000 40000
string GDS_END 42927674
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 39132556
string LEFclass BLOCK
string LEFsymmetry R90
string path 171.875 865.850 171.875 868.725 
<< end >>
