magic
tech sky130B
magscale 1 2
timestamp 1707688321
<< obsli1 >>
rect 224 26 95503 50717
<< obsm1 >>
rect 292 14 95509 50729
<< metal2 >>
rect 17052 0 17221 5923
rect 17249 0 17419 4895
rect 21342 0 21394 270
rect 22018 0 22070 3493
rect 24291 0 24343 9204
rect 25625 0 25677 2035
rect 27035 0 27087 5790
rect 27115 0 27167 7338
rect 28240 0 28309 417
rect 28401 0 28453 1394
rect 28481 0 28533 1996
rect 29443 0 29495 5384
rect 29523 0 29575 9105
rect 29961 0 30013 5650
rect 30682 592 30734 6989
rect 30682 0 30734 456
rect 30762 0 30814 8419
rect 31196 0 31248 6645
rect 31276 0 31328 5791
rect 35398 0 35798 4764
rect 42203 0 42603 4764
rect 46673 0 46725 5791
rect 46753 0 46805 6645
rect 47187 0 47239 8419
rect 47267 0 47319 456
rect 47988 0 48040 5650
rect 48426 0 48478 9105
rect 48506 0 48558 5384
rect 49468 0 49520 1996
rect 49548 0 49600 1394
rect 49692 0 49761 417
rect 50834 0 50886 7338
rect 50914 0 50966 5790
rect 52324 0 52376 2035
rect 53658 0 53710 9204
rect 55931 0 55983 3493
rect 56607 0 56659 270
rect 60582 0 60752 4895
rect 60780 0 60949 5923
rect 80568 0 80620 4506
rect 80999 0 81051 2962
rect 83889 0 83941 885
rect 84538 0 84590 4506
rect 88968 0 89020 3359
rect 89581 0 89633 15042
rect 89731 0 89783 13125
rect 89881 0 89933 16725
rect 90031 0 90083 47202
rect 90181 0 90233 47266
rect 90331 0 90383 47330
rect 90481 0 90533 46836
rect 90631 0 90683 3086
rect 90781 0 90833 3210
rect 92906 0 93034 9087
rect 93206 0 93334 9805
<< obsm2 >>
rect 301 47386 95700 50680
rect 301 47322 90275 47386
rect 301 47258 90125 47322
rect 301 16781 89975 47258
rect 301 15098 89825 16781
rect 301 9260 89525 15098
rect 301 5979 24235 9260
rect 301 0 16996 5979
rect 17277 4951 24235 5979
rect 17475 3549 24235 4951
rect 17475 326 21962 3549
rect 17475 0 21286 326
rect 21450 0 21962 326
rect 22126 0 24235 3549
rect 24399 9161 53602 9260
rect 24399 7394 29467 9161
rect 24399 5846 27059 7394
rect 24399 2091 26979 5846
rect 24399 0 25569 2091
rect 25733 0 26979 2091
rect 27223 5440 29467 7394
rect 27223 2052 29387 5440
rect 27223 1450 28425 2052
rect 27223 473 28345 1450
rect 27223 0 28184 473
rect 28589 0 29387 2052
rect 29631 8475 48370 9161
rect 29631 7045 30706 8475
rect 29631 5706 30626 7045
rect 29631 0 29905 5706
rect 30069 536 30626 5706
rect 30069 512 30706 536
rect 30069 0 30626 512
rect 30870 6701 47131 8475
rect 30870 0 31140 6701
rect 31304 5847 46697 6701
rect 31384 4820 46617 5847
rect 31384 0 35342 4820
rect 35854 0 42147 4820
rect 42659 0 46617 4820
rect 46861 0 47131 6701
rect 47295 5706 48370 8475
rect 47295 512 47932 5706
rect 47375 0 47932 512
rect 48096 0 48370 5706
rect 48534 7394 53602 9161
rect 48534 5440 50778 7394
rect 48614 2052 50778 5440
rect 48614 0 49412 2052
rect 49576 1450 50778 2052
rect 49656 473 50778 1450
rect 49817 0 50778 473
rect 50942 5846 53602 7394
rect 51022 2091 53602 5846
rect 51022 0 52268 2091
rect 52432 0 53602 2091
rect 53766 5979 89525 9260
rect 53766 4951 60724 5979
rect 53766 3549 60526 4951
rect 53766 0 55875 3549
rect 56039 326 60526 3549
rect 56039 0 56551 326
rect 56715 0 60526 326
rect 61005 4562 89525 5979
rect 61005 0 80512 4562
rect 80676 3018 84482 4562
rect 80676 0 80943 3018
rect 81107 941 84482 3018
rect 81107 0 83833 941
rect 83997 0 84482 941
rect 84646 3415 89525 4562
rect 84646 0 88912 3415
rect 89076 0 89525 3415
rect 89689 13181 89825 15098
rect 90439 46892 95700 47386
rect 90589 9861 95700 46892
rect 90589 9143 93150 9861
rect 90589 3266 92850 9143
rect 90589 3142 90725 3266
rect 90889 0 92850 3266
rect 93090 0 93150 9143
rect 93390 0 95700 9861
<< obsm3 >>
rect 60 451 95940 50743
<< metal4 >>
rect 0 45900 254 50743
rect 95746 45900 96000 50743
rect 9867 45548 79857 45580
rect 9867 45480 9967 45548
rect 8963 44576 9867 45480
rect 8124 43737 8963 44576
rect 6941 42554 8124 43737
rect 5886 41499 6941 42554
rect 11602 40293 12210 40901
rect 11069 39790 11602 40293
rect 5852 39760 11602 39790
rect 77594 39853 78642 40901
rect 83642 40615 84822 41795
rect 10829 39550 11069 39760
rect 5852 39520 11069 39550
rect 5852 31877 10829 39520
rect 5150 31856 10829 31877
rect 78642 38503 79992 39853
rect 84822 39209 86228 40615
rect 79992 37333 81162 38503
rect 86228 38009 87428 39209
rect 81162 36133 82362 37333
rect 87428 37325 88112 38009
rect 82362 35263 83232 36133
rect 88800 35335 90102 36637
rect 84252 33493 85002 34243
rect 90102 34062 91375 35335
rect 85632 32173 86322 32863
rect 91375 32859 92578 34062
rect 92578 32178 93259 32859
rect 5150 31175 5852 31856
rect 4764 30789 5150 31175
rect 86802 30973 87522 31693
rect 93259 31490 93947 32178
rect 4080 30105 4764 30789
rect 87522 30343 88152 30973
rect 93947 30547 94890 31490
rect 0 24750 254 29743
rect 3718 29743 4080 30105
rect 88152 29610 88885 30343
rect 94890 29743 95694 30547
rect 95746 24750 96000 29743
rect 0 23560 254 24450
rect 95746 23560 96000 24450
rect 0 22390 254 23280
rect 95746 22390 96000 23280
rect 0 22024 1013 22090
rect 94927 22024 96000 22090
rect 0 21368 89769 21964
rect 89833 21368 96000 21964
rect 0 21072 254 21308
rect 95746 21072 96000 21308
rect 0 20416 89872 21012
rect 89936 20416 96000 21012
rect 0 20290 1013 20356
rect 94927 20290 96000 20356
rect 0 19060 254 19990
rect 95746 19060 96000 19990
rect 0 18090 254 18780
rect 95746 18090 96000 18780
rect 0 17120 254 17810
rect 95746 17120 96000 17810
rect 0 15910 254 16840
rect 95746 15910 96000 16840
rect 0 14700 254 15630
rect 1916 14691 1933 14700
rect 1916 14683 91585 14691
rect 95746 14700 96000 15630
rect 0 13730 193 14420
rect 95807 13730 96000 14420
rect 0 12520 254 13450
rect 95746 12520 96000 13450
rect 0 11150 254 12240
rect 95746 11150 96000 12240
<< obsm4 >>
rect 334 45820 95666 50743
rect 193 45660 95807 45820
rect 193 45560 9787 45660
rect 193 44656 8883 45560
rect 193 43817 8044 44656
rect 79937 45468 95807 45660
rect 10047 45400 95807 45468
rect 193 42634 6861 43817
rect 9947 44496 95807 45400
rect 193 41419 5806 42634
rect 9043 43657 95807 44496
rect 8204 42474 95807 43657
rect 7021 41875 95807 42474
rect 7021 41419 83562 41875
rect 193 40981 83562 41419
rect 193 40373 11522 40981
rect 193 39870 10989 40373
rect 193 39680 5772 39870
rect 12290 40213 77514 40981
rect 11682 39773 77514 40213
rect 78722 40535 83562 40981
rect 84902 40695 95807 41875
rect 78722 39933 84742 40535
rect 193 39630 10749 39680
rect 193 31957 5772 39630
rect 11682 39680 78562 39773
rect 193 31255 5070 31957
rect 11149 39440 78562 39680
rect 10909 38423 78562 39440
rect 80072 39129 84742 39933
rect 86308 39289 95807 40695
rect 80072 38583 86148 39129
rect 10909 37253 79912 38423
rect 81242 37929 86148 38583
rect 87508 38089 95807 39289
rect 81242 37413 87348 37929
rect 10909 36053 81082 37253
rect 82442 37245 87348 37413
rect 88192 37245 95807 38089
rect 82442 36717 95807 37245
rect 82442 36213 88720 36717
rect 10909 35183 82282 36053
rect 83312 35255 88720 36213
rect 90182 35415 95807 36717
rect 83312 35183 90022 35255
rect 10909 34323 90022 35183
rect 10909 33413 84172 34323
rect 85082 33982 90022 34323
rect 91455 34142 95807 35415
rect 85082 33413 91295 33982
rect 10909 32943 91295 33413
rect 10909 32093 85552 32943
rect 86402 32779 91295 32943
rect 92658 32939 95807 34142
rect 86402 32098 92498 32779
rect 93339 32258 95807 32939
rect 86402 32093 93179 32098
rect 193 30869 4684 31255
rect 10909 31776 93179 32093
rect 5932 31773 93179 31776
rect 193 30185 4000 30869
rect 5932 31095 86722 31773
rect 5230 30893 86722 31095
rect 87602 31410 93179 31773
rect 94027 31570 95807 32258
rect 87602 31053 93867 31410
rect 193 29823 3638 30185
rect 5230 30709 87442 30893
rect 4844 30263 87442 30709
rect 88232 30467 93867 31053
rect 94970 30627 95807 31570
rect 88232 30423 94810 30467
rect 334 29663 3638 29823
rect 4844 30025 88072 30263
rect 4160 29663 88072 30025
rect 334 29530 88072 29663
rect 88965 29663 94810 30423
rect 95774 29823 95807 30627
rect 88965 29530 95666 29663
rect 334 24670 95666 29530
rect 193 24530 95807 24670
rect 334 23480 95666 24530
rect 193 23360 95807 23480
rect 334 22310 95666 23360
rect 193 22170 95807 22310
rect 1093 22044 94847 22170
rect 334 21092 95666 21288
rect 1093 20210 94847 20336
rect 193 20070 95807 20210
rect 334 18980 95666 20070
rect 193 18860 95807 18980
rect 334 18010 95666 18860
rect 193 17890 95807 18010
rect 334 17040 95666 17890
rect 193 16920 95807 17040
rect 334 15830 95666 16920
rect 193 15710 95807 15830
rect 334 14780 95666 15710
rect 334 14620 1836 14780
rect 2013 14771 95666 14780
rect 193 14603 1836 14620
rect 91665 14620 95666 14771
rect 91665 14603 95807 14620
rect 193 14500 95807 14603
rect 273 13650 95727 14500
rect 193 13530 95807 13650
rect 334 12440 95666 13530
rect 193 12320 95807 12440
rect 334 11150 95666 12320
<< metal5 >>
rect 0 45900 254 50743
rect 95746 45900 96000 50743
rect 9891 45545 79857 45580
rect 9891 45504 9967 45545
rect 8987 44600 9891 45504
rect 8221 43834 8987 44600
rect 6965 42578 8221 43834
rect 5910 41523 6965 42578
rect 11578 40269 12207 40898
rect 11069 39840 11578 40269
rect 5852 39760 11578 39840
rect 10829 39600 11069 39760
rect 5852 39520 11069 39600
rect 77594 39871 78621 40898
rect 83618 40639 84798 41819
rect 5852 31877 10829 39520
rect 5337 31816 10829 31877
rect 5337 31362 5852 31816
rect 4788 30813 5337 31362
rect 4268 30293 4788 30813
rect 3718 29743 4268 30293
rect 0 24750 254 29740
rect 21438 26397 33978 38920
rect 44023 26397 56563 38920
rect 78621 38514 79978 39871
rect 79978 37314 81178 38514
rect 86204 38033 87404 39233
rect 81178 36153 82339 37314
rect 87404 37349 88088 38033
rect 88776 35359 90078 36661
rect 84218 33554 84938 34274
rect 90078 34086 91351 35359
rect 84938 32882 85610 33554
rect 85610 32194 86298 32882
rect 91351 32883 92554 34086
rect 86298 31704 86788 32194
rect 92554 32202 93235 32883
rect 86788 30966 87526 31704
rect 87526 30354 88138 30966
rect 88142 29740 88752 30350
rect 94866 29740 95697 30571
rect 95725 24750 96000 29740
rect 0 23580 254 24430
rect 0 22410 254 23260
rect 0 20290 254 22090
rect 0 19080 254 19970
rect 0 18111 254 18760
rect 95746 23580 96000 24430
rect 95746 22410 96000 23260
rect 95746 20290 96000 22090
rect 95746 19080 96000 19970
rect 95746 18111 96000 18760
rect 0 17140 254 17790
rect 0 15930 254 16820
rect 0 14720 254 15610
rect 95746 17140 96000 17790
rect 95746 15930 96000 16820
rect 95746 14720 96000 15610
rect 0 13750 193 14400
rect 95807 13750 96000 14400
rect 0 12540 254 13430
rect 0 11170 254 12220
rect 95746 12540 96000 13430
rect 95746 11170 96000 12220
<< obsm5 >>
rect 574 45900 95426 50743
rect 574 45824 9571 45900
rect 574 45580 8667 45824
rect 80177 45580 95426 45900
rect 0 44920 8667 45580
rect 0 44154 7901 44920
rect 80177 45225 96000 45580
rect 10287 45184 96000 45225
rect 0 42898 6645 44154
rect 10211 44280 96000 45184
rect 0 41203 5590 42898
rect 9307 43514 96000 44280
rect 8541 42258 96000 43514
rect 7285 42139 96000 42258
rect 7285 41218 83298 42139
rect 7285 41203 11258 41218
rect 0 40589 11258 41203
rect 0 40160 10749 40589
rect 0 32197 5532 40160
rect 12527 39949 77274 41218
rect 11898 39551 77274 39949
rect 78941 40319 83298 41218
rect 85118 40319 96000 42139
rect 78941 40191 96000 40319
rect 0 31682 5017 32197
rect 11898 39440 78301 39551
rect 11389 39240 78301 39440
rect 11389 39200 21118 39240
rect 0 31133 4468 31682
rect 11149 31496 21118 39200
rect 0 30613 3948 31133
rect 6172 31042 21118 31496
rect 0 30060 3398 30613
rect 5657 30493 21118 31042
rect 574 29743 3398 30060
rect 5108 29973 21118 30493
rect 4588 29743 21118 29973
rect 0 29740 21118 29743
rect 574 29423 3398 29740
rect 4588 29423 21118 29740
rect 574 26077 21118 29423
rect 34298 26077 43703 39240
rect 56883 38194 78301 39240
rect 80298 39553 96000 40191
rect 80298 38834 85884 39553
rect 56883 36994 79658 38194
rect 81498 37713 85884 38834
rect 87724 38353 96000 39553
rect 81498 37634 87084 37713
rect 56883 35833 80858 36994
rect 82659 37029 87084 37634
rect 88408 37029 96000 38353
rect 82659 36981 96000 37029
rect 82659 35833 88456 36981
rect 56883 35039 88456 35833
rect 90398 35679 96000 36981
rect 56883 34594 89758 35039
rect 56883 33234 83898 34594
rect 85258 33874 89758 34594
rect 91671 34406 96000 35679
rect 85930 33766 89758 33874
rect 56883 32562 84618 33234
rect 85930 33202 91031 33766
rect 56883 31874 85290 32562
rect 86618 32563 91031 33202
rect 92874 33203 96000 34406
rect 86618 32514 92234 32563
rect 56883 31384 85978 31874
rect 87108 32024 92234 32514
rect 87846 31882 92234 32024
rect 93555 31882 96000 33203
rect 56883 30646 86468 31384
rect 87846 31286 96000 31882
rect 56883 30034 87206 30646
rect 88458 30891 96000 31286
rect 88458 30670 94546 30891
rect 56883 29420 87822 30034
rect 89072 29420 94546 30670
rect 56883 26077 95405 29420
rect 574 24430 95405 26077
rect 574 18111 95426 24430
rect 0 18110 96000 18111
rect 574 14400 95426 18110
rect 513 13750 95487 14400
rect 574 11170 95426 13750
<< labels >>
rlabel metal5 s 95746 20290 96000 22090 6 vssa
port 1 nsew ground bidirectional
rlabel metal5 s 0 20290 254 22090 6 vssa
port 1 nsew ground bidirectional
rlabel metal5 s 0 18111 254 18760 6 vssa
port 1 nsew ground bidirectional
rlabel metal5 s 95746 18111 96000 18760 6 vssa
port 1 nsew ground bidirectional
rlabel metal4 s 94927 22024 96000 22090 6 vssa
port 1 nsew ground bidirectional
rlabel metal4 s 94927 20290 96000 20356 6 vssa
port 1 nsew ground bidirectional
rlabel metal4 s 95746 21072 96000 21308 6 vssa
port 1 nsew ground bidirectional
rlabel metal4 s 0 18090 254 18780 6 vssa
port 1 nsew ground bidirectional
rlabel metal4 s 0 22024 1013 22090 6 vssa
port 1 nsew ground bidirectional
rlabel metal4 s 0 20290 1013 20356 6 vssa
port 1 nsew ground bidirectional
rlabel metal4 s 95746 18090 96000 18780 6 vssa
port 1 nsew ground bidirectional
rlabel metal4 s 0 21072 254 21308 6 vssa
port 1 nsew ground bidirectional
rlabel metal5 s 95746 14720 96000 15610 6 vddio
port 2 nsew power bidirectional
rlabel metal5 s 95725 24750 96000 29740 6 vddio
port 2 nsew power bidirectional
rlabel metal5 s 0 14720 254 15610 6 vddio
port 2 nsew power bidirectional
rlabel metal5 s 0 24750 254 29740 6 vddio
port 2 nsew power bidirectional
rlabel metal4 s 95746 24750 96000 29743 6 vddio
port 2 nsew power bidirectional
rlabel metal4 s 95746 14700 96000 15630 6 vddio
port 2 nsew power bidirectional
rlabel metal4 s 0 24750 254 29743 6 vddio
port 2 nsew power bidirectional
rlabel metal4 s 0 14700 254 15630 6 vddio
port 2 nsew power bidirectional
rlabel metal5 s 88142 29740 88752 30350 6 vddio
port 2 nsew power bidirectional
rlabel metal5 s 94866 29740 95697 30571 6 vddio
port 2 nsew power bidirectional
rlabel metal5 s 87526 30354 88138 30966 6 vddio
port 2 nsew power bidirectional
rlabel metal5 s 86788 30966 87526 31704 6 vddio
port 2 nsew power bidirectional
rlabel metal5 s 86298 31704 86788 32194 6 vddio
port 2 nsew power bidirectional
rlabel metal5 s 92554 32202 93235 32883 6 vddio
port 2 nsew power bidirectional
rlabel metal5 s 85610 32194 86298 32882 6 vddio
port 2 nsew power bidirectional
rlabel metal5 s 84938 32882 85610 33554 6 vddio
port 2 nsew power bidirectional
rlabel metal5 s 91351 32883 92554 34086 6 vddio
port 2 nsew power bidirectional
rlabel metal5 s 84218 33554 84938 34274 6 vddio
port 2 nsew power bidirectional
rlabel metal5 s 90078 34086 91351 35359 6 vddio
port 2 nsew power bidirectional
rlabel metal5 s 88776 35359 90078 36661 6 vddio
port 2 nsew power bidirectional
rlabel metal5 s 81178 36153 82339 37314 6 vddio
port 2 nsew power bidirectional
rlabel metal5 s 87404 37349 88088 38033 6 vddio
port 2 nsew power bidirectional
rlabel metal5 s 79978 37314 81178 38514 6 vddio
port 2 nsew power bidirectional
rlabel metal5 s 86204 38033 87404 39233 6 vddio
port 2 nsew power bidirectional
rlabel metal5 s 78621 38514 79978 39871 6 vddio
port 2 nsew power bidirectional
rlabel metal5 s 77594 39871 78621 40898 6 vddio
port 2 nsew power bidirectional
rlabel metal5 s 9967 45545 79857 45580 6 vddio
port 2 nsew power bidirectional
rlabel metal5 s 9891 45504 9967 45580 6 vddio
port 2 nsew power bidirectional
rlabel metal5 s 8987 44600 9891 45504 6 vddio
port 2 nsew power bidirectional
rlabel metal5 s 8221 43834 8987 44600 6 vddio
port 2 nsew power bidirectional
rlabel metal5 s 6965 42578 8221 43834 6 vddio
port 2 nsew power bidirectional
rlabel metal5 s 5910 41523 6965 42578 6 vddio
port 2 nsew power bidirectional
rlabel metal5 s 83618 40639 84798 41819 6 vddio
port 2 nsew power bidirectional
rlabel metal5 s 11578 40269 12207 40898 6 vddio
port 2 nsew power bidirectional
rlabel metal5 s 11069 39760 11578 40269 6 vddio
port 2 nsew power bidirectional
rlabel metal5 s 5852 39760 11069 39840 6 vddio
port 2 nsew power bidirectional
rlabel metal5 s 10829 39520 11069 39760 6 vddio
port 2 nsew power bidirectional
rlabel metal5 s 5852 39520 10829 39600 6 vddio
port 2 nsew power bidirectional
rlabel metal5 s 5852 31877 10829 39520 6 vddio
port 2 nsew power bidirectional
rlabel metal5 s 5852 31816 10829 31877 6 vddio
port 2 nsew power bidirectional
rlabel metal5 s 5337 31362 5852 31877 6 vddio
port 2 nsew power bidirectional
rlabel metal5 s 4788 30813 5337 31362 6 vddio
port 2 nsew power bidirectional
rlabel metal5 s 4268 30293 4788 30813 6 vddio
port 2 nsew power bidirectional
rlabel metal5 s 3718 29743 4268 30293 6 vddio
port 2 nsew power bidirectional
rlabel metal4 s 1916 14683 1933 14700 6 vddio
port 2 nsew power bidirectional
rlabel metal4 s 1933 14683 91585 14691 6 vddio
port 2 nsew power bidirectional
rlabel metal4 s 3718 29743 4080 30105 6 vddio
port 2 nsew power bidirectional
rlabel metal4 s 88152 29610 88885 30343 6 vddio
port 2 nsew power bidirectional
rlabel metal4 s 94890 29743 95694 30547 6 vddio
port 2 nsew power bidirectional
rlabel metal4 s 87522 30343 88152 30973 6 vddio
port 2 nsew power bidirectional
rlabel metal4 s 93947 30547 94890 31490 6 vddio
port 2 nsew power bidirectional
rlabel metal4 s 86802 30973 87522 31693 6 vddio
port 2 nsew power bidirectional
rlabel metal4 s 93259 31490 93947 32178 6 vddio
port 2 nsew power bidirectional
rlabel metal4 s 92578 32178 93259 32859 6 vddio
port 2 nsew power bidirectional
rlabel metal4 s 85632 32173 86322 32863 6 vddio
port 2 nsew power bidirectional
rlabel metal4 s 91375 32859 92578 34062 6 vddio
port 2 nsew power bidirectional
rlabel metal4 s 84252 33493 85002 34243 6 vddio
port 2 nsew power bidirectional
rlabel metal4 s 90102 34062 91375 35335 6 vddio
port 2 nsew power bidirectional
rlabel metal4 s 82362 35263 83232 36133 6 vddio
port 2 nsew power bidirectional
rlabel metal4 s 88800 35335 90102 36637 6 vddio
port 2 nsew power bidirectional
rlabel metal4 s 81162 36133 82362 37333 6 vddio
port 2 nsew power bidirectional
rlabel metal4 s 87428 37325 88112 38009 6 vddio
port 2 nsew power bidirectional
rlabel metal4 s 79992 37333 81162 38503 6 vddio
port 2 nsew power bidirectional
rlabel metal4 s 86228 38009 87428 39209 6 vddio
port 2 nsew power bidirectional
rlabel metal4 s 78642 38503 79992 39853 6 vddio
port 2 nsew power bidirectional
rlabel metal4 s 84822 39209 86228 40615 6 vddio
port 2 nsew power bidirectional
rlabel metal4 s 77594 39853 78642 40901 6 vddio
port 2 nsew power bidirectional
rlabel metal4 s 4080 30105 4764 30789 6 vddio
port 2 nsew power bidirectional
rlabel metal4 s 4764 30789 5150 31175 6 vddio
port 2 nsew power bidirectional
rlabel metal4 s 5150 31175 5852 31877 6 vddio
port 2 nsew power bidirectional
rlabel metal4 s 5852 31856 10829 31877 6 vddio
port 2 nsew power bidirectional
rlabel metal4 s 5852 31877 10829 39520 6 vddio
port 2 nsew power bidirectional
rlabel metal4 s 11602 40293 12210 40901 6 vddio
port 2 nsew power bidirectional
rlabel metal4 s 11069 39760 11602 40293 6 vddio
port 2 nsew power bidirectional
rlabel metal4 s 5852 39760 11069 39790 6 vddio
port 2 nsew power bidirectional
rlabel metal4 s 10829 39520 11069 39760 6 vddio
port 2 nsew power bidirectional
rlabel metal4 s 5852 39520 10829 39550 6 vddio
port 2 nsew power bidirectional
rlabel metal4 s 83642 40615 84822 41795 6 vddio
port 2 nsew power bidirectional
rlabel metal4 s 5886 41499 6941 42554 6 vddio
port 2 nsew power bidirectional
rlabel metal4 s 6941 42554 8124 43737 6 vddio
port 2 nsew power bidirectional
rlabel metal4 s 8124 43737 8963 44576 6 vddio
port 2 nsew power bidirectional
rlabel metal4 s 8963 44576 9867 45480 6 vddio
port 2 nsew power bidirectional
rlabel metal4 s 9867 45480 9967 45580 6 vddio
port 2 nsew power bidirectional
rlabel metal4 s 9967 45548 79857 45580 6 vddio
port 2 nsew power bidirectional
rlabel metal5 s 95746 12540 96000 13430 6 vccd
port 3 nsew power bidirectional
rlabel metal5 s 0 12540 254 13430 6 vccd
port 3 nsew power bidirectional
rlabel metal4 s 95746 12520 96000 13450 6 vccd
port 3 nsew power bidirectional
rlabel metal4 s 0 12520 254 13450 6 vccd
port 3 nsew power bidirectional
rlabel metal5 s 95746 11170 96000 12220 6 vcchib
port 4 nsew power bidirectional
rlabel metal5 s 0 11170 254 12220 6 vcchib
port 4 nsew power bidirectional
rlabel metal4 s 95746 11150 96000 12240 6 vcchib
port 4 nsew power bidirectional
rlabel metal4 s 0 11150 254 12240 6 vcchib
port 4 nsew power bidirectional
rlabel metal5 s 95807 13750 96000 14400 6 vdda
port 5 nsew power bidirectional
rlabel metal5 s 0 13750 193 14400 6 vdda
port 5 nsew power bidirectional
rlabel metal4 s 95807 13730 96000 14420 6 vdda
port 5 nsew power bidirectional
rlabel metal4 s 0 13730 193 14420 6 vdda
port 5 nsew power bidirectional
rlabel metal5 s 95746 23580 96000 24430 6 vddio_q
port 6 nsew power bidirectional
rlabel metal5 s 0 23580 254 24430 6 vddio_q
port 6 nsew power bidirectional
rlabel metal4 s 95746 23560 96000 24450 6 vddio_q
port 6 nsew power bidirectional
rlabel metal4 s 0 23560 254 24450 6 vddio_q
port 6 nsew power bidirectional
rlabel metal5 s 0 19080 254 19970 6 vssd
port 7 nsew ground bidirectional
rlabel metal5 s 95746 19080 96000 19970 6 vssd
port 7 nsew ground bidirectional
rlabel metal4 s 95746 19060 96000 19990 6 vssd
port 7 nsew ground bidirectional
rlabel metal4 s 0 19060 254 19990 6 vssd
port 7 nsew ground bidirectional
rlabel metal5 s 0 15930 254 16820 6 vssio
port 8 nsew ground bidirectional
rlabel metal5 s 95746 45900 96000 50743 6 vssio
port 8 nsew ground bidirectional
rlabel metal5 s 0 45900 254 50743 6 vssio
port 8 nsew ground bidirectional
rlabel metal5 s 95746 15930 96000 16820 6 vssio
port 8 nsew ground bidirectional
rlabel metal4 s 95746 15910 96000 16840 6 vssio
port 8 nsew ground bidirectional
rlabel metal4 s 0 15910 254 16840 6 vssio
port 8 nsew ground bidirectional
rlabel metal4 s 95746 45900 96000 50743 6 vssio
port 8 nsew ground bidirectional
rlabel metal4 s 0 45900 254 50743 6 vssio
port 8 nsew ground bidirectional
rlabel metal5 s 0 17140 254 17790 6 vswitch
port 9 nsew power bidirectional
rlabel metal5 s 95746 17140 96000 17790 6 vswitch
port 9 nsew power bidirectional
rlabel metal4 s 95746 17120 96000 17810 6 vswitch
port 9 nsew power bidirectional
rlabel metal4 s 0 17120 254 17810 6 vswitch
port 9 nsew power bidirectional
rlabel metal5 s 0 22410 254 23260 6 vssio_q
port 10 nsew ground bidirectional
rlabel metal5 s 95746 22410 96000 23260 6 vssio_q
port 10 nsew ground bidirectional
rlabel metal4 s 95746 22390 96000 23280 6 vssio_q
port 10 nsew ground bidirectional
rlabel metal4 s 0 22390 254 23280 6 vssio_q
port 10 nsew ground bidirectional
rlabel metal5 s 44023 26397 56563 38920 6 pad<1>
port 11 nsew signal bidirectional
rlabel metal5 s 21438 26397 33978 38920 6 pad<0>
port 12 nsew signal bidirectional
rlabel metal4 s 89936 20416 96000 21012 6 amuxbus_b
port 13 nsew signal bidirectional
rlabel metal4 s 0 20416 89872 21012 6 amuxbus_b
port 13 nsew signal bidirectional
rlabel metal2 s 89731 0 89783 13125 6 amuxbus_b
port 13 nsew signal bidirectional
rlabel metal4 s 89833 21368 96000 21964 6 amuxbus_a
port 14 nsew signal bidirectional
rlabel metal4 s 0 21368 89769 21964 6 amuxbus_a
port 14 nsew signal bidirectional
rlabel metal2 s 89581 0 89633 15042 6 amuxbus_a
port 14 nsew signal bidirectional
rlabel metal2 s 88968 0 89020 3359 6 vreg_en_refgen
port 15 nsew signal input
rlabel metal2 s 80999 0 81051 2962 6 hld_h_n_refgen
port 16 nsew signal input
rlabel metal2 s 89881 0 89933 16725 6 voh_sel<0>
port 17 nsew signal input
rlabel metal2 s 90031 0 90083 47202 6 voh_sel<1>
port 18 nsew signal input
rlabel metal2 s 90181 0 90233 47266 6 voh_sel<2>
port 19 nsew signal input
rlabel metal2 s 83889 0 83941 885 6 vohref
port 20 nsew signal input
rlabel metal2 s 90481 0 90533 46836 6 enable_vdda_h
port 21 nsew signal input
rlabel metal2 s 80568 0 80620 4506 6 vtrip_sel_refgen
port 22 nsew signal input
rlabel metal2 s 90331 0 90383 47330 6 dft_refgen
port 23 nsew signal input
rlabel metal2 s 46753 0 46805 6645 6 dm1<1>
port 24 nsew signal input
rlabel metal2 s 47187 0 47239 8419 6 dm1<2>
port 25 nsew signal input
rlabel metal2 s 46673 0 46725 5791 6 dm1<0>
port 26 nsew signal input
rlabel metal2 s 31276 0 31328 5791 6 dm0<0>
port 27 nsew signal input
rlabel metal2 s 31196 0 31248 6645 6 dm0<1>
port 28 nsew signal input
rlabel metal2 s 30762 0 30814 8419 6 dm0<2>
port 29 nsew signal input
rlabel metal2 s 92906 0 93034 9087 6 voutref_dft
port 30 nsew signal bidirectional
rlabel metal2 s 84538 0 84590 4506 6 ibuf_sel_refgen
port 31 nsew signal input
rlabel metal2 s 90631 0 90683 3086 6 vref_sel<0>
port 32 nsew signal input
rlabel metal2 s 35398 0 35798 4764 6 pad_a_esd_1_h<0>
port 33 nsew signal bidirectional
rlabel metal2 s 50914 0 50966 5790 6 ibuf_sel<1>
port 34 nsew signal input
rlabel metal2 s 93206 0 93334 9805 6 vinref_dft
port 35 nsew signal bidirectional
rlabel metal2 s 42203 0 42603 4764 6 pad_a_esd_1_h<1>
port 36 nsew signal bidirectional
rlabel metal2 s 60780 0 60949 5923 6 pad_a_esd_0_h<1>
port 37 nsew signal bidirectional
rlabel metal2 s 90781 0 90833 3210 6 vref_sel<1>
port 38 nsew signal input
rlabel metal2 s 17052 0 17221 5923 6 pad_a_esd_0_h<0>
port 39 nsew signal bidirectional
rlabel metal2 s 17249 0 17419 4895 6 pad_a_noesd_h<0>
port 40 nsew signal bidirectional
rlabel metal2 s 60582 0 60752 4895 6 pad_a_noesd_h<1>
port 41 nsew signal bidirectional
rlabel metal2 s 56607 0 56659 270 6 inp_dis<1>
port 42 nsew signal input
rlabel metal2 s 21342 0 21394 270 6 inp_dis<0>
port 43 nsew signal input
rlabel metal2 s 22018 0 22070 3493 6 tie_lo_esd<0>
port 44 nsew signal output
rlabel metal2 s 55931 0 55983 3493 6 tie_lo_esd<1>
port 45 nsew signal output
rlabel metal2 s 53658 0 53710 9204 6 out<1>
port 46 nsew signal input
rlabel metal2 s 24291 0 24343 9204 6 out<0>
port 47 nsew signal input
rlabel metal2 s 25625 0 25677 2035 6 vtrip_sel<0>
port 48 nsew signal input
rlabel metal2 s 52324 0 52376 2035 6 vtrip_sel<1>
port 49 nsew signal input
rlabel metal2 s 47267 0 47319 456 6 enable_h
port 50 nsew signal input
rlabel metal2 s 30682 0 30734 456 6 enable_h
port 50 nsew signal input
rlabel metal2 s 30682 605 30734 6989 6 enable_h
port 50 nsew signal input
rlabel metal2 s 30682 592 30734 605 6 enable_h
port 50 nsew signal input
rlabel metal2 s 29961 0 30013 5650 6 vreg_en<0>
port 51 nsew signal input
rlabel metal2 s 47988 0 48040 5650 6 vreg_en<1>
port 52 nsew signal input
rlabel metal2 s 48426 0 48478 9105 6 slow<1>
port 53 nsew signal input
rlabel metal2 s 29523 0 29575 9105 6 slow<0>
port 54 nsew signal input
rlabel metal2 s 29443 0 29495 5384 6 oe_n<0>
port 55 nsew signal input
rlabel metal2 s 48506 0 48558 5384 6 oe_n<1>
port 56 nsew signal input
rlabel metal2 s 49468 0 49520 1996 6 in_h<1>
port 57 nsew signal output
rlabel metal2 s 28481 0 28533 1996 6 in_h<0>
port 58 nsew signal output
rlabel metal2 s 28401 0 28453 1394 6 in<0>
port 59 nsew signal output
rlabel metal2 s 49548 0 49600 1394 6 in<1>
port 60 nsew signal output
rlabel metal2 s 49692 0 49761 417 6 hld_ovr<1>
port 61 nsew signal input
rlabel metal2 s 28240 0 28309 417 6 hld_ovr<0>
port 62 nsew signal input
rlabel metal2 s 50834 0 50886 7338 6 hld_h_n<1>
port 63 nsew signal input
rlabel metal2 s 27115 0 27167 7338 6 hld_h_n<0>
port 64 nsew signal input
rlabel metal2 s 27035 0 27087 5790 6 ibuf_sel<0>
port 65 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 96000 50743
string LEFclass BLOCK
string LEFsymmetry R90
string LEFview TRUE
string GDS_END 112905430
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 102516404
<< end >>
