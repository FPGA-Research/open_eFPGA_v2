magic
tech sky130A
magscale 1 2
timestamp 1707688321
<< nwell >>
rect 8185 2284 8326 2401
rect 8158 2145 8326 2284
rect 8185 1812 8326 2145
rect 8185 1752 8304 1812
tri 8304 1790 8326 1812 nw
rect 8125 1615 8304 1752
rect 7879 1579 8304 1615
rect -177 -134 4673 854
rect 7273 -104 8167 202
<< pwell >>
rect -43 3935 2214 4021
rect 6185 3935 8452 4023
rect -43 1530 43 3935
rect 8364 2871 8452 3935
rect -43 1496 4911 1530
rect -43 1444 5509 1496
rect -43 937 43 1444
rect 4859 1415 5509 1444
rect 5165 1094 5509 1415
rect 6445 1481 7924 1496
rect 6445 1094 8157 1481
rect 6826 1060 8157 1094
rect 6962 1017 8157 1060
rect 6962 972 7184 1017
<< pdiff >>
rect 7104 5277 7116 5319
rect 7622 5277 7634 5319
rect 7104 4861 7116 4903
rect 7622 4861 7634 4903
rect 7369 590 7395 626
rect 8045 590 8071 626
rect 7369 492 7395 528
rect 8045 492 8071 528
<< psubdiff >>
rect 6211 3996 8426 3997
rect -17 3961 17 3995
rect 51 3961 85 3995
rect 119 3961 153 3995
rect 187 3961 221 3995
rect 255 3961 289 3995
rect 323 3961 357 3995
rect 391 3961 425 3995
rect 459 3961 493 3995
rect 527 3961 561 3995
rect 595 3961 629 3995
rect 663 3961 697 3995
rect 731 3961 765 3995
rect 799 3961 833 3995
rect 867 3961 901 3995
rect 935 3961 969 3995
rect 1003 3961 1037 3995
rect 1071 3961 1105 3995
rect 1139 3961 1173 3995
rect 1207 3961 1241 3995
rect 1275 3961 1309 3995
rect 1343 3961 1377 3995
rect 1411 3961 1445 3995
rect 1479 3961 1513 3995
rect 1547 3961 1581 3995
rect 1615 3961 1649 3995
rect 1683 3961 1717 3995
rect 1751 3961 1785 3995
rect 1819 3961 1853 3995
rect 1887 3961 1921 3995
rect 1955 3961 1989 3995
rect 2023 3961 2057 3995
rect 2091 3961 2188 3995
rect 6211 3962 6301 3996
rect 6335 3962 6369 3996
rect 6403 3962 6437 3996
rect 6471 3962 6505 3996
rect 6539 3962 6573 3996
rect 6607 3962 6641 3996
rect 6675 3962 6709 3996
rect 6743 3962 6777 3996
rect 6811 3962 6845 3996
rect 6879 3962 6913 3996
rect 6947 3962 6981 3996
rect 7015 3962 7049 3996
rect 7083 3962 7117 3996
rect 7151 3962 7185 3996
rect 7219 3962 7253 3996
rect 7287 3962 7321 3996
rect 7355 3962 7389 3996
rect 7423 3962 7457 3996
rect 7491 3962 7525 3996
rect 7559 3962 7593 3996
rect 7627 3962 7661 3996
rect 7695 3962 7729 3996
rect 7763 3962 7797 3996
rect 7831 3962 7865 3996
rect 7899 3962 7933 3996
rect 7967 3962 8001 3996
rect 8035 3962 8069 3996
rect 8103 3962 8137 3996
rect 8171 3962 8205 3996
rect 8239 3962 8307 3996
rect 8341 3962 8426 3996
rect 6211 3961 8426 3962
rect 8390 3934 8426 3961
rect -17 2737 17 2825
rect -17 2679 17 2703
rect -17 2483 17 2507
rect -17 2410 17 2449
rect -17 2337 17 2376
rect -17 2264 17 2303
rect -17 2191 17 2230
rect -17 2118 17 2157
rect -17 2045 17 2084
rect -17 1972 17 2011
rect -17 1899 17 1938
rect -17 1593 17 1865
rect -17 1522 17 1559
rect 17 1488 51 1504
rect -17 1470 51 1488
rect 85 1470 120 1504
rect 154 1470 189 1504
rect 223 1470 258 1504
rect 292 1470 327 1504
rect 361 1470 396 1504
rect 430 1470 465 1504
rect 499 1470 534 1504
rect 568 1470 603 1504
rect 637 1470 672 1504
rect 706 1470 741 1504
rect 775 1470 810 1504
rect 844 1470 879 1504
rect 913 1470 948 1504
rect 982 1470 1017 1504
rect 1051 1470 1086 1504
rect 1120 1470 1155 1504
rect 1189 1470 1224 1504
rect 1258 1470 1293 1504
rect 1327 1470 1362 1504
rect 1396 1470 1431 1504
rect 1465 1470 1500 1504
rect 1534 1470 1569 1504
rect 1603 1470 1638 1504
rect 1672 1470 1707 1504
rect 1741 1470 1776 1504
rect 1810 1470 1845 1504
rect 1879 1470 1914 1504
rect 1948 1470 1983 1504
rect 2017 1470 2052 1504
rect 2086 1470 2121 1504
rect 2155 1470 2190 1504
rect 2224 1470 2259 1504
rect 2293 1470 2328 1504
rect 2362 1470 2397 1504
rect 2431 1470 2466 1504
rect 2500 1470 2535 1504
rect 2569 1470 2604 1504
rect 2638 1470 2673 1504
rect 2707 1470 2742 1504
rect 2776 1470 2811 1504
rect 2845 1470 2880 1504
rect 2914 1470 2949 1504
rect 2983 1470 3018 1504
rect 3052 1470 3087 1504
rect 3121 1470 3155 1504
rect 3189 1470 3223 1504
rect 3257 1470 3291 1504
rect 3325 1470 3359 1504
rect 3393 1470 3427 1504
rect 3461 1470 3495 1504
rect 3529 1470 3563 1504
rect 3597 1470 3631 1504
rect 3665 1470 3699 1504
rect 3733 1470 3767 1504
rect 3801 1470 3835 1504
rect 3869 1470 3903 1504
rect 3937 1470 3971 1504
rect 4005 1470 4039 1504
rect 4073 1470 4107 1504
rect 4141 1470 4175 1504
rect 4209 1470 4243 1504
rect 4277 1470 4311 1504
rect 4345 1470 4379 1504
rect 4413 1470 4447 1504
rect 4481 1470 4515 1504
rect 4549 1470 4583 1504
rect 4617 1470 4651 1504
rect 4685 1470 4719 1504
rect 4753 1470 4787 1504
rect 4821 1470 4885 1504
rect -17 1451 17 1470
rect 4885 1441 4971 1470
rect 7084 1455 7898 1470
rect -17 1380 17 1417
rect 7084 1436 8131 1455
rect 7084 1402 7260 1436
rect 7294 1402 7333 1436
rect 7367 1402 7407 1436
rect 7441 1402 7481 1436
rect 7515 1402 7555 1436
rect 7589 1402 7629 1436
rect 7663 1402 7703 1436
rect 7737 1402 7777 1436
rect 7811 1402 7851 1436
rect 7885 1402 7925 1436
rect 7959 1402 7999 1436
rect 8033 1402 8073 1436
rect 8107 1402 8131 1436
rect -17 1322 17 1346
rect 5191 1231 5483 1387
rect 5191 1197 5236 1231
rect 5270 1197 5308 1231
rect 5342 1197 5380 1231
rect 5414 1197 5483 1231
rect 5191 1120 5483 1197
rect 6670 1266 6926 1388
rect 6670 1166 6753 1266
rect 6852 1166 6926 1266
rect 7084 1368 8131 1402
rect 7084 1334 7260 1368
rect 7294 1334 7333 1368
rect 7367 1334 7407 1368
rect 7441 1334 7481 1368
rect 7515 1334 7555 1368
rect 7589 1334 7629 1368
rect 7663 1334 7703 1368
rect 7737 1334 7777 1368
rect 7811 1334 7851 1368
rect 7885 1334 7925 1368
rect 7959 1334 7999 1368
rect 8033 1334 8073 1368
rect 8107 1334 8131 1368
rect 7084 1300 8131 1334
rect 7084 1266 7260 1300
rect 7294 1266 7333 1300
rect 7367 1266 7407 1300
rect 7441 1266 7481 1300
rect 7515 1266 7555 1300
rect 7589 1266 7629 1300
rect 7663 1266 7703 1300
rect 7737 1266 7777 1300
rect 7811 1266 7851 1300
rect 7885 1266 7925 1300
rect 7959 1266 7999 1300
rect 8033 1266 8073 1300
rect 8107 1266 8131 1300
rect 7084 1232 8131 1266
rect 7084 1198 7260 1232
rect 7294 1198 7333 1232
rect 7367 1198 7407 1232
rect 7441 1198 7481 1232
rect 7515 1198 7555 1232
rect 7589 1198 7629 1232
rect 7663 1198 7703 1232
rect 7737 1198 7777 1232
rect 7811 1198 7851 1232
rect 7885 1198 7925 1232
rect 7959 1198 7999 1232
rect 8033 1198 8073 1232
rect 8107 1198 8131 1232
rect 7084 1164 8131 1198
rect 7084 1130 7260 1164
rect 7294 1130 7333 1164
rect 7367 1130 7407 1164
rect 7441 1130 7481 1164
rect 7515 1130 7555 1164
rect 7589 1130 7629 1164
rect 7663 1130 7703 1164
rect 7737 1130 7777 1164
rect 7811 1130 7851 1164
rect 7885 1130 7925 1164
rect 7959 1130 7999 1164
rect 8033 1130 8073 1164
rect 8107 1130 8131 1164
rect 7084 1096 8131 1130
rect 7084 1062 7260 1096
rect 7294 1062 7333 1096
rect 7367 1062 7407 1096
rect 7441 1062 7481 1096
rect 7515 1062 7555 1096
rect 7589 1062 7629 1096
rect 7663 1062 7703 1096
rect 7737 1062 7777 1096
rect 7811 1062 7851 1096
rect 7885 1062 7925 1096
rect 7959 1062 7999 1096
rect 8033 1062 8073 1096
rect 8107 1062 8131 1096
rect 7084 1043 8131 1062
rect 7084 998 7158 1043
<< nsubdiff >>
rect 8203 2213 8283 2284
rect 8203 2179 8225 2213
rect 8259 2179 8283 2213
rect 8203 1833 8283 2179
rect 8125 1651 8159 1685
rect 8193 1651 8238 1685
rect 8097 106 8131 238
rect 7309 104 8131 106
rect 7309 70 7333 104
rect 7367 70 7407 104
rect 7441 70 7481 104
rect 7515 70 7555 104
rect 7589 70 7629 104
rect 7663 70 7703 104
rect 7737 70 7777 104
rect 7811 70 7851 104
rect 7885 70 7925 104
rect 7959 70 7999 104
rect 8033 70 8073 104
rect 8107 70 8131 104
rect 7309 36 8131 70
rect 7309 2 7333 36
rect 7367 2 7407 36
rect 7441 2 7481 36
rect 7515 2 7555 36
rect 7589 2 7629 36
rect 7663 2 7703 36
rect 7737 2 7777 36
rect 7811 2 7851 36
rect 7885 2 7925 36
rect 7959 2 7999 36
rect 8033 2 8073 36
rect 8107 2 8131 36
rect 7309 -32 8131 2
rect 7309 -66 7333 -32
rect 7367 -66 7407 -32
rect 7441 -66 7481 -32
rect 7515 -66 7555 -32
rect 7589 -66 7629 -32
rect 7663 -66 7703 -32
rect 7737 -66 7777 -32
rect 7811 -66 7851 -32
rect 7885 -66 7925 -32
rect 7959 -66 7999 -32
rect 8033 -66 8073 -32
rect 8107 -66 8131 -32
rect 7309 -68 8131 -66
<< mvpsubdiff >>
rect -17 3809 17 3833
rect -17 3738 17 3775
rect -17 3667 17 3704
rect -17 3596 17 3633
rect -17 3525 17 3562
rect -17 3454 17 3491
rect -17 3383 17 3420
rect -17 3312 17 3349
rect -17 3241 17 3278
rect -17 3170 17 3207
rect -17 3099 17 3136
rect -17 3027 17 3065
rect -17 2955 17 2993
rect -17 2897 17 2921
rect 8390 3772 8426 3806
rect 8390 3738 8391 3772
rect 8425 3738 8426 3772
rect 8390 3704 8426 3738
rect 8390 3670 8391 3704
rect 8425 3670 8426 3704
rect 8390 3636 8426 3670
rect 8390 3602 8391 3636
rect 8425 3602 8426 3636
rect 8390 3568 8426 3602
rect 8390 3534 8391 3568
rect 8425 3534 8426 3568
rect 8390 3500 8426 3534
rect 8390 3466 8391 3500
rect 8425 3466 8426 3500
rect 8390 3432 8426 3466
rect 8390 3398 8391 3432
rect 8425 3398 8426 3432
rect 8390 3364 8426 3398
rect 8390 3330 8391 3364
rect 8425 3330 8426 3364
rect 8390 3296 8426 3330
rect 8390 3262 8391 3296
rect 8425 3262 8426 3296
rect 8390 3228 8426 3262
rect 8390 3194 8391 3228
rect 8425 3194 8426 3228
rect 8390 3160 8426 3194
rect 8390 3126 8391 3160
rect 8425 3126 8426 3160
rect 8390 3092 8426 3126
rect 8390 3058 8391 3092
rect 8425 3058 8426 3092
rect 8390 3024 8426 3058
rect 8390 2990 8391 3024
rect 8425 2990 8426 3024
rect 8390 2897 8426 2990
rect -17 1226 17 1250
rect -17 1158 17 1192
rect -17 1090 17 1124
rect -17 1021 17 1056
rect -17 963 17 987
<< mvnsubdiff >>
rect -17 674 17 698
rect -17 603 17 640
rect -17 532 17 569
rect -17 461 17 498
rect -17 390 17 427
rect -17 319 17 356
rect -17 248 17 285
rect -17 177 17 214
rect -17 106 17 143
rect -17 34 17 72
rect -17 -34 17 0
rect 4571 72 4607 98
rect 4571 46 4572 72
rect 4606 46 4607 72
rect 4571 -34 4607 46
rect -17 -68 7 -34
rect 41 -68 76 -34
rect 110 -68 145 -34
rect 179 -68 214 -34
rect 248 -68 283 -34
rect 317 -68 352 -34
rect 386 -68 421 -34
rect 455 -68 490 -34
rect 524 -68 559 -34
rect 593 -68 628 -34
rect 662 -68 697 -34
rect 731 -68 766 -34
rect 800 -68 835 -34
rect 869 -68 904 -34
rect 938 -68 973 -34
rect 1007 -68 1042 -34
rect 1076 -68 1111 -34
rect 1145 -68 1180 -34
rect 1214 -68 1249 -34
rect 1283 -68 1318 -34
rect 1352 -68 1387 -34
rect 1421 -68 1456 -34
rect 1490 -68 1525 -34
rect 1559 -68 1594 -34
rect 1628 -68 1663 -34
rect 1697 -68 1732 -34
rect 1766 -68 1801 -34
rect 1835 -68 1870 -34
rect 1904 -68 1939 -34
rect 1973 -68 2008 -34
rect 2042 -68 2077 -34
rect 2111 -68 2146 -34
rect 2180 -68 2215 -34
rect 2249 -68 2284 -34
rect 2318 -68 2353 -34
rect 2387 -68 2422 -34
rect 2456 -68 2491 -34
rect 2525 -68 2560 -34
rect 2594 -68 2629 -34
rect 2663 -68 2698 -34
rect 2732 -68 2767 -34
rect 2801 -68 2836 -34
rect 2870 -68 2905 -34
rect 2939 -68 2974 -34
rect 3008 -68 3043 -34
rect 3077 -68 3112 -34
rect 3146 -68 3181 -34
rect 3215 -68 3250 -34
rect 3284 -68 3319 -34
rect 3353 -68 3388 -34
rect 3422 -68 3457 -34
rect 3491 -68 3526 -34
rect 3560 -68 3595 -34
rect 3629 -68 3664 -34
rect 3698 -68 3733 -34
rect 3767 -68 3801 -34
rect 3835 -68 3869 -34
rect 3903 -68 3937 -34
rect 3971 -68 4005 -34
rect 4039 -68 4073 -34
rect 4107 -68 4141 -34
rect 4175 -68 4209 -34
rect 4243 -68 4277 -34
rect 4311 -68 4345 -34
rect 4379 -68 4413 -34
rect 4447 -68 4481 -34
rect 4515 -68 4549 -34
rect 4583 -68 4607 -34
<< psubdiffcont >>
rect 17 3961 51 3995
rect 85 3961 119 3995
rect 153 3961 187 3995
rect 221 3961 255 3995
rect 289 3961 323 3995
rect 357 3961 391 3995
rect 425 3961 459 3995
rect 493 3961 527 3995
rect 561 3961 595 3995
rect 629 3961 663 3995
rect 697 3961 731 3995
rect 765 3961 799 3995
rect 833 3961 867 3995
rect 901 3961 935 3995
rect 969 3961 1003 3995
rect 1037 3961 1071 3995
rect 1105 3961 1139 3995
rect 1173 3961 1207 3995
rect 1241 3961 1275 3995
rect 1309 3961 1343 3995
rect 1377 3961 1411 3995
rect 1445 3961 1479 3995
rect 1513 3961 1547 3995
rect 1581 3961 1615 3995
rect 1649 3961 1683 3995
rect 1717 3961 1751 3995
rect 1785 3961 1819 3995
rect 1853 3961 1887 3995
rect 1921 3961 1955 3995
rect 1989 3961 2023 3995
rect 2057 3961 2091 3995
rect 6301 3962 6335 3996
rect 6369 3962 6403 3996
rect 6437 3962 6471 3996
rect 6505 3962 6539 3996
rect 6573 3962 6607 3996
rect 6641 3962 6675 3996
rect 6709 3962 6743 3996
rect 6777 3962 6811 3996
rect 6845 3962 6879 3996
rect 6913 3962 6947 3996
rect 6981 3962 7015 3996
rect 7049 3962 7083 3996
rect 7117 3962 7151 3996
rect 7185 3962 7219 3996
rect 7253 3962 7287 3996
rect 7321 3962 7355 3996
rect 7389 3962 7423 3996
rect 7457 3962 7491 3996
rect 7525 3962 7559 3996
rect 7593 3962 7627 3996
rect 7661 3962 7695 3996
rect 7729 3962 7763 3996
rect 7797 3962 7831 3996
rect 7865 3962 7899 3996
rect 7933 3962 7967 3996
rect 8001 3962 8035 3996
rect 8069 3962 8103 3996
rect 8137 3962 8171 3996
rect 8205 3962 8239 3996
rect 8307 3962 8341 3996
rect -17 2703 17 2737
rect -17 2449 17 2483
rect -17 2376 17 2410
rect -17 2303 17 2337
rect -17 2230 17 2264
rect -17 2157 17 2191
rect -17 2084 17 2118
rect -17 2011 17 2045
rect -17 1938 17 1972
rect -17 1865 17 1899
rect -17 1559 17 1593
rect -17 1488 17 1522
rect 51 1470 85 1504
rect 120 1470 154 1504
rect 189 1470 223 1504
rect 258 1470 292 1504
rect 327 1470 361 1504
rect 396 1470 430 1504
rect 465 1470 499 1504
rect 534 1470 568 1504
rect 603 1470 637 1504
rect 672 1470 706 1504
rect 741 1470 775 1504
rect 810 1470 844 1504
rect 879 1470 913 1504
rect 948 1470 982 1504
rect 1017 1470 1051 1504
rect 1086 1470 1120 1504
rect 1155 1470 1189 1504
rect 1224 1470 1258 1504
rect 1293 1470 1327 1504
rect 1362 1470 1396 1504
rect 1431 1470 1465 1504
rect 1500 1470 1534 1504
rect 1569 1470 1603 1504
rect 1638 1470 1672 1504
rect 1707 1470 1741 1504
rect 1776 1470 1810 1504
rect 1845 1470 1879 1504
rect 1914 1470 1948 1504
rect 1983 1470 2017 1504
rect 2052 1470 2086 1504
rect 2121 1470 2155 1504
rect 2190 1470 2224 1504
rect 2259 1470 2293 1504
rect 2328 1470 2362 1504
rect 2397 1470 2431 1504
rect 2466 1470 2500 1504
rect 2535 1470 2569 1504
rect 2604 1470 2638 1504
rect 2673 1470 2707 1504
rect 2742 1470 2776 1504
rect 2811 1470 2845 1504
rect 2880 1470 2914 1504
rect 2949 1470 2983 1504
rect 3018 1470 3052 1504
rect 3087 1470 3121 1504
rect 3155 1470 3189 1504
rect 3223 1470 3257 1504
rect 3291 1470 3325 1504
rect 3359 1470 3393 1504
rect 3427 1470 3461 1504
rect 3495 1470 3529 1504
rect 3563 1470 3597 1504
rect 3631 1470 3665 1504
rect 3699 1470 3733 1504
rect 3767 1470 3801 1504
rect 3835 1470 3869 1504
rect 3903 1470 3937 1504
rect 3971 1470 4005 1504
rect 4039 1470 4073 1504
rect 4107 1470 4141 1504
rect 4175 1470 4209 1504
rect 4243 1470 4277 1504
rect 4311 1470 4345 1504
rect 4379 1470 4413 1504
rect 4447 1470 4481 1504
rect 4515 1470 4549 1504
rect 4583 1470 4617 1504
rect 4651 1470 4685 1504
rect 4719 1470 4753 1504
rect 4787 1470 4821 1504
rect -17 1417 17 1451
rect 7260 1402 7294 1436
rect 7333 1402 7367 1436
rect 7407 1402 7441 1436
rect 7481 1402 7515 1436
rect 7555 1402 7589 1436
rect 7629 1402 7663 1436
rect 7703 1402 7737 1436
rect 7777 1402 7811 1436
rect 7851 1402 7885 1436
rect 7925 1402 7959 1436
rect 7999 1402 8033 1436
rect 8073 1402 8107 1436
rect -17 1346 17 1380
rect 5236 1197 5270 1231
rect 5308 1197 5342 1231
rect 5380 1197 5414 1231
rect 7260 1334 7294 1368
rect 7333 1334 7367 1368
rect 7407 1334 7441 1368
rect 7481 1334 7515 1368
rect 7555 1334 7589 1368
rect 7629 1334 7663 1368
rect 7703 1334 7737 1368
rect 7777 1334 7811 1368
rect 7851 1334 7885 1368
rect 7925 1334 7959 1368
rect 7999 1334 8033 1368
rect 8073 1334 8107 1368
rect 7260 1266 7294 1300
rect 7333 1266 7367 1300
rect 7407 1266 7441 1300
rect 7481 1266 7515 1300
rect 7555 1266 7589 1300
rect 7629 1266 7663 1300
rect 7703 1266 7737 1300
rect 7777 1266 7811 1300
rect 7851 1266 7885 1300
rect 7925 1266 7959 1300
rect 7999 1266 8033 1300
rect 8073 1266 8107 1300
rect 7260 1198 7294 1232
rect 7333 1198 7367 1232
rect 7407 1198 7441 1232
rect 7481 1198 7515 1232
rect 7555 1198 7589 1232
rect 7629 1198 7663 1232
rect 7703 1198 7737 1232
rect 7777 1198 7811 1232
rect 7851 1198 7885 1232
rect 7925 1198 7959 1232
rect 7999 1198 8033 1232
rect 8073 1198 8107 1232
rect 7260 1130 7294 1164
rect 7333 1130 7367 1164
rect 7407 1130 7441 1164
rect 7481 1130 7515 1164
rect 7555 1130 7589 1164
rect 7629 1130 7663 1164
rect 7703 1130 7737 1164
rect 7777 1130 7811 1164
rect 7851 1130 7885 1164
rect 7925 1130 7959 1164
rect 7999 1130 8033 1164
rect 8073 1130 8107 1164
rect 7260 1062 7294 1096
rect 7333 1062 7367 1096
rect 7407 1062 7441 1096
rect 7481 1062 7515 1096
rect 7555 1062 7589 1096
rect 7629 1062 7663 1096
rect 7703 1062 7737 1096
rect 7777 1062 7811 1096
rect 7851 1062 7885 1096
rect 7925 1062 7959 1096
rect 7999 1062 8033 1096
rect 8073 1062 8107 1096
<< nsubdiffcont >>
rect 8225 2179 8259 2213
rect 8159 1651 8193 1685
rect 7333 70 7367 104
rect 7407 70 7441 104
rect 7481 70 7515 104
rect 7555 70 7589 104
rect 7629 70 7663 104
rect 7703 70 7737 104
rect 7777 70 7811 104
rect 7851 70 7885 104
rect 7925 70 7959 104
rect 7999 70 8033 104
rect 8073 70 8107 104
rect 7333 2 7367 36
rect 7407 2 7441 36
rect 7481 2 7515 36
rect 7555 2 7589 36
rect 7629 2 7663 36
rect 7703 2 7737 36
rect 7777 2 7811 36
rect 7851 2 7885 36
rect 7925 2 7959 36
rect 7999 2 8033 36
rect 8073 2 8107 36
rect 7333 -66 7367 -32
rect 7407 -66 7441 -32
rect 7481 -66 7515 -32
rect 7555 -66 7589 -32
rect 7629 -66 7663 -32
rect 7703 -66 7737 -32
rect 7777 -66 7811 -32
rect 7851 -66 7885 -32
rect 7925 -66 7959 -32
rect 7999 -66 8033 -32
rect 8073 -66 8107 -32
<< mvpsubdiffcont >>
rect -17 3775 17 3809
rect -17 3704 17 3738
rect -17 3633 17 3667
rect -17 3562 17 3596
rect -17 3491 17 3525
rect -17 3420 17 3454
rect -17 3349 17 3383
rect -17 3278 17 3312
rect -17 3207 17 3241
rect -17 3136 17 3170
rect -17 3065 17 3099
rect -17 2993 17 3027
rect -17 2921 17 2955
rect 8391 3738 8425 3772
rect 8391 3670 8425 3704
rect 8391 3602 8425 3636
rect 8391 3534 8425 3568
rect 8391 3466 8425 3500
rect 8391 3398 8425 3432
rect 8391 3330 8425 3364
rect 8391 3262 8425 3296
rect 8391 3194 8425 3228
rect 8391 3126 8425 3160
rect 8391 3058 8425 3092
rect 8391 2990 8425 3024
rect -17 1192 17 1226
rect -17 1124 17 1158
rect -17 1056 17 1090
rect -17 987 17 1021
<< mvnsubdiffcont >>
rect -17 640 17 674
rect -17 569 17 603
rect -17 498 17 532
rect -17 427 17 461
rect -17 356 17 390
rect -17 285 17 319
rect -17 214 17 248
rect -17 143 17 177
rect 4572 114 4606 148
rect -17 72 17 106
rect -17 0 17 34
rect 4572 46 4606 72
rect 7 -68 41 -34
rect 76 -68 110 -34
rect 145 -68 179 -34
rect 214 -68 248 -34
rect 283 -68 317 -34
rect 352 -68 386 -34
rect 421 -68 455 -34
rect 490 -68 524 -34
rect 559 -68 593 -34
rect 628 -68 662 -34
rect 697 -68 731 -34
rect 766 -68 800 -34
rect 835 -68 869 -34
rect 904 -68 938 -34
rect 973 -68 1007 -34
rect 1042 -68 1076 -34
rect 1111 -68 1145 -34
rect 1180 -68 1214 -34
rect 1249 -68 1283 -34
rect 1318 -68 1352 -34
rect 1387 -68 1421 -34
rect 1456 -68 1490 -34
rect 1525 -68 1559 -34
rect 1594 -68 1628 -34
rect 1663 -68 1697 -34
rect 1732 -68 1766 -34
rect 1801 -68 1835 -34
rect 1870 -68 1904 -34
rect 1939 -68 1973 -34
rect 2008 -68 2042 -34
rect 2077 -68 2111 -34
rect 2146 -68 2180 -34
rect 2215 -68 2249 -34
rect 2284 -68 2318 -34
rect 2353 -68 2387 -34
rect 2422 -68 2456 -34
rect 2491 -68 2525 -34
rect 2560 -68 2594 -34
rect 2629 -68 2663 -34
rect 2698 -68 2732 -34
rect 2767 -68 2801 -34
rect 2836 -68 2870 -34
rect 2905 -68 2939 -34
rect 2974 -68 3008 -34
rect 3043 -68 3077 -34
rect 3112 -68 3146 -34
rect 3181 -68 3215 -34
rect 3250 -68 3284 -34
rect 3319 -68 3353 -34
rect 3388 -68 3422 -34
rect 3457 -68 3491 -34
rect 3526 -68 3560 -34
rect 3595 -68 3629 -34
rect 3664 -68 3698 -34
rect 3733 -68 3767 -34
rect 3801 -68 3835 -34
rect 3869 -68 3903 -34
rect 3937 -68 3971 -34
rect 4005 -68 4039 -34
rect 4073 -68 4107 -34
rect 4141 -68 4175 -34
rect 4209 -68 4243 -34
rect 4277 -68 4311 -34
rect 4345 -68 4379 -34
rect 4413 -68 4447 -34
rect 4481 -68 4515 -34
rect 4549 -68 4583 -34
<< locali >>
rect 6808 4609 6842 4647
rect 7114 4620 7162 4624
rect 7080 4552 7114 4590
rect 7610 4590 7642 4624
rect 7576 4552 7642 4590
rect 7610 4518 7642 4552
rect 6598 3997 7816 4032
rect 6068 3996 8426 3997
rect -17 3809 17 3995
rect 51 3961 85 3995
rect 119 3961 153 3995
rect 187 3961 221 3995
rect 255 3961 289 3995
rect 323 3961 357 3995
rect 391 3961 425 3995
rect 459 3961 493 3995
rect 527 3961 561 3995
rect 595 3961 629 3995
rect 663 3961 697 3995
rect 731 3961 765 3995
rect 799 3961 833 3995
rect 867 3961 901 3995
rect 935 3961 969 3995
rect 1003 3961 1037 3995
rect 1071 3961 1105 3995
rect 1139 3961 1173 3995
rect 1207 3961 1241 3995
rect 1275 3961 1309 3995
rect 1343 3961 1377 3995
rect 1411 3961 1445 3995
rect 1479 3961 1513 3995
rect 1547 3961 1581 3995
rect 1615 3961 1649 3995
rect 1683 3961 1717 3995
rect 1751 3961 1785 3995
rect 1819 3961 1853 3995
rect 1887 3961 1921 3995
rect 1955 3961 1989 3995
rect 2023 3961 2057 3995
rect 2091 3961 2188 3995
rect 6068 3962 6301 3996
rect 6335 3962 6369 3996
rect 6403 3962 6437 3996
rect 6471 3962 6505 3996
rect 6539 3962 6573 3996
rect 6607 3962 6641 3996
rect 6675 3962 6709 3996
rect 6743 3962 6777 3996
rect 6811 3962 6845 3996
rect 6879 3962 6913 3996
rect 6947 3962 6981 3996
rect 7015 3962 7049 3996
rect 7083 3962 7117 3996
rect 7151 3962 7185 3996
rect 7219 3962 7253 3996
rect 7287 3962 7321 3996
rect 7355 3962 7389 3996
rect 7423 3962 7457 3996
rect 7491 3962 7525 3996
rect 7559 3962 7593 3996
rect 7627 3962 7661 3996
rect 7695 3962 7729 3996
rect 7763 3962 7797 3996
rect 7831 3962 7865 3996
rect 7899 3962 7933 3996
rect 7967 3962 8001 3996
rect 8035 3962 8069 3996
rect 8103 3962 8137 3996
rect 8171 3962 8205 3996
rect 8239 3995 8307 3996
rect 8341 3995 8426 3996
rect 8270 3962 8307 3995
rect 6068 3961 8236 3962
rect 8270 3961 8308 3962
rect 8342 3961 8380 3995
rect 8414 3961 8426 3995
rect 6068 3960 8426 3961
rect 245 3877 283 3911
rect 435 3877 473 3911
rect 549 3861 1256 3911
rect -17 3738 17 3775
rect -17 3667 17 3704
rect -17 3596 17 3633
rect -17 3525 17 3561
rect -17 3454 17 3489
rect -17 3383 17 3420
rect 1150 3443 1256 3861
rect 1184 3409 1222 3443
rect 2948 3861 3655 3911
rect 3731 3877 3769 3911
rect 3921 3877 3959 3911
rect 4449 3877 4487 3911
rect 4639 3877 4677 3911
rect 4753 3861 5460 3911
rect 2948 3443 3054 3861
rect 2982 3409 3020 3443
rect 5354 3443 5460 3861
rect 5388 3409 5426 3443
rect 7152 3861 7859 3911
rect 7927 3877 7965 3911
rect 8125 3877 8163 3911
rect 7152 3443 7258 3861
rect 7186 3409 7224 3443
rect 8390 3772 8426 3960
rect 8390 3738 8391 3772
rect 8425 3738 8426 3772
rect 8390 3704 8426 3738
rect 8390 3670 8391 3704
rect 8425 3670 8426 3704
rect 8390 3636 8426 3670
rect 8390 3602 8391 3636
rect 8425 3602 8426 3636
rect 8390 3568 8426 3602
rect 8390 3534 8391 3568
rect 8425 3534 8426 3568
rect 8390 3500 8426 3534
rect 8390 3466 8391 3500
rect 8425 3466 8426 3500
rect 8390 3432 8426 3466
rect -17 3312 17 3349
rect -17 3241 17 3278
rect -17 3170 17 3207
rect -17 3099 17 3136
rect -17 3027 17 3065
rect -17 2955 17 2993
rect -17 2897 17 2921
rect 8390 3398 8391 3432
rect 8425 3398 8426 3432
rect 8390 3364 8426 3398
rect 8390 3330 8391 3364
rect 8425 3330 8426 3364
rect 8390 3296 8426 3330
rect 8390 3262 8391 3296
rect 8425 3262 8426 3296
rect 8390 3228 8426 3262
rect 8390 3194 8391 3228
rect 8425 3194 8426 3228
rect 8390 3160 8426 3194
rect 8390 3126 8391 3160
rect 8425 3126 8426 3160
rect 8390 3092 8426 3126
rect 8390 3058 8391 3092
rect 8425 3058 8426 3092
rect 8390 3024 8426 3058
rect 8390 2990 8391 3024
rect 8425 2990 8426 3024
rect 8390 2897 8426 2990
rect -17 2737 17 2825
rect -17 2679 17 2703
rect -17 2483 17 2507
rect -17 2410 17 2449
rect -17 2337 17 2376
rect -17 2264 17 2303
rect -17 2191 17 2230
rect -17 2118 17 2157
rect 8225 2264 8259 2284
rect 8225 2213 8259 2230
rect 8225 2145 8259 2158
rect -17 2045 17 2084
rect -17 1972 17 2011
rect -17 1899 17 1938
rect -17 1841 17 1865
rect 8125 1651 8159 1685
rect 8193 1651 8238 1685
rect -17 1593 17 1617
rect -17 1522 17 1559
rect 17 1488 51 1504
rect -17 1470 51 1488
rect 85 1470 120 1504
rect 154 1470 189 1504
rect 223 1470 258 1504
rect 292 1470 327 1504
rect 361 1470 396 1504
rect 430 1470 465 1504
rect 499 1470 534 1504
rect 568 1470 603 1504
rect 637 1470 672 1504
rect 706 1470 741 1504
rect 775 1470 810 1504
rect 844 1470 879 1504
rect 913 1470 948 1504
rect 982 1470 1017 1504
rect 1051 1470 1086 1504
rect 1120 1470 1155 1504
rect 1189 1470 1224 1504
rect 1258 1470 1293 1504
rect 1327 1470 1362 1504
rect 1396 1470 1431 1504
rect 1465 1470 1500 1504
rect 1534 1470 1569 1504
rect 1603 1470 1638 1504
rect 1672 1470 1707 1504
rect 1741 1470 1776 1504
rect 1810 1470 1845 1504
rect 1879 1470 1914 1504
rect 1948 1470 1983 1504
rect 2017 1470 2052 1504
rect 2086 1470 2121 1504
rect 2155 1470 2190 1504
rect 2224 1470 2259 1504
rect 2293 1470 2328 1504
rect 2362 1470 2397 1504
rect 2431 1470 2466 1504
rect 2500 1470 2535 1504
rect 2569 1470 2604 1504
rect 2638 1470 2673 1504
rect 2707 1470 2742 1504
rect 2776 1470 2811 1504
rect 2845 1470 2880 1504
rect 2914 1470 2949 1504
rect 2983 1470 3018 1504
rect 3052 1470 3087 1504
rect 3121 1470 3155 1504
rect 3189 1470 3223 1504
rect 3257 1470 3291 1504
rect 3325 1470 3359 1504
rect 3393 1470 3427 1504
rect 3461 1470 3495 1504
rect 3529 1470 3563 1504
rect 3597 1470 3631 1504
rect 3665 1470 3699 1504
rect 3733 1470 3767 1504
rect 3801 1470 3835 1504
rect 3869 1470 3903 1504
rect 3937 1470 3971 1504
rect 4005 1470 4039 1504
rect 4073 1470 4107 1504
rect 4141 1470 4175 1504
rect 4209 1470 4243 1504
rect 4277 1470 4311 1504
rect 4345 1470 4379 1504
rect 4413 1470 4447 1504
rect 4481 1470 4515 1504
rect 4549 1470 4583 1504
rect 4617 1470 4651 1504
rect 4685 1470 4719 1504
rect 4753 1470 4787 1504
rect 4821 1470 4885 1504
rect -17 1451 17 1470
rect -17 1380 17 1417
rect -17 1226 17 1346
rect 493 1332 505 1348
rect 187 1298 225 1332
rect 527 1298 565 1332
rect 493 1282 505 1298
rect -17 1158 17 1192
rect -17 1090 17 1124
rect -17 1021 17 1056
rect 4572 1250 5449 1470
rect -17 920 17 958
rect 275 920 309 958
rect 913 920 947 958
rect 1617 920 1651 958
rect 4433 920 4467 958
rect 4572 946 4759 1250
rect 5201 1231 5449 1250
rect 5201 1197 5236 1231
rect 5270 1197 5308 1231
rect 5342 1197 5380 1231
rect 5414 1197 5449 1231
rect 5201 1120 5449 1197
rect 6472 1455 7935 1470
rect 6472 1449 8131 1455
rect 6472 1436 8097 1449
rect 6472 1402 7260 1436
rect 7294 1402 7333 1436
rect 7367 1402 7407 1436
rect 7441 1402 7481 1436
rect 7515 1402 7555 1436
rect 7589 1402 7629 1436
rect 7663 1402 7703 1436
rect 7737 1402 7777 1436
rect 7811 1402 7851 1436
rect 7885 1402 7925 1436
rect 7959 1402 7999 1436
rect 8033 1402 8073 1436
rect 8107 1402 8131 1415
rect 6472 1377 8131 1402
rect 6472 1368 8097 1377
rect 6472 1334 7260 1368
rect 7294 1334 7333 1368
rect 7367 1334 7407 1368
rect 7441 1334 7481 1368
rect 7515 1334 7555 1368
rect 7589 1334 7629 1368
rect 7663 1334 7703 1368
rect 7737 1334 7777 1368
rect 7811 1334 7851 1368
rect 7885 1334 7925 1368
rect 7959 1334 7999 1368
rect 8033 1334 8073 1368
rect 8107 1334 8131 1343
rect 6472 1305 8131 1334
rect 6472 1300 8097 1305
rect 6472 1266 7260 1300
rect 7294 1266 7333 1300
rect 7367 1266 7407 1300
rect 7441 1266 7481 1300
rect 7515 1266 7555 1300
rect 7589 1266 7629 1300
rect 7663 1266 7703 1300
rect 7737 1266 7777 1300
rect 7811 1266 7851 1300
rect 7885 1266 7925 1300
rect 7959 1266 7999 1300
rect 8033 1266 8073 1300
rect 8107 1266 8131 1271
rect 6472 1120 6745 1266
rect 6852 1233 8131 1266
rect 6852 1232 8097 1233
rect 6852 1198 7260 1232
rect 7294 1198 7333 1232
rect 7367 1198 7407 1232
rect 7441 1198 7481 1232
rect 7515 1198 7555 1232
rect 7589 1198 7629 1232
rect 7663 1198 7703 1232
rect 7737 1198 7777 1232
rect 7811 1198 7851 1232
rect 7885 1198 7925 1232
rect 7959 1198 7999 1232
rect 8033 1198 8073 1232
rect 8107 1198 8131 1199
rect 6852 1164 8131 1198
rect 6852 1130 7260 1164
rect 7294 1130 7333 1164
rect 7367 1130 7407 1164
rect 7441 1130 7481 1164
rect 7515 1130 7555 1164
rect 7589 1130 7629 1164
rect 7663 1130 7703 1164
rect 7737 1130 7777 1164
rect 7811 1130 7851 1164
rect 7885 1130 7925 1164
rect 7959 1130 7999 1164
rect 8033 1130 8073 1164
rect 8107 1161 8131 1164
rect 6852 1127 8097 1130
rect 6852 1096 8131 1127
rect 6852 1086 7260 1096
rect 6988 1062 7260 1086
rect 7294 1062 7333 1096
rect 7367 1062 7407 1096
rect 7441 1062 7481 1096
rect 7515 1062 7555 1096
rect 7589 1062 7629 1096
rect 7663 1062 7703 1096
rect 7737 1062 7777 1096
rect 7811 1062 7851 1096
rect 7885 1062 7925 1096
rect 7959 1062 7999 1096
rect 8033 1062 8073 1096
rect 8107 1089 8131 1096
rect 6988 1055 8097 1062
rect 6988 1043 8131 1055
rect 6988 998 7037 1043
rect 275 770 309 808
rect 913 770 947 808
rect 1265 770 1299 808
rect 1617 770 1651 808
rect 1969 770 2003 808
rect 2321 770 2355 808
rect 2673 770 2707 808
rect 3025 770 3059 808
rect 3377 770 3411 808
rect 4081 770 4115 808
rect 4433 770 4467 808
rect 4572 770 4606 808
rect -17 674 17 698
rect -17 603 17 640
rect -17 532 17 569
rect -17 461 17 498
rect 7333 442 7367 476
rect -17 390 17 427
rect -17 319 17 356
rect -17 248 17 285
rect 5109 228 6837 272
rect -17 177 17 214
rect -17 106 17 143
rect 7309 106 7343 240
rect 8097 106 8131 238
rect 7309 104 8131 106
rect -17 34 17 72
rect -17 -34 17 0
rect 4572 72 4606 100
rect 4572 -34 4606 46
rect 7309 70 7333 104
rect 7367 70 7407 104
rect 7441 70 7481 104
rect 7515 70 7555 104
rect 7589 70 7629 104
rect 7663 70 7703 104
rect 7737 70 7777 104
rect 7811 70 7851 104
rect 7885 70 7925 104
rect 7959 70 7999 104
rect 8033 70 8073 104
rect 8107 70 8131 104
rect 7309 36 8131 70
rect 7309 2 7333 36
rect 7367 2 7407 36
rect 7441 2 7481 36
rect 7515 2 7555 36
rect 7589 2 7629 36
rect 7663 2 7703 36
rect 7737 2 7777 36
rect 7811 2 7851 36
rect 7885 2 7925 36
rect 7959 2 7999 36
rect 8033 2 8073 36
rect 8107 2 8131 36
rect 7309 -32 8131 2
rect -17 -68 7 -34
rect 41 -68 76 -34
rect 110 -68 145 -34
rect 179 -68 214 -34
rect 248 -68 283 -34
rect 317 -68 352 -34
rect 386 -68 421 -34
rect 455 -68 490 -34
rect 524 -68 559 -34
rect 593 -68 628 -34
rect 662 -68 697 -34
rect 731 -68 766 -34
rect 800 -68 835 -34
rect 869 -68 904 -34
rect 938 -68 973 -34
rect 1007 -68 1042 -34
rect 1076 -68 1111 -34
rect 1145 -68 1180 -34
rect 1214 -68 1249 -34
rect 1283 -68 1318 -34
rect 1352 -68 1387 -34
rect 1421 -68 1456 -34
rect 1490 -68 1525 -34
rect 1559 -68 1594 -34
rect 1628 -68 1663 -34
rect 1697 -68 1732 -34
rect 1766 -68 1801 -34
rect 1835 -68 1870 -34
rect 1904 -68 1939 -34
rect 1973 -68 2008 -34
rect 2042 -68 2077 -34
rect 2111 -68 2146 -34
rect 2180 -68 2215 -34
rect 2249 -68 2284 -34
rect 2318 -68 2353 -34
rect 2387 -68 2422 -34
rect 2456 -68 2491 -34
rect 2525 -68 2560 -34
rect 2594 -68 2629 -34
rect 2663 -68 2698 -34
rect 2732 -68 2767 -34
rect 2801 -68 2836 -34
rect 2870 -68 2905 -34
rect 2939 -68 2974 -34
rect 3008 -68 3043 -34
rect 3077 -68 3112 -34
rect 3146 -68 3181 -34
rect 3215 -68 3250 -34
rect 3284 -68 3319 -34
rect 3353 -68 3388 -34
rect 3422 -68 3457 -34
rect 3491 -68 3526 -34
rect 3560 -68 3595 -34
rect 3629 -68 3664 -34
rect 3698 -68 3733 -34
rect 3767 -68 3801 -34
rect 3835 -68 3869 -34
rect 3903 -68 3937 -34
rect 3971 -68 4005 -34
rect 4039 -68 4073 -34
rect 4107 -68 4141 -34
rect 4175 -68 4209 -34
rect 4243 -68 4277 -34
rect 4311 -68 4345 -34
rect 4379 -68 4413 -34
rect 4447 -68 4481 -34
rect 4515 -68 4549 -34
rect 4583 -68 4607 -34
rect 7309 -66 7333 -32
rect 7367 -66 7407 -32
rect 7441 -66 7481 -32
rect 7515 -66 7555 -32
rect 7589 -66 7629 -32
rect 7663 -66 7703 -32
rect 7737 -66 7777 -32
rect 7811 -66 7851 -32
rect 7885 -66 7925 -32
rect 7959 -66 7999 -32
rect 8033 -66 8073 -32
rect 8107 -66 8131 -32
rect 7309 -68 8131 -66
<< viali >>
rect 6808 4647 6842 4681
rect 6808 4575 6842 4609
rect 7080 4590 7114 4624
rect 7080 4518 7114 4552
rect 7576 4590 7610 4624
rect 7576 4518 7610 4552
rect 8236 3962 8239 3995
rect 8239 3962 8270 3995
rect 8308 3962 8341 3995
rect 8341 3962 8342 3995
rect 8236 3961 8270 3962
rect 8308 3961 8342 3962
rect 8380 3961 8414 3995
rect 211 3877 245 3911
rect 283 3877 317 3911
rect 401 3877 435 3911
rect 473 3877 507 3911
rect -17 3562 17 3595
rect -17 3561 17 3562
rect -17 3491 17 3523
rect -17 3489 17 3491
rect 1150 3409 1184 3443
rect 1222 3409 1256 3443
rect 3697 3877 3731 3911
rect 3769 3877 3803 3911
rect 3887 3877 3921 3911
rect 3959 3877 3993 3911
rect 4415 3877 4449 3911
rect 4487 3877 4521 3911
rect 4605 3877 4639 3911
rect 4677 3877 4711 3911
rect 2948 3409 2982 3443
rect 3020 3409 3054 3443
rect 5354 3409 5388 3443
rect 5426 3409 5460 3443
rect 7893 3877 7927 3911
rect 7965 3877 7999 3911
rect 8091 3877 8125 3911
rect 8163 3877 8197 3911
rect 7152 3409 7186 3443
rect 7224 3409 7258 3443
rect 8225 2230 8259 2264
rect 8225 2179 8259 2192
rect 8225 2158 8259 2179
rect 153 1298 187 1332
rect 225 1298 259 1332
rect 493 1298 527 1332
rect 565 1298 599 1332
rect -17 987 17 992
rect -17 958 17 987
rect -17 886 17 920
rect 275 958 309 992
rect 275 886 309 920
rect 913 958 947 992
rect 913 886 947 920
rect 1617 958 1651 992
rect 1617 886 1651 920
rect 4433 958 4467 992
rect 8097 1436 8131 1449
rect 8097 1415 8107 1436
rect 8107 1415 8131 1436
rect 8097 1368 8131 1377
rect 8097 1343 8107 1368
rect 8107 1343 8131 1368
rect 8097 1300 8131 1305
rect 8097 1271 8107 1300
rect 8107 1271 8131 1300
rect 8097 1232 8131 1233
rect 8097 1199 8107 1232
rect 8107 1199 8131 1232
rect 8097 1130 8107 1161
rect 8107 1130 8131 1161
rect 8097 1127 8131 1130
rect 8097 1062 8107 1089
rect 8107 1062 8131 1089
rect 8097 1055 8131 1062
rect 4433 886 4467 920
rect 275 808 309 842
rect 275 736 309 770
rect 913 808 947 842
rect 913 736 947 770
rect 1265 808 1299 842
rect 1265 736 1299 770
rect 1617 808 1651 842
rect 1617 736 1651 770
rect 1969 808 2003 842
rect 1969 736 2003 770
rect 2321 808 2355 842
rect 2321 736 2355 770
rect 2673 808 2707 842
rect 2673 736 2707 770
rect 3025 808 3059 842
rect 3025 736 3059 770
rect 3377 808 3411 842
rect 3377 736 3411 770
rect 4081 808 4115 842
rect 4081 736 4115 770
rect 4433 808 4467 842
rect 4433 736 4467 770
rect 4572 808 4606 842
rect 4572 736 4606 770
<< metal1 >>
tri 7307 5593 7383 5669 se
rect 7383 5663 7435 5669
rect 7383 5599 7435 5611
tri 6477 5541 6529 5593 se
rect 6529 5547 7383 5593
rect 6529 5541 7435 5547
tri 7765 5541 7819 5595 se
rect 7819 5589 7871 5595
tri 6455 5519 6477 5541 se
rect 6477 5519 6529 5541
tri 6529 5519 6551 5541 nw
tri 7743 5519 7765 5541 se
rect 7765 5537 7819 5541
rect 7765 5525 7871 5537
rect 7765 5519 7819 5525
tri 6449 5513 6455 5519 se
rect 6455 5513 6523 5519
tri 6523 5513 6529 5519 nw
tri 7737 5513 7743 5519 se
rect 7743 5513 7819 5519
tri 6404 5468 6449 5513 se
rect 6449 5479 6489 5513
tri 6489 5479 6523 5513 nw
tri 6529 5479 6563 5513 se
rect 6563 5479 7819 5513
rect 6449 5468 6478 5479
tri 6478 5468 6489 5479 nw
tri 6518 5468 6529 5479 se
rect 6529 5473 7819 5479
rect 6529 5468 7871 5473
rect 6091 5467 6477 5468
tri 6477 5467 6478 5468 nw
tri 6517 5467 6518 5468 se
rect 6518 5467 7871 5468
rect 6091 5447 6457 5467
tri 6457 5447 6477 5467 nw
tri 6497 5447 6517 5467 se
rect 6517 5447 6563 5467
tri 6563 5447 6583 5467 nw
rect 6091 5428 6438 5447
tri 6438 5428 6457 5447 nw
tri 6478 5428 6497 5447 se
rect 6091 5416 6426 5428
tri 6426 5416 6438 5428 nw
tri 6466 5416 6478 5428 se
rect 6478 5416 6497 5428
tri 6431 5381 6466 5416 se
rect 6466 5381 6497 5416
tri 6497 5381 6563 5447 nw
tri 6402 5352 6431 5381 se
rect 6431 5352 6468 5381
tri 6468 5352 6497 5381 nw
tri 6167 5232 6243 5308 se
rect 6243 5302 6295 5308
rect 6243 5238 6295 5250
rect 6094 5186 6243 5232
rect 6094 5180 6295 5186
tri 6352 5180 6402 5230 se
rect 6402 5210 6448 5352
tri 6448 5332 6468 5352 nw
tri 6336 5164 6352 5180 se
rect 6352 5164 6402 5180
tri 6402 5164 6448 5210 nw
tri 6270 5098 6336 5164 se
tri 6336 5098 6402 5164 nw
tri 6259 5087 6270 5098 se
rect 6270 5087 6325 5098
tri 6325 5087 6336 5098 nw
tri 6244 5072 6259 5087 se
rect 6259 5072 6310 5087
tri 6310 5072 6325 5087 nw
rect 6094 5026 6264 5072
tri 6264 5026 6310 5072 nw
rect 6050 4917 6094 4988
tri 6094 4917 6165 4988 sw
rect 7778 4945 8068 5235
tri 8402 5072 8417 5087 se
rect 8417 5072 8423 5087
tri 8356 5026 8402 5072 se
rect 8402 5035 8423 5072
rect 8475 5035 8481 5087
rect 8402 5026 8481 5035
tri 8318 4988 8356 5026 se
rect 8356 5023 8481 5026
rect 8356 4988 8423 5023
tri 8275 4945 8318 4988 se
rect 8318 4971 8423 4988
rect 8475 4971 8481 5023
rect 8318 4959 8481 4971
rect 8318 4945 8423 4959
tri 8247 4917 8275 4945 se
rect 8275 4917 8423 4945
rect 6050 4715 6904 4917
rect 7778 4907 8423 4917
rect 8475 4907 8481 4959
rect 7778 4895 8481 4907
rect 7778 4843 8423 4895
rect 8475 4843 8481 4895
rect 7778 4831 8481 4843
rect 7778 4779 8423 4831
rect 8475 4779 8481 4831
rect 7778 4767 8481 4779
rect 7778 4715 8423 4767
rect 8475 4715 8481 4767
rect 6050 4687 6137 4715
tri 6137 4687 6165 4715 nw
rect 6050 4681 6131 4687
tri 6131 4681 6137 4687 nw
rect 6050 4647 6097 4681
tri 6097 4647 6131 4681 nw
rect 6050 4641 6091 4647
tri 6091 4641 6097 4647 nw
rect 6793 4635 6799 4687
rect 6851 4635 6857 4687
rect 6793 4623 6857 4635
rect 6793 4571 6799 4623
rect 6851 4571 6857 4623
rect 6793 4569 6857 4571
rect 7071 4630 7123 4636
rect 7071 4566 7123 4578
rect 7071 4506 7123 4514
rect 7463 4630 7616 4636
rect 7515 4624 7616 4630
rect 7515 4590 7576 4624
rect 7610 4590 7616 4624
rect 7515 4578 7616 4590
rect 7463 4566 7616 4578
rect 7515 4552 7616 4566
rect 7515 4518 7576 4552
rect 7610 4518 7616 4552
rect 7515 4514 7616 4518
rect 7463 4506 7616 4514
tri 8146 4471 8156 4481 se
tri 7038 4465 7044 4471 se
rect 6094 4419 6584 4465
rect 7044 4419 7050 4471
rect 7102 4419 7114 4471
rect 7166 4419 7172 4471
tri 7172 4465 7178 4471 sw
tri 8140 4465 8146 4471 se
rect 8146 4465 8156 4471
rect 7827 4419 8156 4465
rect 6094 4391 8156 4419
rect 6094 4189 6599 4391
rect 7233 4211 7239 4391
rect 7355 4211 7361 4391
rect 7827 4189 8156 4391
rect 6094 4161 8156 4189
rect 6094 4109 6587 4161
rect 7044 4109 7050 4161
rect 7102 4109 7114 4161
rect 7166 4109 7172 4161
rect 7827 4109 8156 4161
rect 6094 4029 8563 4081
rect 7807 3957 8229 4001
rect 7807 3955 7952 3957
tri 7952 3955 7954 3957 nw
tri 8215 3955 8217 3957 ne
rect 8217 3955 8229 3957
rect 6094 3949 6415 3955
tri 6415 3949 6421 3955 nw
tri 8217 3949 8223 3955 ne
rect 8223 3949 8229 3955
rect 8281 3949 8293 4001
rect 8345 3995 8426 4001
rect 8345 3961 8380 3995
rect 8414 3961 8426 3995
rect 8345 3949 8426 3961
rect 8033 3923 8203 3929
rect 7594 3917 8005 3923
rect 199 3865 207 3917
rect 259 3865 271 3917
rect 323 3865 329 3917
rect 389 3911 456 3917
rect 389 3877 401 3911
rect 435 3877 456 3911
rect 389 3865 456 3877
rect 508 3865 520 3917
rect 572 3865 578 3917
rect 3626 3865 3632 3917
rect 3684 3865 3696 3917
rect 3748 3911 3815 3917
rect 3748 3877 3769 3911
rect 3803 3877 3815 3911
rect 3748 3865 3815 3877
rect 3875 3865 3881 3917
rect 3933 3865 3945 3917
rect 3997 3865 4005 3917
rect 4403 3865 4411 3917
rect 4463 3865 4475 3917
rect 4527 3865 4533 3917
rect 4593 3911 4660 3917
rect 4593 3877 4605 3911
rect 4639 3877 4660 3911
rect 4593 3865 4660 3877
rect 4712 3865 4724 3917
rect 4776 3865 4782 3917
rect 7594 3865 7600 3917
rect 7652 3865 7664 3917
rect 7716 3911 8005 3917
rect 7716 3877 7893 3911
rect 7927 3877 7965 3911
rect 7999 3877 8005 3911
rect 7716 3865 8005 3877
rect 8085 3911 8097 3923
rect 8149 3911 8203 3923
rect 8085 3877 8091 3911
rect 8149 3877 8163 3911
rect 8197 3877 8203 3911
rect 8085 3871 8097 3877
rect 8149 3871 8203 3877
rect 8033 3865 8203 3871
tri 8403 3865 8417 3879 se
tri 8375 3837 8403 3865 se
rect 8403 3837 8417 3865
rect -23 3606 23 3607
rect -23 3600 30 3606
rect -23 3548 -22 3600
rect -23 3536 30 3548
rect -23 3484 -22 3536
rect -23 3477 30 3484
rect 2143 3600 2345 3607
rect 2143 3548 2149 3600
rect 2201 3548 2218 3600
rect 2270 3548 2287 3600
rect 2339 3548 2345 3600
rect 2143 3536 2345 3548
rect 2143 3484 2149 3536
rect 2201 3484 2218 3536
rect 2270 3484 2287 3536
rect 2339 3484 2345 3536
rect 2143 3477 2345 3484
rect 4031 3600 4233 3607
rect 4031 3548 4037 3600
rect 4089 3548 4106 3600
rect 4158 3548 4175 3600
rect 4227 3548 4233 3600
rect 4031 3536 4233 3548
rect 4031 3484 4037 3536
rect 4089 3484 4106 3536
rect 4158 3484 4175 3536
rect 4227 3484 4233 3536
rect 4031 3477 4233 3484
rect 5177 3600 5543 3607
rect 5177 3548 5183 3600
rect 5235 3548 5259 3600
rect 5311 3548 5335 3600
rect 5387 3548 5410 3600
rect 5462 3548 5485 3600
rect 5537 3548 5543 3600
rect 5177 3536 5543 3548
rect 5177 3484 5183 3536
rect 5235 3484 5259 3536
rect 5311 3484 5335 3536
rect 5387 3484 5410 3536
rect 5462 3484 5485 3536
rect 5537 3484 5543 3536
rect 5177 3477 5543 3484
rect 5974 3599 6090 3605
rect 5974 3477 6090 3483
rect 6152 3600 6413 3607
rect 6152 3548 6158 3600
rect 6210 3548 6224 3600
rect 6276 3548 6290 3600
rect 6342 3548 6355 3600
rect 6407 3548 6413 3600
rect 6152 3536 6413 3548
rect 6152 3484 6158 3536
rect 6210 3484 6224 3536
rect 6276 3484 6290 3536
rect 6342 3484 6355 3536
rect 6407 3484 6413 3536
rect 6152 3477 6413 3484
rect 7200 3600 7387 3607
rect 7200 3548 7206 3600
rect 7258 3548 7329 3600
rect 7381 3548 7387 3600
rect 7200 3536 7387 3548
rect 7200 3484 7206 3536
rect 7258 3484 7329 3536
rect 7381 3484 7387 3536
rect 8152 3491 8158 3607
rect 8338 3491 8344 3607
rect 7200 3477 7387 3484
rect 1138 3443 3506 3449
rect 1138 3409 1150 3443
rect 1184 3409 1222 3443
rect 1256 3409 2948 3443
rect 2982 3409 3020 3443
rect 3054 3409 3506 3443
rect 1138 3397 3506 3409
rect 3558 3397 3570 3449
rect 3622 3443 7270 3449
rect 3622 3409 5354 3443
rect 5388 3409 5426 3443
rect 5460 3409 7152 3443
rect 7186 3409 7224 3443
rect 7258 3409 7270 3443
rect 3622 3397 7270 3409
rect 7670 3443 7722 3449
rect 7670 3379 7722 3391
tri 7645 3351 7670 3376 se
rect 59 3345 136 3351
rect 138 3350 174 3351
rect 111 3299 136 3345
rect 137 3300 175 3350
rect 176 3345 278 3351
rect 138 3299 174 3300
rect 176 3299 201 3345
rect 59 3281 111 3293
tri 111 3274 136 3299 nw
tri 176 3274 201 3299 ne
rect 253 3299 278 3345
rect 279 3300 280 3350
rect 316 3300 317 3350
rect 318 3299 426 3351
rect 428 3350 464 3351
rect 427 3300 465 3350
rect 466 3345 568 3351
rect 428 3299 464 3300
rect 466 3299 491 3345
rect 201 3281 253 3293
rect 59 3223 111 3229
tri 253 3274 278 3299 nw
tri 318 3274 343 3299 ne
rect 343 3268 401 3299
tri 401 3274 426 3299 nw
tri 466 3274 491 3299 ne
rect 543 3299 568 3345
rect 569 3300 570 3350
rect 606 3300 607 3350
rect 608 3344 3596 3351
rect 608 3299 855 3344
rect 491 3281 543 3293
rect 201 3223 253 3229
tri 543 3274 568 3299 nw
tri 830 3274 855 3299 ne
rect 907 3299 3596 3344
rect 3597 3300 3598 3350
rect 3634 3300 3635 3350
rect 3636 3345 3738 3351
rect 3740 3350 3776 3351
rect 3636 3299 3661 3345
rect 855 3280 907 3292
rect 491 3223 543 3229
tri 907 3274 932 3299 nw
tri 3636 3274 3661 3299 ne
rect 3713 3299 3738 3345
rect 3739 3300 3777 3350
rect 3740 3299 3776 3300
rect 3778 3299 3886 3351
rect 3887 3300 3888 3350
rect 3924 3300 3925 3350
rect 3926 3345 4028 3351
rect 4030 3350 4066 3351
rect 3926 3299 3951 3345
rect 3661 3281 3713 3293
rect 855 3222 907 3228
rect 1700 3264 1752 3270
rect 2373 3264 2425 3270
rect 1700 3200 1752 3212
tri 1752 3199 1777 3224 nw
tri 3713 3274 3738 3299 nw
tri 3778 3274 3803 3299 ne
rect 3803 3268 3861 3299
tri 3861 3274 3886 3299 nw
tri 3926 3274 3951 3299 ne
rect 4003 3299 4028 3345
rect 4029 3300 4067 3350
rect 4068 3345 4340 3351
rect 4342 3350 4378 3351
rect 4030 3299 4066 3300
rect 4068 3299 4262 3345
rect 3951 3281 4003 3293
rect 2425 3223 2449 3224
tri 2449 3223 2450 3224 nw
rect 3661 3223 3713 3229
tri 4003 3274 4028 3299 nw
tri 4237 3274 4262 3299 ne
rect 4314 3299 4340 3345
rect 4341 3300 4379 3350
rect 4380 3345 4482 3351
rect 4342 3299 4378 3300
rect 4380 3299 4405 3345
rect 4262 3281 4314 3293
rect 3951 3223 4003 3229
tri 4314 3274 4339 3299 nw
tri 4380 3274 4405 3299 ne
rect 4457 3299 4482 3345
rect 4483 3300 4484 3350
rect 4520 3300 4521 3350
rect 4522 3299 4630 3351
rect 4632 3350 4668 3351
rect 4631 3300 4669 3350
rect 4670 3345 4772 3351
rect 4632 3299 4668 3300
rect 4670 3299 4695 3345
rect 4405 3281 4457 3293
rect 4262 3223 4314 3229
tri 4457 3274 4482 3299 nw
tri 4522 3274 4547 3299 ne
rect 4547 3268 4605 3299
tri 4605 3274 4630 3299 nw
tri 4670 3274 4695 3299 ne
rect 4747 3299 4772 3345
rect 4773 3300 4774 3350
rect 4810 3300 4811 3350
rect 4812 3345 7605 3351
rect 4812 3299 5059 3345
rect 4695 3281 4747 3293
rect 4405 3223 4457 3229
tri 4747 3274 4772 3299 nw
tri 5034 3274 5059 3299 ne
rect 5111 3299 7605 3345
rect 7606 3300 7607 3350
rect 7643 3300 7644 3350
rect 7645 3327 7670 3351
rect 8007 3443 8258 3449
rect 8260 3448 8296 3449
rect 8059 3391 8071 3443
rect 8123 3391 8258 3443
rect 8007 3385 8258 3391
rect 8259 3386 8297 3448
rect 8298 3443 8375 3449
rect 8298 3391 8323 3443
rect 8260 3385 8296 3386
rect 8298 3385 8375 3391
tri 7722 3351 7747 3376 sw
rect 7722 3327 7749 3351
rect 7751 3350 7787 3351
rect 7645 3299 7749 3327
rect 7750 3300 7788 3350
rect 7789 3349 7855 3351
tri 7855 3349 7857 3351 sw
rect 7789 3337 7857 3349
tri 7857 3337 7869 3349 sw
rect 8007 3339 8065 3385
tri 8065 3360 8090 3385 nw
tri 8298 3360 8323 3385 ne
rect 8323 3379 8375 3385
rect 8008 3337 8064 3338
rect 7789 3321 7869 3337
tri 7869 3321 7885 3337 sw
rect 8323 3321 8375 3327
rect 7789 3301 7885 3321
tri 7885 3301 7905 3321 sw
rect 7751 3299 7787 3300
rect 7789 3299 7905 3301
tri 7905 3299 7907 3301 sw
rect 8008 3300 8064 3301
rect 5059 3281 5111 3293
rect 4695 3223 4747 3229
tri 5111 3274 5136 3299 nw
tri 7832 3274 7857 3299 ne
rect 7857 3274 7907 3299
tri 7907 3274 7932 3299 sw
tri 7982 3274 8007 3299 se
rect 8007 3274 8065 3299
tri 7857 3270 7861 3274 ne
rect 7861 3270 8065 3274
rect 5059 3223 5111 3229
rect 5884 3264 5936 3270
rect 2373 3200 2425 3212
rect 1700 3142 1752 3148
tri 2425 3199 2449 3223 nw
rect 6676 3264 6728 3270
rect 5884 3200 5936 3212
rect 2373 3142 2425 3148
tri 5936 3199 5961 3224 nw
tri 6651 3199 6676 3224 ne
tri 7861 3247 7884 3270 ne
rect 7884 3247 8065 3270
tri 7884 3222 7909 3247 ne
rect 7909 3222 8007 3247
rect 6676 3200 6728 3212
rect 5884 3142 5936 3148
tri 7982 3197 8007 3222 ne
rect 6676 3142 6728 3148
rect 59 2952 111 2958
rect 4029 2952 4081 2958
tri 57 2888 59 2890 se
rect 59 2888 111 2900
tri 111 2888 136 2913 sw
rect 4262 2952 4314 2958
rect 4029 2889 4081 2900
tri 4081 2889 4105 2913 sw
rect 8233 2927 8525 2933
rect 4029 2888 4105 2889
tri 4105 2888 4106 2889 sw
tri 4261 2888 4262 2889 se
rect 4262 2888 4314 2900
tri 4314 2888 4339 2913 sw
rect 59 2830 111 2836
rect 4029 2830 4081 2836
rect 8233 2883 8473 2927
tri 8351 2858 8376 2883 nw
tri 8448 2858 8473 2883 ne
rect 8473 2863 8525 2875
rect 4262 2830 4314 2836
rect 8473 2805 8525 2811
rect -161 2486 34 2688
rect 3806 2678 3922 2684
rect 3806 2492 3922 2498
rect 4114 2676 4230 2682
rect 7228 2497 7234 2677
rect 7350 2497 7356 2677
rect 4114 2490 4230 2496
rect 1990 2452 4466 2458
rect 1990 2412 4414 2452
tri 4072 2387 4097 2412 nw
tri 4304 2387 4329 2412 ne
rect 4329 2400 4414 2412
rect 6194 2412 6484 2458
rect 4329 2388 4466 2400
rect 4329 2336 4414 2388
tri 4466 2387 4491 2412 nw
rect 4329 2330 4466 2336
rect 8219 2264 8482 2276
rect 8219 2230 8225 2264
rect 8259 2230 8482 2264
rect 8219 2192 8482 2230
rect 8219 2158 8225 2192
rect 8259 2158 8482 2192
rect 8219 2146 8482 2158
tri 8420 2118 8448 2146 ne
rect 185 1841 219 2043
rect 6836 1863 6842 2043
rect 6958 1863 6964 2043
tri 8420 1813 8448 1841 se
rect 8448 1813 8482 2146
rect 0 1695 34 1813
rect 8437 1695 8482 1813
rect -29 1615 3564 1667
rect 3616 1615 3628 1667
rect 3680 1615 7965 1667
rect -29 1535 4428 1587
rect 4480 1535 4492 1587
rect 4544 1535 7897 1587
rect 7949 1535 7961 1587
rect 8013 1535 8019 1587
rect -17 1455 1530 1507
rect 1582 1455 1594 1507
rect 1646 1455 2558 1507
rect 2610 1455 2622 1507
rect 2674 1455 5734 1507
rect 5786 1455 5798 1507
rect 5850 1455 8255 1507
tri 8043 1449 8049 1455 ne
rect 8049 1449 8255 1455
tri 8049 1415 8083 1449 ne
rect 8083 1415 8097 1449
rect 8131 1415 8255 1449
tri 8083 1407 8091 1415 ne
rect 8091 1377 8255 1415
rect 139 1286 145 1338
rect 197 1286 209 1338
rect 261 1286 271 1338
rect 481 1292 488 1344
rect 540 1292 552 1344
rect 604 1292 611 1344
rect 8091 1343 8097 1377
rect 8131 1343 8255 1377
rect 8091 1305 8255 1343
rect 8091 1271 8097 1305
rect 8131 1271 8255 1305
rect 8091 1233 8255 1271
rect -161 1026 116 1228
rect 3806 1221 3922 1227
rect 3806 1035 3922 1041
rect 4115 1221 4231 1227
rect 4115 1035 4231 1041
rect 7231 1037 7237 1217
rect 7353 1037 7359 1217
rect 8091 1199 8097 1233
rect 8131 1199 8255 1233
rect 8091 1161 8255 1199
rect 8091 1127 8097 1161
rect 8131 1127 8255 1161
rect 8091 1089 8255 1127
rect 8091 1055 8097 1089
rect 8131 1055 8255 1089
rect 8091 1043 8255 1055
tri 8091 1037 8097 1043 ne
rect 8097 1037 8139 1043
tri 8097 1035 8099 1037 ne
rect 8099 1035 8139 1037
tri 8099 1026 8108 1035 ne
rect 8108 1026 8139 1035
tri 8108 998 8136 1026 ne
rect 8136 998 8139 1026
rect -29 992 116 998
rect -29 958 -17 992
rect 17 958 116 992
rect -29 952 116 958
rect 263 992 321 998
rect 263 958 275 992
rect 309 958 321 992
tri -54 927 -29 952 ne
rect -29 920 29 952
tri 29 927 54 952 nw
tri 238 927 263 952 ne
rect -29 886 -17 920
rect 17 886 29 920
rect -29 880 29 886
rect 263 920 321 958
rect 901 992 959 998
rect 901 958 913 992
rect 947 958 959 992
tri 321 927 346 952 nw
tri 876 927 901 952 ne
rect 263 886 275 920
rect 309 886 321 920
rect 263 880 321 886
rect 901 920 959 958
rect 1605 992 1663 998
rect 1605 958 1617 992
rect 1651 958 1663 992
tri 959 927 984 952 nw
tri 1580 927 1605 952 ne
rect 901 886 913 920
rect 947 886 959 920
rect 901 880 959 886
rect 1605 920 1663 958
rect 4421 992 4479 998
tri 8136 995 8139 998 ne
rect 4421 958 4433 992
rect 4467 958 4479 992
rect 4421 952 4479 958
tri 1663 927 1688 952 nw
tri 4396 927 4421 952 ne
rect 4421 944 4496 952
tri 4496 944 4504 952 nw
rect 1605 886 1617 920
rect 1651 886 1663 920
rect 1605 880 1663 886
tri 3597 853 3622 878 ne
rect 3622 872 3628 924
rect 3680 872 3686 924
rect 4421 920 4479 944
tri 4479 927 4496 944 nw
rect 7885 938 8019 946
rect 4421 886 4433 920
rect 4467 886 4479 920
rect 4421 880 4479 886
rect 7885 886 7967 938
rect 3622 860 3686 872
rect 263 842 321 848
rect 263 808 275 842
rect 309 808 321 842
tri 238 776 263 801 se
rect -285 500 116 776
rect 263 770 321 808
rect 901 842 959 848
rect 901 808 913 842
rect 947 808 959 842
tri 321 776 346 801 sw
tri 876 776 901 801 se
rect 263 736 275 770
rect 309 736 321 770
rect 263 730 321 736
rect 901 770 959 808
rect 1253 842 1311 848
rect 1253 808 1265 842
rect 1299 808 1311 842
tri 959 776 984 801 sw
tri 1228 776 1253 801 se
rect 901 736 913 770
rect 947 736 959 770
rect 901 730 959 736
rect 1253 770 1311 808
rect 1605 842 1663 848
rect 1605 808 1617 842
rect 1651 808 1663 842
tri 1311 776 1336 801 sw
tri 1580 776 1605 801 se
rect 1253 736 1265 770
rect 1299 736 1311 770
rect 1253 730 1311 736
rect 1605 770 1663 808
rect 1957 842 2015 848
rect 1957 808 1969 842
rect 2003 808 2015 842
tri 1663 776 1688 801 sw
tri 1932 776 1957 801 se
rect 1605 736 1617 770
rect 1651 736 1663 770
rect 1605 730 1663 736
rect 1957 770 2015 808
rect 2309 842 2367 848
rect 2309 808 2321 842
rect 2355 808 2367 842
tri 2015 776 2040 801 sw
tri 2284 776 2309 801 se
rect 1957 736 1969 770
rect 2003 736 2015 770
rect 1957 730 2015 736
rect 2309 770 2367 808
rect 2661 842 2719 848
rect 2661 808 2673 842
rect 2707 808 2719 842
tri 2367 776 2392 801 sw
tri 2636 776 2661 801 se
rect 2309 736 2321 770
rect 2355 736 2367 770
rect 2309 730 2367 736
rect 2661 770 2719 808
rect 3013 842 3071 848
rect 3013 808 3025 842
rect 3059 808 3071 842
tri 2719 776 2744 801 sw
tri 2988 776 3013 801 se
rect 2661 736 2673 770
rect 2707 736 2719 770
rect 2661 730 2719 736
rect 3013 770 3071 808
rect 3365 842 3423 848
rect 3365 808 3377 842
rect 3411 808 3423 842
rect 3622 808 3628 860
rect 3680 808 3686 860
tri 3686 853 3711 878 nw
rect 7885 874 8019 886
rect 4069 842 4127 848
rect 4069 808 4081 842
rect 4115 808 4127 842
tri 3071 776 3096 801 sw
tri 3340 776 3365 801 se
rect 3013 736 3025 770
rect 3059 736 3071 770
rect 3013 730 3071 736
rect 3365 770 3423 808
tri 3423 776 3448 801 sw
tri 4044 776 4069 801 se
rect 3365 736 3377 770
rect 3411 736 3423 770
rect 3365 730 3423 736
rect 4069 770 4127 808
rect 4421 842 4618 848
rect 4421 808 4433 842
rect 4467 808 4572 842
rect 4606 808 4618 842
rect 7885 822 7967 874
rect 7885 816 8019 822
tri 4127 776 4152 801 sw
tri 4396 776 4421 801 se
rect 4421 776 4618 808
rect 4069 736 4081 770
rect 4115 736 4127 770
rect 4069 730 4127 736
rect 4421 770 4479 776
rect 4421 736 4433 770
rect 4467 736 4479 770
rect 4421 730 4479 736
rect 4560 770 4618 776
rect 4560 736 4572 770
rect 4606 736 4618 770
rect 4560 730 4618 736
tri 8114 625 8139 650 se
rect -285 -2 -23 500
rect 23 498 171 500
tri 171 498 173 500 nw
rect 23 444 117 498
tri 117 444 171 498 nw
tri 4620 444 4674 498 se
rect 4674 444 5089 545
tri 23 350 117 444 nw
rect 3290 330 5089 444
rect 6836 365 6842 545
rect 6958 365 6964 545
rect 3290 264 5056 330
tri 5056 264 5122 330 nw
tri 6838 278 6844 284 se
tri 6844 207 6869 232 nw
rect 8323 126 8375 132
tri 8298 56 8323 81 se
rect 8323 62 8375 74
rect 139 4 145 56
rect 197 4 209 56
rect 261 4 785 56
rect 837 4 849 56
rect 901 4 4348 56
rect 4400 4 4412 56
rect 4464 4 4989 56
rect 5041 4 5053 56
rect 5105 46 6956 56
tri 6956 46 6966 56 sw
tri 7184 46 7194 56 se
rect 7194 46 8323 56
rect 5105 10 8323 46
rect 5105 4 8375 10
rect -285 -74 23 -2
tri 23 -28 48 -3 sw
<< rmetal1 >>
rect 136 3350 138 3351
rect 174 3350 176 3351
rect 136 3300 137 3350
rect 175 3300 176 3350
rect 278 3350 280 3351
rect 136 3299 138 3300
rect 174 3299 176 3300
rect 278 3300 279 3350
rect 278 3299 280 3300
rect 316 3350 318 3351
rect 317 3300 318 3350
rect 316 3299 318 3300
rect 426 3350 428 3351
rect 464 3350 466 3351
rect 426 3300 427 3350
rect 465 3300 466 3350
rect 568 3350 570 3351
rect 426 3299 428 3300
rect 464 3299 466 3300
rect 568 3300 569 3350
rect 568 3299 570 3300
rect 606 3350 608 3351
rect 607 3300 608 3350
rect 3596 3350 3598 3351
rect 606 3299 608 3300
rect 3596 3300 3597 3350
rect 3596 3299 3598 3300
rect 3634 3350 3636 3351
rect 3635 3300 3636 3350
rect 3738 3350 3740 3351
rect 3776 3350 3778 3351
rect 3634 3299 3636 3300
rect 3738 3300 3739 3350
rect 3777 3300 3778 3350
rect 3738 3299 3740 3300
rect 3776 3299 3778 3300
rect 3886 3350 3888 3351
rect 3886 3300 3887 3350
rect 3886 3299 3888 3300
rect 3924 3350 3926 3351
rect 3925 3300 3926 3350
rect 4028 3350 4030 3351
rect 4066 3350 4068 3351
rect 3924 3299 3926 3300
rect 4028 3300 4029 3350
rect 4067 3300 4068 3350
rect 4340 3350 4342 3351
rect 4378 3350 4380 3351
rect 4028 3299 4030 3300
rect 4066 3299 4068 3300
rect 4340 3300 4341 3350
rect 4379 3300 4380 3350
rect 4482 3350 4484 3351
rect 4340 3299 4342 3300
rect 4378 3299 4380 3300
rect 4482 3300 4483 3350
rect 4482 3299 4484 3300
rect 4520 3350 4522 3351
rect 4521 3300 4522 3350
rect 4520 3299 4522 3300
rect 4630 3350 4632 3351
rect 4668 3350 4670 3351
rect 4630 3300 4631 3350
rect 4669 3300 4670 3350
rect 4772 3350 4774 3351
rect 4630 3299 4632 3300
rect 4668 3299 4670 3300
rect 4772 3300 4773 3350
rect 4772 3299 4774 3300
rect 4810 3350 4812 3351
rect 4811 3300 4812 3350
rect 7605 3350 7607 3351
rect 4810 3299 4812 3300
rect 7605 3300 7606 3350
rect 7605 3299 7607 3300
rect 7643 3350 7645 3351
rect 7644 3300 7645 3350
rect 8258 3448 8260 3449
rect 8296 3448 8298 3449
rect 8258 3386 8259 3448
rect 8297 3386 8298 3448
rect 8258 3385 8260 3386
rect 8296 3385 8298 3386
rect 7749 3350 7751 3351
rect 7787 3350 7789 3351
rect 7643 3299 7645 3300
rect 7749 3300 7750 3350
rect 7788 3300 7789 3350
rect 8007 3338 8065 3339
rect 8007 3337 8008 3338
rect 8064 3337 8065 3338
rect 7749 3299 7751 3300
rect 7787 3299 7789 3300
rect 8007 3300 8008 3301
rect 8064 3300 8065 3301
rect 8007 3299 8065 3300
<< via1 >>
rect 7383 5611 7435 5663
rect 7383 5547 7435 5599
rect 7819 5537 7871 5589
rect 7819 5473 7871 5525
rect 6243 5250 6295 5302
rect 6243 5186 6295 5238
rect 8423 5035 8475 5087
rect 8423 4971 8475 5023
rect 8423 4907 8475 4959
rect 8423 4843 8475 4895
rect 8423 4779 8475 4831
rect 8423 4715 8475 4767
rect 6799 4681 6851 4687
rect 6799 4647 6808 4681
rect 6808 4647 6842 4681
rect 6842 4647 6851 4681
rect 6799 4635 6851 4647
rect 6799 4609 6851 4623
rect 6799 4575 6808 4609
rect 6808 4575 6842 4609
rect 6842 4575 6851 4609
rect 6799 4571 6851 4575
rect 7071 4624 7123 4630
rect 7071 4590 7080 4624
rect 7080 4590 7114 4624
rect 7114 4590 7123 4624
rect 7071 4578 7123 4590
rect 7071 4552 7123 4566
rect 7071 4518 7080 4552
rect 7080 4518 7114 4552
rect 7114 4518 7123 4552
rect 7071 4514 7123 4518
rect 7463 4578 7515 4630
rect 7463 4514 7515 4566
rect 7050 4419 7102 4471
rect 7114 4419 7166 4471
rect 7239 4211 7355 4391
rect 7050 4109 7102 4161
rect 7114 4109 7166 4161
rect 8229 3995 8281 4001
rect 8229 3961 8236 3995
rect 8236 3961 8270 3995
rect 8270 3961 8281 3995
rect 8229 3949 8281 3961
rect 8293 3995 8345 4001
rect 8293 3961 8308 3995
rect 8308 3961 8342 3995
rect 8342 3961 8345 3995
rect 8293 3949 8345 3961
rect 207 3911 259 3917
rect 207 3877 211 3911
rect 211 3877 245 3911
rect 245 3877 259 3911
rect 207 3865 259 3877
rect 271 3911 323 3917
rect 271 3877 283 3911
rect 283 3877 317 3911
rect 317 3877 323 3911
rect 271 3865 323 3877
rect 456 3911 508 3917
rect 456 3877 473 3911
rect 473 3877 507 3911
rect 507 3877 508 3911
rect 456 3865 508 3877
rect 520 3865 572 3917
rect 3632 3865 3684 3917
rect 3696 3911 3748 3917
rect 3696 3877 3697 3911
rect 3697 3877 3731 3911
rect 3731 3877 3748 3911
rect 3696 3865 3748 3877
rect 3881 3911 3933 3917
rect 3881 3877 3887 3911
rect 3887 3877 3921 3911
rect 3921 3877 3933 3911
rect 3881 3865 3933 3877
rect 3945 3911 3997 3917
rect 3945 3877 3959 3911
rect 3959 3877 3993 3911
rect 3993 3877 3997 3911
rect 3945 3865 3997 3877
rect 4411 3911 4463 3917
rect 4411 3877 4415 3911
rect 4415 3877 4449 3911
rect 4449 3877 4463 3911
rect 4411 3865 4463 3877
rect 4475 3911 4527 3917
rect 4475 3877 4487 3911
rect 4487 3877 4521 3911
rect 4521 3877 4527 3911
rect 4475 3865 4527 3877
rect 4660 3911 4712 3917
rect 4660 3877 4677 3911
rect 4677 3877 4711 3911
rect 4711 3877 4712 3911
rect 4660 3865 4712 3877
rect 4724 3865 4776 3917
rect 7600 3865 7652 3917
rect 7664 3865 7716 3917
rect 8033 3871 8085 3923
rect 8097 3911 8149 3923
rect 8097 3877 8125 3911
rect 8125 3877 8149 3911
rect 8097 3871 8149 3877
rect -22 3595 30 3600
rect -22 3561 -17 3595
rect -17 3561 17 3595
rect 17 3561 30 3595
rect -22 3548 30 3561
rect -22 3523 30 3536
rect -22 3489 -17 3523
rect -17 3489 17 3523
rect 17 3489 30 3523
rect -22 3484 30 3489
rect 2149 3548 2201 3600
rect 2218 3548 2270 3600
rect 2287 3548 2339 3600
rect 2149 3484 2201 3536
rect 2218 3484 2270 3536
rect 2287 3484 2339 3536
rect 4037 3548 4089 3600
rect 4106 3548 4158 3600
rect 4175 3548 4227 3600
rect 4037 3484 4089 3536
rect 4106 3484 4158 3536
rect 4175 3484 4227 3536
rect 5183 3548 5235 3600
rect 5259 3548 5311 3600
rect 5335 3548 5387 3600
rect 5410 3548 5462 3600
rect 5485 3548 5537 3600
rect 5183 3484 5235 3536
rect 5259 3484 5311 3536
rect 5335 3484 5387 3536
rect 5410 3484 5462 3536
rect 5485 3484 5537 3536
rect 5974 3483 6090 3599
rect 6158 3548 6210 3600
rect 6224 3548 6276 3600
rect 6290 3548 6342 3600
rect 6355 3548 6407 3600
rect 6158 3484 6210 3536
rect 6224 3484 6276 3536
rect 6290 3484 6342 3536
rect 6355 3484 6407 3536
rect 7206 3548 7258 3600
rect 7329 3548 7381 3600
rect 7206 3484 7258 3536
rect 7329 3484 7381 3536
rect 8158 3491 8338 3607
rect 3506 3397 3558 3449
rect 3570 3397 3622 3449
rect 7670 3391 7722 3443
rect 59 3293 111 3345
rect 59 3229 111 3281
rect 201 3293 253 3345
rect 201 3229 253 3281
rect 491 3293 543 3345
rect 491 3229 543 3281
rect 855 3292 907 3344
rect 855 3228 907 3280
rect 3661 3293 3713 3345
rect 1700 3212 1752 3264
rect 1700 3148 1752 3200
rect 2373 3212 2425 3264
rect 3661 3229 3713 3281
rect 3951 3293 4003 3345
rect 3951 3229 4003 3281
rect 4262 3293 4314 3345
rect 4262 3229 4314 3281
rect 4405 3293 4457 3345
rect 4405 3229 4457 3281
rect 4695 3293 4747 3345
rect 4695 3229 4747 3281
rect 5059 3293 5111 3345
rect 7670 3327 7722 3379
rect 8007 3391 8059 3443
rect 8071 3391 8123 3443
rect 8323 3391 8375 3443
rect 8323 3327 8375 3379
rect 5059 3229 5111 3281
rect 2373 3148 2425 3200
rect 5884 3212 5936 3264
rect 5884 3148 5936 3200
rect 6676 3212 6728 3264
rect 6676 3148 6728 3200
rect 59 2900 111 2952
rect 4029 2900 4081 2952
rect 4262 2900 4314 2952
rect 59 2836 111 2888
rect 4029 2836 4081 2888
rect 4262 2836 4314 2888
rect 8473 2875 8525 2927
rect 8473 2811 8525 2863
rect 3806 2498 3922 2678
rect 4114 2496 4230 2676
rect 7234 2497 7350 2677
rect 4414 2400 4466 2452
rect 4414 2336 4466 2388
rect 6842 1863 6958 2043
rect 3564 1615 3616 1667
rect 3628 1615 3680 1667
rect 4428 1535 4480 1587
rect 4492 1535 4544 1587
rect 7897 1535 7949 1587
rect 7961 1535 8013 1587
rect 1530 1455 1582 1507
rect 1594 1455 1646 1507
rect 2558 1455 2610 1507
rect 2622 1455 2674 1507
rect 5734 1455 5786 1507
rect 5798 1455 5850 1507
rect 145 1332 197 1338
rect 145 1298 153 1332
rect 153 1298 187 1332
rect 187 1298 197 1332
rect 145 1286 197 1298
rect 209 1332 261 1338
rect 209 1298 225 1332
rect 225 1298 259 1332
rect 259 1298 261 1332
rect 209 1286 261 1298
rect 488 1332 540 1344
rect 488 1298 493 1332
rect 493 1298 527 1332
rect 527 1298 540 1332
rect 488 1292 540 1298
rect 552 1332 604 1344
rect 552 1298 565 1332
rect 565 1298 599 1332
rect 599 1298 604 1332
rect 552 1292 604 1298
rect 3806 1041 3922 1221
rect 4115 1041 4231 1221
rect 7237 1037 7353 1217
rect 3628 872 3680 924
rect 7967 886 8019 938
rect 3628 808 3680 860
rect 7967 822 8019 874
rect 6842 365 6958 545
rect 8323 74 8375 126
rect 145 4 197 56
rect 209 4 261 56
rect 785 4 837 56
rect 849 4 901 56
rect 4348 4 4400 56
rect 4412 4 4464 56
rect 4989 4 5041 56
rect 5053 4 5105 56
rect 8323 10 8375 62
<< metal2 >>
rect 7383 5663 7435 5669
rect 6147 5143 6215 5638
rect 6243 5302 6295 5638
rect 6243 5238 6295 5250
rect 6243 5180 6295 5186
tri 6215 5143 6240 5168 sw
tri 6298 5143 6323 5168 se
rect 6323 5143 6415 5638
rect -197 4068 185 4162
rect -197 4001 118 4068
tri 118 4001 185 4068 nw
rect -197 3949 66 4001
tri 66 3949 118 4001 nw
rect -197 3923 40 3949
tri 40 3923 66 3949 nw
rect -197 3917 34 3923
tri 34 3917 40 3923 nw
rect -197 3600 31 3917
tri 31 3914 34 3917 nw
rect -197 3548 -22 3600
rect 30 3548 31 3600
rect -197 3536 31 3548
rect -197 3484 -22 3536
rect 30 3484 31 3536
tri -237 3094 -197 3134 se
rect -197 3094 31 3484
rect 201 3865 207 3917
rect 259 3865 271 3917
rect 323 3865 329 3917
rect 450 3865 456 3917
rect 508 3865 520 3917
rect 572 3865 578 3917
tri 837 3865 847 3875 se
rect 847 3865 979 4162
tri -264 3067 -237 3094 se
rect -237 3067 31 3094
tri -285 3046 -264 3067 se
rect -264 3046 31 3067
rect 59 3345 111 3351
rect 59 3281 111 3293
rect 59 3134 111 3229
rect 201 3345 253 3865
tri 253 3840 278 3865 nw
tri 466 3840 491 3865 ne
rect 201 3281 253 3293
rect 201 3223 253 3229
rect 491 3345 543 3865
tri 543 3840 568 3865 nw
tri 812 3840 837 3865 se
rect 837 3840 979 3865
tri 787 3815 812 3840 se
rect 812 3815 979 3840
tri 961 3548 1007 3594 se
rect 1007 3548 1323 4162
rect 3939 4023 4471 4049
rect 3939 4021 4469 4023
tri 4469 4021 4471 4023 nw
tri 949 3536 961 3548 se
rect 961 3536 1323 3548
tri 935 3522 949 3536 se
rect 949 3522 1323 3536
rect 491 3281 543 3293
rect 491 3223 543 3229
rect 855 3344 907 3350
rect 855 3280 907 3292
tri 111 3134 116 3139 sw
rect 59 3116 116 3134
tri 59 3059 116 3116 ne
tri 116 3059 191 3134 sw
rect -285 2236 31 3046
tri 116 3036 139 3059 ne
tri -285 2148 -197 2236 ne
rect -197 -50 31 2236
rect 59 2952 111 2958
rect 59 2888 111 2900
rect 59 -94 111 2836
rect 139 1344 191 3059
tri 191 1344 210 1363 sw
rect 139 1338 210 1344
tri 210 1338 216 1344 sw
rect 139 1286 145 1338
rect 197 1286 209 1338
rect 261 1286 267 1338
rect 482 1292 488 1344
rect 540 1292 552 1344
rect 604 1292 610 1344
tri 482 1286 488 1292 ne
rect 488 1286 542 1292
rect 139 74 191 1286
tri 191 1261 216 1286 nw
tri 488 1284 490 1286 ne
tri 191 74 198 81 sw
rect 139 62 198 74
tri 198 62 210 74 sw
rect 139 56 210 62
tri 210 56 216 62 sw
rect 139 4 145 56
rect 197 4 209 56
rect 261 4 267 56
tri 190 -21 215 4 ne
rect 215 -94 267 4
rect 490 -94 542 1286
tri 542 1267 567 1292 nw
tri 848 74 855 81 se
rect 855 74 907 3228
tri 836 62 848 74 se
rect 848 62 907 74
tri 830 56 836 62 se
rect 836 56 907 62
rect 779 4 785 56
rect 837 4 849 56
rect 901 4 907 56
rect 935 -50 1323 3522
rect 1444 3270 1496 4021
tri 1496 3270 1507 3281 sw
rect 1444 3264 1507 3270
tri 1507 3264 1513 3270 sw
rect 1700 3264 1752 4021
rect 1444 3256 1513 3264
tri 1513 3256 1521 3264 sw
rect 1444 3212 1496 3256
rect 1700 3200 1752 3212
rect 2143 3600 2345 4021
rect 2143 3548 2149 3600
rect 2201 3548 2218 3600
rect 2270 3548 2287 3600
rect 2339 3548 2345 3600
rect 2143 3536 2345 3548
rect 2143 3484 2149 3536
rect 2201 3484 2218 3536
rect 2270 3484 2287 3536
rect 2339 3484 2345 3536
tri 2131 3148 2143 3160 se
rect 2143 3148 2345 3484
rect 1700 3142 1752 3148
tri 2125 3142 2131 3148 se
rect 2131 3142 2345 3148
rect 2373 3264 2425 4021
tri 2504 3723 2520 3739 se
rect 2520 3723 2572 4021
rect 2373 3200 2425 3212
rect 2373 3142 2425 3148
tri 2460 3679 2504 3723 se
rect 2504 3679 2512 3723
tri 2050 3067 2125 3142 se
rect 2125 3067 2345 3142
tri 2029 3046 2050 3067 se
rect 2050 3046 2345 3067
rect 1524 1507 1652 2716
rect 2029 2236 2345 3046
tri 2029 2122 2143 2236 ne
rect 1524 1455 1530 1507
rect 1582 1455 1594 1507
rect 1646 1455 1652 1507
rect 2143 -50 2345 2236
rect 2460 1310 2512 3679
tri 2512 3663 2572 3723 nw
rect 2632 3270 2684 4021
rect 2790 3560 3152 4021
rect 3180 3594 3496 4021
tri 3939 4001 3959 4021 ne
rect 3959 4001 4449 4021
tri 4449 4001 4469 4021 nw
tri 3959 3949 4011 4001 ne
rect 4011 3949 4397 4001
tri 4397 3949 4449 4001 nw
tri 4011 3929 4031 3949 ne
rect 4031 3929 4377 3949
tri 4377 3929 4397 3949 nw
rect 4031 3923 4371 3929
tri 4371 3923 4377 3929 nw
rect 4031 3917 4365 3923
tri 4365 3917 4371 3923 nw
rect 3626 3865 3632 3917
rect 3684 3865 3696 3917
rect 3748 3865 3754 3917
rect 3875 3865 3881 3917
rect 3933 3865 3945 3917
rect 3997 3865 4003 3917
tri 3636 3840 3661 3865 ne
tri 3180 3582 3192 3594 ne
rect 3192 3582 3496 3594
tri 3152 3560 3174 3582 sw
tri 3192 3566 3208 3582 ne
tri 2684 3270 2695 3281 sw
rect 2632 3256 2695 3270
tri 2695 3256 2709 3270 sw
rect 2632 3218 2684 3256
rect 2552 1507 2680 2716
rect 2552 1455 2558 1507
rect 2610 1455 2622 1507
rect 2674 1455 2680 1507
rect 2790 1875 3174 3560
rect 3208 3525 3496 3582
rect 3208 3484 3455 3525
tri 3455 3484 3496 3525 nw
rect 3208 3483 3454 3484
tri 3454 3483 3455 3484 nw
rect 3208 3449 3420 3483
tri 3420 3449 3454 3483 nw
rect 3208 3397 3368 3449
tri 3368 3397 3420 3449 nw
rect 3500 3397 3506 3449
rect 3558 3397 3570 3449
rect 3622 3397 3628 3449
rect 3208 3391 3362 3397
tri 3362 3391 3368 3397 nw
tri 3539 3391 3545 3397 ne
rect 3545 3391 3628 3397
rect 3208 1955 3358 3391
tri 3358 3387 3362 3391 nw
tri 3545 3387 3549 3391 ne
rect 3549 3387 3628 3391
tri 3549 3379 3557 3387 ne
rect 3557 3379 3628 3387
tri 3557 3372 3564 3379 ne
rect 3564 3200 3628 3379
rect 3661 3345 3713 3865
tri 3713 3840 3738 3865 nw
tri 3926 3840 3951 3865 ne
rect 3661 3281 3713 3293
rect 3661 3223 3713 3229
rect 3951 3345 4003 3865
rect 3951 3281 4003 3293
rect 3951 3223 4003 3229
rect 4031 3865 4313 3917
tri 4313 3865 4365 3917 nw
rect 4405 3865 4411 3917
rect 4463 3865 4475 3917
rect 4527 3865 4533 3917
rect 4654 3865 4660 3917
rect 4712 3865 4724 3917
rect 4776 3865 4782 3917
rect 4031 3600 4236 3865
tri 4236 3788 4313 3865 nw
rect 4405 3854 4471 3865
tri 4471 3854 4482 3865 nw
tri 4670 3854 4681 3865 ne
rect 4681 3854 4747 3865
rect 4031 3548 4037 3600
rect 4089 3548 4106 3600
rect 4158 3548 4175 3600
rect 4227 3548 4236 3600
rect 4031 3536 4236 3548
rect 4031 3484 4037 3536
rect 4089 3484 4106 3536
rect 4158 3484 4175 3536
rect 4227 3484 4236 3536
rect 4031 3416 4236 3484
tri 3628 3200 3634 3206 sw
rect 3564 3179 3634 3200
tri 3564 3148 3595 3179 ne
rect 3595 3148 3634 3179
tri 3634 3148 3686 3200 sw
tri 3595 3121 3622 3148 ne
tri 3208 1909 3254 1955 ne
rect 3254 1909 3358 1955
tri 3358 1909 3468 2019 sw
tri 3174 1875 3208 1909 sw
tri 3254 1881 3282 1909 ne
rect 3282 1881 3468 1909
tri 3468 1881 3496 1909 sw
tri 3282 1875 3288 1881 ne
rect 3288 1875 3496 1881
rect 2790 1863 3208 1875
tri 3208 1863 3220 1875 sw
tri 3288 1863 3300 1875 ne
rect 3300 1863 3496 1875
rect 2790 1817 3220 1863
tri 3220 1817 3266 1863 sw
tri 3300 1817 3346 1863 ne
rect 2790 1793 3266 1817
tri 3266 1793 3290 1817 sw
tri 2460 1266 2504 1310 ne
rect 2504 1266 2512 1310
tri 2512 1266 2572 1326 sw
tri 2504 1258 2512 1266 ne
rect 2512 1258 2572 1266
tri 2512 1250 2520 1258 ne
rect 2520 -94 2572 1258
tri 2778 455 2790 467 se
rect 2790 455 3290 1793
rect 2778 264 3290 455
tri 2778 252 2790 264 ne
rect 2790 -50 3290 264
rect 3346 -50 3496 1863
tri 3597 1667 3622 1692 se
rect 3622 1667 3686 3148
rect 4031 3003 4234 3416
tri 4234 3414 4236 3416 nw
rect 4262 3345 4314 3351
rect 4262 3281 4314 3293
rect 4262 3172 4314 3229
rect 4405 3345 4457 3854
tri 4457 3840 4471 3854 nw
tri 4681 3840 4695 3854 ne
rect 4405 3281 4457 3293
rect 4405 3223 4457 3229
rect 4695 3345 4747 3854
tri 4747 3840 4772 3865 nw
rect 5175 3600 5547 4021
rect 5175 3548 5183 3600
rect 5235 3548 5259 3600
rect 5311 3548 5335 3600
rect 5387 3548 5410 3600
rect 5462 3548 5485 3600
rect 5537 3548 5547 3600
rect 5175 3536 5547 3548
rect 5175 3484 5183 3536
rect 5235 3484 5259 3536
rect 5311 3484 5335 3536
rect 5387 3484 5410 3536
rect 5462 3484 5485 3536
rect 5537 3484 5547 3536
rect 4695 3281 4747 3293
rect 4695 3223 4747 3229
rect 5059 3345 5111 3351
rect 5059 3281 5111 3293
tri 4314 3172 4336 3194 sw
tri 4262 3166 4268 3172 ne
rect 4268 3166 4336 3172
tri 4336 3166 4342 3172 sw
tri 4268 3148 4286 3166 ne
rect 4286 3148 4342 3166
tri 4342 3148 4360 3166 sw
tri 4286 3092 4342 3148 ne
rect 4342 3114 4360 3148
tri 4360 3114 4394 3148 sw
tri 4084 2978 4109 3003 ne
rect 4029 2952 4081 2958
rect 4029 2888 4081 2900
tri 3858 2684 3883 2709 sw
rect 3558 1615 3564 1667
rect 3616 1615 3628 1667
rect 3680 1615 3686 1667
tri 3597 1590 3622 1615 ne
rect 3622 924 3686 1615
rect 3806 2678 3922 2684
rect 3806 1221 3922 2498
rect 3806 1035 3922 1041
rect 3622 872 3628 924
rect 3680 872 3686 924
rect 3622 860 3686 872
rect 3622 808 3628 860
rect 3680 808 3686 860
rect 4029 -94 4081 2836
rect 4109 2676 4234 3003
rect 4109 2496 4114 2676
rect 4230 2496 4234 2676
rect 4109 1221 4234 2496
rect 4109 1041 4115 1221
rect 4231 1041 4234 1221
rect 4109 -50 4234 1041
rect 4262 2952 4314 2958
rect 4262 2888 4314 2900
rect 4262 -94 4314 2836
rect 4342 2480 4394 3114
rect 4342 2307 4386 2480
tri 4386 2472 4394 2480 nw
rect 4414 2452 4474 2458
rect 4466 2400 4474 2452
rect 4414 2388 4474 2400
rect 4466 2336 4474 2388
rect 4414 2330 4474 2336
tri 4414 2322 4422 2330 ne
tri 4386 2307 4394 2315 sw
rect 4342 74 4394 2307
rect 4422 1587 4474 2330
tri 4474 1587 4499 1612 sw
rect 4422 1535 4428 1587
rect 4480 1535 4492 1587
rect 4544 1535 4550 1587
rect 4624 332 4944 2043
tri 4394 74 4401 81 sw
tri 5052 74 5059 81 se
rect 5059 74 5111 3229
rect 4342 62 4401 74
tri 4401 62 4413 74 sw
tri 5040 62 5052 74 se
rect 5052 62 5111 74
rect 4342 56 4413 62
tri 4413 56 4419 62 sw
tri 5034 56 5040 62 se
rect 5040 56 5111 62
rect 4342 4 4348 56
rect 4400 4 4412 56
rect 4464 4 4470 56
rect 4983 4 4989 56
rect 5041 4 5053 56
rect 5105 4 5111 56
rect 5175 -50 5547 3484
rect 5648 3270 5700 4021
tri 5700 3270 5711 3281 sw
rect 5648 3264 5711 3270
tri 5711 3264 5717 3270 sw
rect 5884 3264 5936 4021
rect 5648 3256 5717 3264
tri 5717 3256 5725 3264 sw
rect 5648 3212 5700 3256
rect 5884 3200 5936 3212
rect 5884 3142 5936 3148
rect 5974 3599 6090 3607
tri 5948 3114 5974 3140 se
rect 5974 3114 6090 3483
rect 5948 3092 6090 3114
rect 6147 3600 6415 5143
rect 6147 3548 6158 3600
rect 6210 3548 6224 3600
rect 6276 3548 6290 3600
rect 6342 3548 6355 3600
rect 6407 3548 6415 3600
rect 6147 3536 6415 3548
rect 6147 3484 6158 3536
rect 6210 3484 6224 3536
rect 6276 3484 6290 3536
rect 6342 3484 6355 3536
rect 6407 3484 6415 3536
rect 5728 1507 5856 2716
rect 5948 1507 6064 3092
tri 6064 3066 6090 3092 nw
tri 6119 3066 6147 3094 se
rect 6147 3066 6415 3484
tri 6099 3046 6119 3066 se
rect 6119 3046 6415 3066
rect 6099 2236 6415 3046
tri 6099 2188 6147 2236 ne
rect 5728 1455 5734 1507
rect 5786 1455 5798 1507
rect 5850 1455 5856 1507
rect 6147 -50 6415 2236
rect 6471 2677 6648 5638
rect 6676 3264 6728 5638
tri 6793 4687 6799 4693 se
rect 6799 4687 6851 5638
tri 6851 4687 6857 4693 sw
rect 6793 4635 6799 4687
rect 6851 4635 6857 4687
rect 6793 4623 6857 4635
rect 6793 4571 6799 4623
rect 6851 4571 6857 4623
tri 6887 3256 6912 3281 se
rect 6912 3212 6964 5638
rect 7071 4630 7123 5638
rect 7151 5473 7327 5638
rect 7383 5599 7435 5611
rect 7383 5541 7435 5547
tri 7327 5473 7370 5516 sw
rect 7151 5456 7370 5473
tri 7370 5456 7387 5473 sw
rect 7151 5382 7387 5456
tri 7151 5333 7200 5382 ne
rect 7071 4566 7123 4578
rect 7071 4508 7123 4514
rect 7044 4419 7050 4471
rect 7102 4419 7114 4471
rect 7166 4419 7172 4471
rect 7044 4161 7172 4419
rect 7044 4109 7050 4161
rect 7102 4109 7114 4161
rect 7166 4109 7172 4161
rect 6676 3200 6728 3212
rect 6676 3142 6728 3148
tri 6648 2677 6733 2762 sw
rect 6471 2619 6733 2677
tri 6733 2619 6791 2677 sw
rect 6471 -50 6791 2619
rect 6836 1863 6842 2043
rect 6958 1863 6964 2043
rect 6836 545 6964 1863
rect 7044 1507 7172 4109
rect 7200 4391 7387 5382
rect 7463 4630 7515 5638
rect 7463 4566 7515 4578
rect 7463 4508 7515 4514
tri 7518 4391 7543 4416 se
rect 7543 4391 7711 5638
rect 7819 5589 7871 5638
rect 7819 5525 7871 5537
rect 7819 5467 7871 5473
rect 7200 4211 7239 4391
rect 7355 4211 7387 4391
rect 7434 4211 7711 4391
tri 7860 5325 7899 5364 se
rect 7899 5325 8083 5638
tri 7826 4282 7860 4316 se
rect 7860 4282 8083 5325
tri 7755 4211 7826 4282 se
rect 7826 4211 8083 4282
rect 7200 3600 7387 4211
tri 7716 4172 7755 4211 se
rect 7755 4172 8083 4211
rect 7200 3548 7206 3600
rect 7258 3548 7329 3600
rect 7381 3548 7387 3600
rect 7200 3536 7387 3548
rect 7200 3484 7206 3536
rect 7258 3484 7329 3536
rect 7381 3484 7387 3536
rect 7200 2677 7387 3484
rect 7200 2497 7234 2677
rect 7350 2497 7387 2677
rect 6836 365 6842 545
rect 6958 365 6964 545
rect 7200 1217 7387 2497
rect 7200 1037 7237 1217
rect 7353 1037 7387 1217
rect 7200 -50 7387 1037
rect 7415 4069 8083 4172
rect 7415 4009 8023 4069
tri 8023 4009 8083 4069 nw
rect 8139 4047 8361 5638
tri 8139 4009 8177 4047 ne
rect 7415 4001 8015 4009
tri 8015 4001 8023 4009 nw
rect 8177 4001 8361 4047
rect 7415 3958 7973 4001
tri 7973 3959 8015 4001 nw
rect 7415 3949 7580 3958
tri 7580 3949 7589 3958 nw
tri 7723 3949 7732 3958 ne
rect 7732 3949 7973 3958
rect 7415 2030 7562 3949
tri 7562 3931 7580 3949 nw
tri 7732 3931 7750 3949 ne
rect 7594 3865 7600 3917
rect 7652 3865 7664 3917
rect 7716 3865 7722 3917
tri 7645 3840 7670 3865 ne
rect 7670 3443 7722 3865
rect 7670 3379 7722 3391
rect 7670 3321 7722 3327
rect 7750 2440 7973 3949
rect 8177 3949 8229 4001
rect 8281 3949 8293 4001
rect 8345 3949 8361 4001
rect 8033 3923 8149 3929
rect 8085 3871 8097 3923
rect 8033 3865 8149 3871
rect 8033 3840 8124 3865
tri 8124 3840 8149 3865 nw
rect 8033 3475 8085 3840
tri 8085 3801 8124 3840 nw
tri 8151 3808 8177 3834 se
rect 8177 3808 8361 3949
rect 8151 3607 8361 3808
rect 8151 3491 8158 3607
rect 8338 3491 8361 3607
rect 8417 5087 8728 5638
rect 8417 5035 8423 5087
rect 8475 5035 8728 5087
rect 8417 5023 8728 5035
rect 8417 4971 8423 5023
rect 8475 4971 8728 5023
rect 8417 4959 8728 4971
rect 8417 4907 8423 4959
rect 8475 4907 8728 4959
rect 8417 4895 8728 4907
rect 8417 4843 8423 4895
rect 8475 4843 8728 4895
rect 8417 4831 8728 4843
rect 8417 4779 8423 4831
rect 8475 4779 8728 4831
rect 8417 4767 8728 4779
rect 8417 4715 8423 4767
rect 8475 4715 8728 4767
rect 8151 3487 8321 3491
tri 8321 3487 8325 3491 nw
tri 8085 3475 8097 3487 sw
rect 8151 3475 8309 3487
tri 8309 3475 8321 3487 nw
tri 8007 3449 8033 3475 se
rect 8033 3449 8097 3475
tri 8097 3449 8123 3475 sw
rect 8007 3443 8123 3449
rect 8059 3391 8071 3443
rect 8007 3385 8123 3391
tri 7750 2364 7826 2440 ne
tri 7781 2059 7826 2104 se
rect 7826 2059 7973 2440
tri 7562 2030 7591 2059 sw
tri 7752 2030 7781 2059 se
rect 7781 2030 7973 2059
rect 7415 1896 7973 2030
rect 7415 878 7731 1896
tri 7731 1654 7973 1896 nw
tri 8139 3361 8151 3373 se
rect 8151 3361 8295 3475
tri 8295 3461 8309 3475 nw
rect 7891 1535 7897 1587
rect 7949 1535 7961 1587
rect 8013 1535 8019 1587
tri 7942 1510 7967 1535 ne
rect 7415 874 7727 878
tri 7727 874 7731 878 nw
rect 7967 938 8019 1535
rect 7967 874 8019 886
rect 7415 822 7675 874
tri 7675 822 7727 874 nw
rect 7415 816 7669 822
tri 7669 816 7675 822 nw
rect 7967 816 8019 822
rect 7415 -50 7599 816
tri 7599 746 7669 816 nw
rect 8139 -50 8295 3361
rect 8323 3443 8375 3449
rect 8323 3379 8375 3391
rect 8323 126 8375 3327
rect 8417 2964 8728 4715
rect 8323 62 8375 74
rect 8323 4 8375 10
rect 8459 2927 8525 2933
rect 8459 2875 8473 2927
rect 8459 2863 8525 2875
rect 8459 2811 8473 2863
rect 8459 2805 8525 2811
rect 8459 -94 8511 2805
tri 8511 2791 8525 2805 nw
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_0
timestamp 1707688321
transform 0 1 7893 1 0 3877
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_1
timestamp 1707688321
transform 0 1 8091 1 0 3877
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_2
timestamp 1707688321
transform 1 0 1969 0 -1 842
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_3
timestamp 1707688321
transform 1 0 2321 0 -1 842
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_4
timestamp 1707688321
transform 1 0 2673 0 -1 842
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_5
timestamp 1707688321
transform 1 0 3025 0 -1 842
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_6
timestamp 1707688321
transform 1 0 3377 0 -1 842
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_7
timestamp 1707688321
transform 1 0 4081 0 -1 842
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_8
timestamp 1707688321
transform 1 0 4433 0 -1 842
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_9
timestamp 1707688321
transform 1 0 4572 0 -1 842
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_10
timestamp 1707688321
transform 1 0 1617 0 -1 842
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_11
timestamp 1707688321
transform 1 0 1265 0 -1 842
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_12
timestamp 1707688321
transform 1 0 913 0 -1 842
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_13
timestamp 1707688321
transform 1 0 275 0 -1 842
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_14
timestamp 1707688321
transform 1 0 -17 0 1 886
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_15
timestamp 1707688321
transform 1 0 4433 0 1 886
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_16
timestamp 1707688321
transform 1 0 1617 0 1 886
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_17
timestamp 1707688321
transform 1 0 913 0 1 886
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_18
timestamp 1707688321
transform 1 0 275 0 1 886
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_19
timestamp 1707688321
transform 1 0 6808 0 1 4575
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_0
timestamp 1707688321
transform 0 -1 7114 -1 0 4624
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_1
timestamp 1707688321
transform 0 -1 17 -1 0 3595
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_2
timestamp 1707688321
transform 0 -1 7610 -1 0 4624
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_3
timestamp 1707688321
transform -1 0 3993 0 1 3877
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_4
timestamp 1707688321
transform -1 0 3803 0 1 3877
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_5
timestamp 1707688321
transform 0 -1 8259 1 0 2158
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_6
timestamp 1707688321
transform 1 0 493 0 1 1298
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_7
timestamp 1707688321
transform 1 0 401 0 1 3877
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_8
timestamp 1707688321
transform 1 0 211 0 1 3877
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_9
timestamp 1707688321
transform 1 0 4415 0 1 3877
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_10
timestamp 1707688321
transform 1 0 4605 0 1 3877
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_11
timestamp 1707688321
transform 1 0 1150 0 1 3409
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_12
timestamp 1707688321
transform 1 0 2948 0 1 3409
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_13
timestamp 1707688321
transform 1 0 5354 0 1 3409
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_14
timestamp 1707688321
transform 1 0 7152 0 1 3409
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_15
timestamp 1707688321
transform 1 0 153 0 1 1298
box 0 0 1 1
use L1M1_CDNS_5246887918590  L1M1_CDNS_5246887918590_0
timestamp 1707688321
transform -1 0 8414 0 1 3961
box 0 0 1 1
use L1M1_CDNS_52468879185194  L1M1_CDNS_52468879185194_0
timestamp 1707688321
transform 0 -1 17 -1 0 764
box -12 -6 766 40
use L1M1_CDNS_52468879185308  L1M1_CDNS_52468879185308_0
timestamp 1707688321
transform 0 -1 8131 1 0 1055
box 0 0 1 1
use L1M1_CDNS_52468879185501  L1M1_CDNS_52468879185501_0
timestamp 1707688321
transform 1 0 -17 0 1 958
box 0 0 1 1
use L1M1_CDNS_52468879185945  L1M1_CDNS_52468879185945_0
timestamp 1707688321
transform 1 0 6106 0 1 3961
box -12 -6 1846 40
use L1M1_CDNS_524688791851104  L1M1_CDNS_524688791851104_0
timestamp 1707688321
transform 1 0 10 0 1 -68
box -12 -6 4582 40
use L1M1_CDNS_524688791851153  L1M1_CDNS_524688791851153_0
timestamp 1707688321
transform -1 0 4847 0 1 1467
box -12 -6 4798 40
use L1M1_CDNS_524688791851154  L1M1_CDNS_524688791851154_0
timestamp 1707688321
transform 1 0 5142 0 -1 272
box -12 -6 1702 112
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_0
timestamp 1707688321
transform 0 -1 4081 -1 0 2958
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_1
timestamp 1707688321
transform 0 -1 8375 -1 0 132
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_2
timestamp 1707688321
transform 0 -1 5936 -1 0 3270
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_3
timestamp 1707688321
transform 0 -1 4314 -1 0 2958
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_4
timestamp 1707688321
transform 0 1 4414 -1 0 2458
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_5
timestamp 1707688321
transform 0 1 59 -1 0 2958
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_6
timestamp 1707688321
transform 0 1 7071 -1 0 4636
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_7
timestamp 1707688321
transform 0 1 7463 -1 0 4636
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_8
timestamp 1707688321
transform -1 0 3628 0 1 3397
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_9
timestamp 1707688321
transform -1 0 4003 0 1 3865
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_10
timestamp 1707688321
transform -1 0 3754 0 1 3865
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_11
timestamp 1707688321
transform -1 0 7722 0 1 3865
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_12
timestamp 1707688321
transform -1 0 8351 0 1 3949
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_13
timestamp 1707688321
transform -1 0 3686 0 -1 1667
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_14
timestamp 1707688321
transform -1 0 4550 0 -1 1587
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_15
timestamp 1707688321
transform 0 1 8473 1 0 2805
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_16
timestamp 1707688321
transform 0 1 3951 1 0 3223
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_17
timestamp 1707688321
transform 0 1 3661 1 0 3223
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_18
timestamp 1707688321
transform 0 1 7670 1 0 3321
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_19
timestamp 1707688321
transform 0 1 8323 1 0 3321
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_20
timestamp 1707688321
transform 0 -1 7871 1 0 5467
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_21
timestamp 1707688321
transform 0 -1 8019 1 0 816
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_22
timestamp 1707688321
transform 0 -1 1752 1 0 3142
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_23
timestamp 1707688321
transform 0 -1 543 1 0 3223
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_24
timestamp 1707688321
transform 0 -1 253 1 0 3223
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_25
timestamp 1707688321
transform 0 -1 4457 1 0 3223
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_26
timestamp 1707688321
transform 0 -1 4747 1 0 3223
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_27
timestamp 1707688321
transform 0 -1 111 1 0 3223
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_28
timestamp 1707688321
transform 0 -1 4314 1 0 3223
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_29
timestamp 1707688321
transform 0 -1 907 1 0 3222
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_30
timestamp 1707688321
transform 0 -1 5111 1 0 3223
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_31
timestamp 1707688321
transform 0 -1 6295 1 0 5180
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_32
timestamp 1707688321
transform 0 -1 7435 1 0 5541
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_33
timestamp 1707688321
transform 0 -1 6728 1 0 3142
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_34
timestamp 1707688321
transform 0 -1 2425 1 0 3142
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_35
timestamp 1707688321
transform 1 0 7891 0 -1 1587
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_36
timestamp 1707688321
transform 1 0 7044 0 1 4419
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_37
timestamp 1707688321
transform 1 0 7044 0 1 4109
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_38
timestamp 1707688321
transform 1 0 450 0 1 3865
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_39
timestamp 1707688321
transform 1 0 201 0 1 3865
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_40
timestamp 1707688321
transform 1 0 4405 0 1 3865
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_41
timestamp 1707688321
transform 1 0 4654 0 1 3865
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_42
timestamp 1707688321
transform 1 0 139 0 1 4
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_43
timestamp 1707688321
transform 1 0 4342 0 1 4
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_44
timestamp 1707688321
transform 1 0 779 0 1 4
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_45
timestamp 1707688321
transform 1 0 4983 0 1 4
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_46
timestamp 1707688321
transform 1 0 5728 0 1 1455
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_47
timestamp 1707688321
transform 1 0 2552 0 1 1455
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_48
timestamp 1707688321
transform 1 0 1524 0 1 1455
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_49
timestamp 1707688321
transform 1 0 482 0 1 1292
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_50
timestamp 1707688321
transform 1 0 139 0 1 1286
box 0 0 1 1
use M1M2_CDNS_52468879185198  M1M2_CDNS_52468879185198_0
timestamp 1707688321
transform 0 1 3806 -1 0 1227
box 0 0 1 1
use M1M2_CDNS_52468879185198  M1M2_CDNS_52468879185198_1
timestamp 1707688321
transform 0 1 3806 -1 0 2684
box 0 0 1 1
use M1M2_CDNS_52468879185198  M1M2_CDNS_52468879185198_2
timestamp 1707688321
transform 0 1 4114 1 0 2490
box 0 0 1 1
use M1M2_CDNS_52468879185198  M1M2_CDNS_52468879185198_3
timestamp 1707688321
transform 0 1 4115 1 0 1035
box 0 0 1 1
use M1M2_CDNS_52468879185198  M1M2_CDNS_52468879185198_4
timestamp 1707688321
transform 1 0 8152 0 1 3491
box 0 0 1 1
use M1M2_CDNS_52468879185199  M1M2_CDNS_52468879185199_0
timestamp 1707688321
transform 0 1 5974 1 0 3477
box 0 0 1 1
use M1M2_CDNS_52468879185200  M1M2_CDNS_52468879185200_0
timestamp 1707688321
transform 1 0 7233 0 -1 4391
box 0 0 1 1
use M1M2_CDNS_52468879185200  M1M2_CDNS_52468879185200_1
timestamp 1707688321
transform 1 0 6836 0 -1 545
box 0 0 1 1
use M1M2_CDNS_52468879185200  M1M2_CDNS_52468879185200_2
timestamp 1707688321
transform 1 0 6836 0 -1 2043
box 0 0 1 1
use M1M2_CDNS_52468879185200  M1M2_CDNS_52468879185200_3
timestamp 1707688321
transform 1 0 7228 0 1 2497
box 0 0 1 1
use M1M2_CDNS_52468879185200  M1M2_CDNS_52468879185200_4
timestamp 1707688321
transform 1 0 7231 0 1 1037
box 0 0 1 1
use M1M2_CDNS_52468879185201  M1M2_CDNS_52468879185201_0
timestamp 1707688321
transform 1 0 6471 0 -1 278
box 0 0 320 116
use M1M2_CDNS_52468879185201  M1M2_CDNS_52468879185201_1
timestamp 1707688321
transform 1 0 6471 0 -1 1813
box 0 0 320 116
use M1M2_CDNS_52468879185208  M1M2_CDNS_52468879185208_0
timestamp 1707688321
transform 1 0 7876 0 1 4970
box 0 0 192 244
use M1M2_CDNS_52468879185209  M1M2_CDNS_52468879185209_0
timestamp 1707688321
transform 1 0 935 0 -1 776
box 0 0 128 244
use M1M2_CDNS_52468879185209  M1M2_CDNS_52468879185209_1
timestamp 1707688321
transform 1 0 3359 0 1 514
box 0 0 128 244
use M1M2_CDNS_52468879185209  M1M2_CDNS_52468879185209_2
timestamp 1707688321
transform 1 0 8417 0 1 3635
box 0 0 128 244
use M1M2_CDNS_52468879185369  M1M2_CDNS_52468879185369_0
timestamp 1707688321
transform -1 0 6857 0 1 4571
box 0 0 1 1
use M1M2_CDNS_52468879185369  M1M2_CDNS_52468879185369_1
timestamp 1707688321
transform 0 -1 8149 1 0 3865
box 0 0 1 1
use M1M2_CDNS_52468879185369  M1M2_CDNS_52468879185369_2
timestamp 1707688321
transform 0 -1 8123 1 0 3385
box 0 0 1 1
use M1M2_CDNS_52468879185369  M1M2_CDNS_52468879185369_3
timestamp 1707688321
transform 1 0 3622 0 -1 924
box 0 0 1 1
use M1M2_CDNS_52468879185959  M1M2_CDNS_52468879185959_0
timestamp 1707688321
transform 1 0 8417 0 1 4715
box 0 0 1 1
use M1M2_CDNS_52468879185975  M1M2_CDNS_52468879185975_0
timestamp 1707688321
transform -1 0 979 0 1 3635
box 0 0 192 180
use M1M2_CDNS_52468879185975  M1M2_CDNS_52468879185975_1
timestamp 1707688321
transform -1 0 31 0 1 1037
box 0 0 192 180
use M1M2_CDNS_52468879185975  M1M2_CDNS_52468879185975_2
timestamp 1707688321
transform -1 0 31 0 1 2497
box 0 0 192 180
use M1M2_CDNS_52468879185975  M1M2_CDNS_52468879185975_3
timestamp 1707688321
transform 1 0 2148 0 1 2497
box 0 0 192 180
use M1M2_CDNS_52468879185975  M1M2_CDNS_52468879185975_4
timestamp 1707688321
transform 1 0 2148 0 1 1037
box 0 0 192 180
use M1M2_CDNS_524688791851032  M1M2_CDNS_524688791851032_0
timestamp 1707688321
transform -1 0 8348 0 1 4109
box 0 0 192 372
use M1M2_CDNS_524688791851077  M1M2_CDNS_524688791851077_0
timestamp 1707688321
transform 1 0 4624 0 -1 2043
box 0 0 320 180
use M1M2_CDNS_524688791851077  M1M2_CDNS_524688791851077_1
timestamp 1707688321
transform 1 0 5201 0 1 1037
box 0 0 320 180
use M1M2_CDNS_524688791851077  M1M2_CDNS_524688791851077_2
timestamp 1707688321
transform 1 0 5201 0 1 2497
box 0 0 320 180
use M1M2_CDNS_524688791851081  M1M2_CDNS_524688791851081_0
timestamp 1707688321
transform 1 0 4674 0 -1 518
box 0 0 256 180
use M1M2_CDNS_524688791851081  M1M2_CDNS_524688791851081_1
timestamp 1707688321
transform 1 0 7441 0 -1 4391
box 0 0 256 180
use M1M2_CDNS_524688791851081  M1M2_CDNS_524688791851081_2
timestamp 1707688321
transform 1 0 6152 0 -1 4391
box 0 0 256 180
use M1M2_CDNS_524688791851081  M1M2_CDNS_524688791851081_3
timestamp 1707688321
transform 1 0 6154 0 1 2497
box 0 0 256 180
use M1M2_CDNS_524688791851081  M1M2_CDNS_524688791851081_4
timestamp 1707688321
transform 1 0 6154 0 1 1037
box 0 0 256 180
use M1M2_CDNS_524688791851144  M1M2_CDNS_524688791851144_0
timestamp 1707688321
transform 1 0 2790 0 1 1853
box 0 0 384 180
use M1M2_CDNS_524688791851150  M1M2_CDNS_524688791851150_0
timestamp 1707688321
transform 1 0 1063 0 -1 776
box 0 0 256 244
use M1M2_CDNS_524688791851151  M1M2_CDNS_524688791851151_0
timestamp 1707688321
transform 1 0 2778 0 1 264
box 0 0 512 180
use M1M2_CDNS_524688791851152  M1M2_CDNS_524688791851152_0
timestamp 1707688321
transform 0 1 8139 1 0 573
box 0 0 896 116
use sky130_fd_io__refgen_com_ctl_hld_refgen  sky130_fd_io__refgen_com_ctl_hld_refgen_0
timestamp 1707688321
transform 1 0 -38 0 1 -25
box 63 12 8211 1555
use sky130_fd_io__refgen_com_ctl_ls  sky130_fd_io__refgen_com_ctl_ls_0
timestamp 1707688321
transform -1 0 2102 0 -1 3927
box -91 0 2150 2319
use sky130_fd_io__refgen_com_ctl_ls  sky130_fd_io__refgen_com_ctl_ls_1
timestamp 1707688321
transform -1 0 6306 0 -1 3927
box -91 0 2150 2319
use sky130_fd_io__refgen_com_ctl_ls  sky130_fd_io__refgen_com_ctl_ls_2
timestamp 1707688321
transform 1 0 2102 0 -1 3927
box -91 0 2150 2319
use sky130_fd_io__refgen_com_ctl_ls  sky130_fd_io__refgen_com_ctl_ls_3
timestamp 1707688321
transform 1 0 6306 0 -1 3927
box -91 0 2150 2319
use sky130_fd_io__refgen_em1o_CDNS_524688791851126  sky130_fd_io__refgen_em1o_CDNS_524688791851126_0
timestamp 1707688321
transform 0 1 8007 -1 0 3391
box 0 0 1 1
use sky130_fd_io__refgen_em1o_CDNS_524688791851127  sky130_fd_io__refgen_em1o_CDNS_524688791851127_0
timestamp 1707688321
transform -1 0 660 0 1 3299
box 0 0 1 1
use sky130_fd_io__refgen_em1o_CDNS_524688791851127  sky130_fd_io__refgen_em1o_CDNS_524688791851127_1
timestamp 1707688321
transform -1 0 4864 0 1 3299
box 0 0 1 1
use sky130_fd_io__refgen_em1o_CDNS_524688791851127  sky130_fd_io__refgen_em1o_CDNS_524688791851127_2
timestamp 1707688321
transform -1 0 3978 0 -1 3351
box 0 0 1 1
use sky130_fd_io__refgen_em1o_CDNS_524688791851127  sky130_fd_io__refgen_em1o_CDNS_524688791851127_3
timestamp 1707688321
transform 1 0 226 0 -1 3351
box 0 0 1 1
use sky130_fd_io__refgen_em1o_CDNS_524688791851127  sky130_fd_io__refgen_em1o_CDNS_524688791851127_4
timestamp 1707688321
transform 1 0 4430 0 -1 3351
box 0 0 1 1
use sky130_fd_io__refgen_em1o_CDNS_524688791851127  sky130_fd_io__refgen_em1o_CDNS_524688791851127_5
timestamp 1707688321
transform 1 0 3544 0 1 3299
box 0 0 1 1
use sky130_fd_io__refgen_em1o_CDNS_524688791851127  sky130_fd_io__refgen_em1o_CDNS_524688791851127_6
timestamp 1707688321
transform 1 0 7553 0 1 3299
box 0 0 1 1
use sky130_fd_io__refgen_em1s_CDNS_524688791851128  sky130_fd_io__refgen_em1s_CDNS_524688791851128_0
timestamp 1707688321
transform -1 0 518 0 1 3299
box 0 0 1 1
use sky130_fd_io__refgen_em1s_CDNS_524688791851128  sky130_fd_io__refgen_em1s_CDNS_524688791851128_1
timestamp 1707688321
transform -1 0 4722 0 1 3299
box 0 0 1 1
use sky130_fd_io__refgen_em1s_CDNS_524688791851128  sky130_fd_io__refgen_em1s_CDNS_524688791851128_2
timestamp 1707688321
transform -1 0 4120 0 1 3299
box 0 0 1 1
use sky130_fd_io__refgen_em1s_CDNS_524688791851128  sky130_fd_io__refgen_em1s_CDNS_524688791851128_3
timestamp 1707688321
transform 1 0 84 0 1 3299
box 0 0 1 1
use sky130_fd_io__refgen_em1s_CDNS_524688791851128  sky130_fd_io__refgen_em1s_CDNS_524688791851128_4
timestamp 1707688321
transform 1 0 3686 0 1 3299
box 0 0 1 1
use sky130_fd_io__refgen_em1s_CDNS_524688791851128  sky130_fd_io__refgen_em1s_CDNS_524688791851128_5
timestamp 1707688321
transform 1 0 4288 0 1 3299
box 0 0 1 1
use sky130_fd_io__refgen_em1s_CDNS_524688791851128  sky130_fd_io__refgen_em1s_CDNS_524688791851128_6
timestamp 1707688321
transform 1 0 7697 0 1 3299
box 0 0 1 1
use sky130_fd_io__refgen_em1s_CDNS_524688791851166  sky130_fd_io__refgen_em1s_CDNS_524688791851166_0
timestamp 1707688321
transform -1 0 8350 0 1 3385
box 0 0 1 1
use sky130_fd_io__refgen_vpwrka_ls  sky130_fd_io__refgen_vpwrka_ls_0
timestamp 1707688321
transform -1 0 7695 0 -1 5302
box -147 -161 1123 1332
<< labels >>
flabel comment s 7417 5612 7417 5612 3 FreeSans 200 270 0 0 vohref_0p5
flabel comment s 7852 5609 7852 5609 3 FreeSans 200 270 0 0 sel_vohref_op5
flabel comment s 6265 5614 6265 5614 3 FreeSans 200 270 0 0 sel_vcc_io_0p4
flabel comment s 911 4141 911 4141 0 FreeSans 200 0 0 0 vcc_a
flabel metal1 s 0 2486 34 2688 0 FreeSans 200 0 0 0 vgnd_io
port 2 nsew
flabel metal1 s 0 1695 34 1813 0 FreeSans 200 0 0 0 vpb
port 3 nsew
flabel metal1 s 185 1841 219 2043 0 FreeSans 200 0 0 0 vpwr
port 4 nsew
flabel metal2 s 8171 5600 8339 5638 3 FreeSans 200 270 0 0 vgnd_io
port 2 nsew
flabel metal2 s 7151 5608 7327 5638 3 FreeSans 200 270 0 0 vgnd_io
port 2 nsew
flabel metal2 s 7463 5600 7515 5638 3 FreeSans 200 270 0 0 ls_in_h
port 5 nsew
flabel metal2 s 7899 5599 8083 5638 3 FreeSans 200 270 0 0 vpwr_ka
port 6 nsew
flabel metal2 s 8417 5600 8563 5638 3 FreeSans 200 270 0 0 vcc_a
port 7 nsew
flabel metal2 s 3346 4001 3496 4021 3 FreeSans 200 270 0 0 vcc_io
port 8 nsew
flabel metal2 s 1007 4136 1323 4162 3 FreeSans 200 270 0 0 vcc_io
port 8 nsew
flabel metal2 s 6471 -50 6791 -28 3 FreeSans 200 90 0 0 vpb
port 3 nsew
flabel metal2 s 6147 -50 6415 -28 3 FreeSans 200 90 0 0 vgnd_io
port 2 nsew
flabel metal2 s 5176 -50 5547 -28 3 FreeSans 200 90 0 0 vgnd_io
port 2 nsew
flabel metal2 s 4109 -50 4234 -28 3 FreeSans 200 90 0 0 vgnd_io
port 2 nsew
flabel metal2 s 2143 -50 2345 -28 3 FreeSans 200 90 0 0 vgnd_io
port 2 nsew
flabel metal2 s -197 -50 31 -28 3 FreeSans 200 90 0 0 vgnd_io
port 2 nsew
flabel metal2 s -197 4136 185 4162 3 FreeSans 200 270 0 0 vgnd_io
port 2 nsew
flabel metal2 s 2143 4001 2345 4021 3 FreeSans 200 270 0 0 vgnd_io
port 2 nsew
flabel metal2 s 2790 3991 3152 4021 3 FreeSans 200 270 0 0 vpwr
port 4 nsew
flabel metal2 s 5175 4001 5547 4021 3 FreeSans 200 270 0 0 vgnd_io
port 2 nsew
flabel metal2 s 6147 5600 6215 5638 3 FreeSans 200 270 0 0 vgnd_io
port 2 nsew
flabel metal2 s 6799 5608 6851 5638 3 FreeSans 200 270 0 0 biasen_n
port 9 nsew
flabel metal2 s 6471 5600 6648 5638 3 FreeSans 200 270 0 0 vpb
port 3 nsew
flabel metal2 s 6323 5600 6415 5638 3 FreeSans 200 270 0 0 vgnd_io
port 2 nsew
flabel metal2 s 7071 5608 7123 5638 3 FreeSans 200 270 0 0 ls_in_h_n
port 10 nsew
flabel metal2 s 7543 5600 7711 5638 3 FreeSans 200 270 0 0 vgnd_io
port 2 nsew
flabel metal2 s 215 -94 267 -74 2 FreeSans 200 90 0 0 od_h
port 11 nsew
flabel metal2 s 490 -94 542 -74 3 FreeSans 200 90 0 0 hld_h_n
port 12 nsew
flabel metal2 s 2632 3991 2684 4021 0 FreeSans 200 0 0 0 ibuf_sel_h
port 13 nsew
flabel metal2 s 2373 3987 2425 4021 0 FreeSans 200 0 0 0 ibuf_sel_h_n
port 14 nsew
flabel metal2 s 5648 3991 5700 4021 0 FreeSans 200 0 0 0 vref_sel_h
port 15 nsew
flabel metal2 s 5884 3987 5936 4021 0 FreeSans 200 0 0 0 vref_sel_h_n
port 16 nsew
flabel metal2 s 6912 5608 6964 5638 0 FreeSans 200 0 0 0 vreg_en_h
port 17 nsew
flabel metal2 s 6676 5608 6728 5638 0 FreeSans 200 0 0 0 vreg_en_h_n
port 18 nsew
flabel metal2 s 1444 3995 1496 4021 0 FreeSans 200 0 0 0 vtrip_sel_h
port 19 nsew
flabel metal2 s 1700 3995 1752 4021 0 FreeSans 200 0 0 0 vtrip_sel_h_n
port 20 nsew
flabel metal2 s 4029 -94 4081 -74 3 FreeSans 200 90 0 0 ibuf_sel
port 21 nsew
flabel metal2 s 4262 -94 4314 -74 3 FreeSans 200 90 0 0 vref_sel
port 22 nsew
flabel metal2 s 8459 -94 8511 -74 3 FreeSans 200 90 0 0 vreg_en
port 23 nsew
flabel metal2 s 59 -94 111 -74 3 FreeSans 200 90 0 0 vtrip_sel
port 24 nsew
<< properties >>
string GDS_END 79823946
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 79759312
string path 53.575 88.550 58.625 88.550 
<< end >>
