magic
tech sky130B
magscale 1 2
timestamp 1707688321
<< obsli1 >>
rect 140 287 682 303
rect 140 253 142 287
rect 176 253 214 287
rect 248 253 286 287
rect 320 253 358 287
rect 392 253 430 287
rect 464 253 502 287
rect 536 253 574 287
rect 608 253 646 287
rect 680 253 682 287
rect 140 235 682 253
rect 50 173 84 189
rect 50 101 84 139
rect 50 51 84 67
rect 136 51 170 189
rect 222 173 256 189
rect 222 101 256 139
rect 222 51 256 67
rect 308 51 342 189
rect 394 173 428 189
rect 394 101 428 139
rect 394 51 428 67
rect 480 51 514 189
rect 566 173 600 189
rect 566 101 600 139
rect 566 51 600 67
rect 652 51 686 189
rect 738 173 772 189
rect 738 101 772 139
rect 738 51 772 67
<< obsli1c >>
rect 142 253 176 287
rect 214 253 248 287
rect 286 253 320 287
rect 358 253 392 287
rect 430 253 464 287
rect 502 253 536 287
rect 574 253 608 287
rect 646 253 680 287
rect 50 139 84 173
rect 50 67 84 101
rect 222 139 256 173
rect 222 67 256 101
rect 394 139 428 173
rect 394 67 428 101
rect 566 139 600 173
rect 566 67 600 101
rect 738 139 772 173
rect 738 67 772 101
<< metal1 >>
rect 130 287 692 299
rect 130 253 142 287
rect 176 253 214 287
rect 248 253 286 287
rect 320 253 358 287
rect 392 253 430 287
rect 464 253 502 287
rect 536 253 574 287
rect 608 253 646 287
rect 680 253 692 287
rect 130 241 692 253
rect 44 173 90 189
rect 44 139 50 173
rect 84 139 90 173
rect 44 101 90 139
rect 44 67 50 101
rect 84 67 90 101
rect 44 -29 90 67
rect 216 173 262 189
rect 216 139 222 173
rect 256 139 262 173
rect 216 101 262 139
rect 216 67 222 101
rect 256 67 262 101
rect 216 -29 262 67
rect 388 173 434 189
rect 388 139 394 173
rect 428 139 434 173
rect 388 101 434 139
rect 388 67 394 101
rect 428 67 434 101
rect 388 -29 434 67
rect 560 173 606 189
rect 560 139 566 173
rect 600 139 606 173
rect 560 101 606 139
rect 560 67 566 101
rect 600 67 606 101
rect 560 -29 606 67
rect 732 173 778 189
rect 732 139 738 173
rect 772 139 778 173
rect 732 101 778 139
rect 732 67 738 101
rect 772 67 778 101
rect 732 -29 778 67
rect 44 -89 778 -29
<< obsm1 >>
rect 127 51 179 189
rect 299 51 351 189
rect 471 51 523 189
rect 643 51 695 189
<< obsm2 >>
rect 120 43 186 197
rect 292 43 358 197
rect 464 43 530 197
rect 636 43 702 197
<< metal3 >>
rect 120 131 702 197
rect 120 43 186 131
rect 292 43 358 131
rect 464 43 530 131
rect 636 43 702 131
<< labels >>
rlabel metal3 s 636 43 702 131 6 DRAIN
port 1 nsew
rlabel metal3 s 464 43 530 131 6 DRAIN
port 1 nsew
rlabel metal3 s 292 43 358 131 6 DRAIN
port 1 nsew
rlabel metal3 s 120 131 702 197 6 DRAIN
port 1 nsew
rlabel metal3 s 120 43 186 131 6 DRAIN
port 1 nsew
rlabel metal1 s 130 241 692 299 6 GATE
port 2 nsew
rlabel metal1 s 732 -29 778 189 6 SOURCE
port 3 nsew
rlabel metal1 s 560 -29 606 189 6 SOURCE
port 3 nsew
rlabel metal1 s 388 -29 434 189 6 SOURCE
port 3 nsew
rlabel metal1 s 216 -29 262 189 6 SOURCE
port 3 nsew
rlabel metal1 s 44 -29 90 189 6 SOURCE
port 3 nsew
rlabel metal1 s 44 -89 778 -29 8 SOURCE
port 3 nsew
<< properties >>
string FIXED_BBOX 0 -89 816 303
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 9214434
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_pr/gds/sky130_fd_pr.gds
string GDS_START 9202506
<< end >>
