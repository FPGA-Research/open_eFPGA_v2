magic
tech sky130A
timestamp 1707688321
<< properties >>
string GDS_END 98003654
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 98002950
<< end >>
