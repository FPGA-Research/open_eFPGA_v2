magic
tech sky130B
magscale 1 2
timestamp 1707688321
<< nwell >>
rect 0 487 95 5063
rect 6352 3344 8395 3346
rect 5603 3254 8395 3344
rect 5438 3088 12253 3254
rect 5438 3027 11329 3088
rect 5439 2933 5605 3027
rect 4097 554 4263 1623
rect 4097 383 4275 554
<< pwell >>
rect 10979 1374 11927 1732
rect 10979 1312 11827 1374
rect 14084 149 14170 801
rect 14010 63 14170 149
<< pdiff >>
rect 6682 1314 6702 1732
rect 11873 82 11893 116
rect 11954 82 11960 116
<< psubdiff >>
rect 11005 1672 11093 1706
rect 11127 1672 11162 1706
rect 11196 1672 11231 1706
rect 11005 1638 11231 1672
rect 11005 1604 11093 1638
rect 11127 1604 11162 1638
rect 11196 1604 11231 1638
rect 11005 1570 11231 1604
rect 11005 1536 11093 1570
rect 11127 1536 11162 1570
rect 11196 1536 11231 1570
rect 11005 1502 11231 1536
rect 11005 1468 11093 1502
rect 11127 1468 11162 1502
rect 11196 1468 11231 1502
rect 11005 1434 11231 1468
rect 11005 1400 11093 1434
rect 11127 1400 11162 1434
rect 11196 1400 11231 1434
rect 11877 1400 11901 1706
rect 11005 1338 11801 1400
<< mvpsubdiff >>
rect 14110 751 14144 775
rect 14110 675 14144 717
rect 14110 599 14144 641
rect 14110 523 14144 565
rect 14110 447 14144 489
rect 14110 372 14144 413
rect 14110 297 14144 338
rect 14110 222 14144 263
rect 14110 147 14144 188
rect 14036 113 14110 123
rect 14036 89 14144 113
<< mvnsubdiff >>
rect 5669 3244 5693 3278
rect 5727 3244 5762 3278
rect 5796 3244 5831 3278
rect 5865 3244 5900 3278
rect 5934 3244 5969 3278
rect 6003 3244 6038 3278
rect 6072 3244 6106 3278
rect 6140 3244 6174 3278
rect 6208 3244 6242 3278
rect 6276 3244 6300 3278
rect 6474 3246 6498 3280
rect 6532 3246 6568 3280
rect 6602 3246 6638 3280
rect 6672 3246 6708 3280
rect 6742 3246 6778 3280
rect 6812 3246 6848 3280
rect 6882 3246 6918 3280
rect 6952 3246 6987 3280
rect 7021 3246 7056 3280
rect 7090 3246 7114 3280
rect 7288 3246 7312 3280
rect 7346 3246 7380 3280
rect 7414 3246 7448 3280
rect 7482 3246 7516 3280
rect 7550 3246 7584 3280
rect 7618 3246 7652 3280
rect 7686 3246 7720 3280
rect 7754 3246 7788 3280
rect 7822 3246 7857 3280
rect 7891 3246 7926 3280
rect 7960 3246 7995 3280
rect 8029 3246 8064 3280
rect 8098 3246 8133 3280
rect 8167 3246 8202 3280
rect 8236 3246 8271 3280
rect 8305 3246 8329 3280
rect 5504 3154 5529 3188
rect 5563 3154 5604 3188
rect 5638 3154 5860 3188
rect 5894 3154 5937 3188
rect 5971 3154 6014 3188
rect 6048 3154 6090 3188
rect 6124 3154 6166 3188
rect 6200 3154 6242 3188
rect 6276 3154 6498 3188
rect 6532 3154 6568 3188
rect 6602 3154 6638 3188
rect 6672 3154 6708 3188
rect 6742 3154 6778 3188
rect 6812 3154 6848 3188
rect 6882 3154 6918 3188
rect 6952 3154 6987 3188
rect 7021 3154 7056 3188
rect 7090 3154 7312 3188
rect 7346 3154 7384 3188
rect 7418 3154 7455 3188
rect 7489 3154 7526 3188
rect 7560 3154 7597 3188
rect 7631 3154 7668 3188
rect 7702 3154 7739 3188
rect 7773 3154 7810 3188
rect 7844 3154 7881 3188
rect 7915 3154 7952 3188
rect 7986 3154 8023 3188
rect 8057 3154 8094 3188
rect 8128 3154 8165 3188
rect 8199 3154 8236 3188
rect 8270 3154 8307 3188
rect 8341 3154 8378 3188
rect 8412 3154 8449 3188
rect 8483 3154 8520 3188
rect 8554 3154 8591 3188
rect 8625 3154 8662 3188
rect 8696 3154 8733 3188
rect 8767 3154 8804 3188
rect 8838 3154 9112 3188
rect 9146 3154 9185 3188
rect 9219 3154 9258 3188
rect 9292 3154 9510 3188
rect 9544 3154 9578 3188
rect 9612 3154 9646 3188
rect 9680 3154 9714 3188
rect 9748 3154 9783 3188
rect 9817 3154 9852 3188
rect 9886 3154 9921 3188
rect 9955 3154 9990 3188
rect 10024 3154 10059 3188
rect 10093 3154 10128 3188
rect 10162 3154 10197 3188
rect 10231 3154 10266 3188
rect 10300 3154 10335 3188
rect 10369 3154 10404 3188
rect 10438 3154 10473 3188
rect 10507 3154 10542 3188
rect 10576 3154 10611 3188
rect 10645 3154 10680 3188
rect 10714 3154 10749 3188
rect 10783 3154 10818 3188
rect 10852 3154 10887 3188
rect 10921 3154 10956 3188
rect 10990 3154 11025 3188
rect 11059 3154 11094 3188
rect 11128 3154 11163 3188
rect 11197 3154 11232 3188
rect 11266 3154 11301 3188
rect 11335 3154 11370 3188
rect 11404 3154 11439 3188
rect 11473 3154 11508 3188
rect 11542 3154 11577 3188
rect 11611 3154 11646 3188
rect 11680 3154 11715 3188
rect 11749 3154 11784 3188
rect 11818 3154 11853 3188
rect 11887 3154 11922 3188
rect 11956 3154 11991 3188
rect 12025 3154 12060 3188
rect 12094 3154 12129 3188
rect 12163 3154 12187 3188
rect 5504 3057 5540 3154
rect 5504 3023 5505 3057
rect 5539 3023 5540 3057
rect 11393 3031 12187 3154
rect 5504 3016 5540 3023
rect 5505 2999 5539 3016
rect 4163 1533 4197 1557
rect 4163 1461 4197 1499
rect 4163 1389 4197 1427
rect 4163 1317 4197 1355
rect 4163 1245 4197 1283
rect 4163 1173 4197 1211
rect 4163 1101 4197 1139
rect 4163 1029 4197 1067
rect 4163 957 4197 995
rect 4163 885 4197 923
rect 4163 813 4197 851
rect 4163 741 4197 779
rect 4163 669 4197 707
rect 4163 598 4197 635
rect 4163 527 4197 564
rect 4163 483 4197 493
rect 4163 449 4280 483
<< psubdiffcont >>
rect 11093 1672 11127 1706
rect 11162 1672 11196 1706
rect 11093 1604 11127 1638
rect 11162 1604 11196 1638
rect 11093 1536 11127 1570
rect 11162 1536 11196 1570
rect 11093 1468 11127 1502
rect 11162 1468 11196 1502
rect 11093 1400 11127 1434
rect 11162 1400 11196 1434
rect 11231 1400 11877 1706
<< mvpsubdiffcont >>
rect 14110 717 14144 751
rect 14110 641 14144 675
rect 14110 565 14144 599
rect 14110 489 14144 523
rect 14110 413 14144 447
rect 14110 338 14144 372
rect 14110 263 14144 297
rect 14110 188 14144 222
rect 14110 113 14144 147
<< mvnsubdiffcont >>
rect 5693 3244 5727 3278
rect 5762 3244 5796 3278
rect 5831 3244 5865 3278
rect 5900 3244 5934 3278
rect 5969 3244 6003 3278
rect 6038 3244 6072 3278
rect 6106 3244 6140 3278
rect 6174 3244 6208 3278
rect 6242 3244 6276 3278
rect 6498 3246 6532 3280
rect 6568 3246 6602 3280
rect 6638 3246 6672 3280
rect 6708 3246 6742 3280
rect 6778 3246 6812 3280
rect 6848 3246 6882 3280
rect 6918 3246 6952 3280
rect 6987 3246 7021 3280
rect 7056 3246 7090 3280
rect 7312 3246 7346 3280
rect 7380 3246 7414 3280
rect 7448 3246 7482 3280
rect 7516 3246 7550 3280
rect 7584 3246 7618 3280
rect 7652 3246 7686 3280
rect 7720 3246 7754 3280
rect 7788 3246 7822 3280
rect 7857 3246 7891 3280
rect 7926 3246 7960 3280
rect 7995 3246 8029 3280
rect 8064 3246 8098 3280
rect 8133 3246 8167 3280
rect 8202 3246 8236 3280
rect 8271 3246 8305 3280
rect 5529 3154 5563 3188
rect 5604 3154 5638 3188
rect 5860 3154 5894 3188
rect 5937 3154 5971 3188
rect 6014 3154 6048 3188
rect 6090 3154 6124 3188
rect 6166 3154 6200 3188
rect 6242 3154 6276 3188
rect 6498 3154 6532 3188
rect 6568 3154 6602 3188
rect 6638 3154 6672 3188
rect 6708 3154 6742 3188
rect 6778 3154 6812 3188
rect 6848 3154 6882 3188
rect 6918 3154 6952 3188
rect 6987 3154 7021 3188
rect 7056 3154 7090 3188
rect 7312 3154 7346 3188
rect 7384 3154 7418 3188
rect 7455 3154 7489 3188
rect 7526 3154 7560 3188
rect 7597 3154 7631 3188
rect 7668 3154 7702 3188
rect 7739 3154 7773 3188
rect 7810 3154 7844 3188
rect 7881 3154 7915 3188
rect 7952 3154 7986 3188
rect 8023 3154 8057 3188
rect 8094 3154 8128 3188
rect 8165 3154 8199 3188
rect 8236 3154 8270 3188
rect 8307 3154 8341 3188
rect 8378 3154 8412 3188
rect 8449 3154 8483 3188
rect 8520 3154 8554 3188
rect 8591 3154 8625 3188
rect 8662 3154 8696 3188
rect 8733 3154 8767 3188
rect 8804 3154 8838 3188
rect 9112 3154 9146 3188
rect 9185 3154 9219 3188
rect 9258 3154 9292 3188
rect 9510 3154 9544 3188
rect 9578 3154 9612 3188
rect 9646 3154 9680 3188
rect 9714 3154 9748 3188
rect 9783 3154 9817 3188
rect 9852 3154 9886 3188
rect 9921 3154 9955 3188
rect 9990 3154 10024 3188
rect 10059 3154 10093 3188
rect 10128 3154 10162 3188
rect 10197 3154 10231 3188
rect 10266 3154 10300 3188
rect 10335 3154 10369 3188
rect 10404 3154 10438 3188
rect 10473 3154 10507 3188
rect 10542 3154 10576 3188
rect 10611 3154 10645 3188
rect 10680 3154 10714 3188
rect 10749 3154 10783 3188
rect 10818 3154 10852 3188
rect 10887 3154 10921 3188
rect 10956 3154 10990 3188
rect 11025 3154 11059 3188
rect 11094 3154 11128 3188
rect 11163 3154 11197 3188
rect 11232 3154 11266 3188
rect 11301 3154 11335 3188
rect 11370 3154 11404 3188
rect 11439 3154 11473 3188
rect 11508 3154 11542 3188
rect 11577 3154 11611 3188
rect 11646 3154 11680 3188
rect 11715 3154 11749 3188
rect 11784 3154 11818 3188
rect 11853 3154 11887 3188
rect 11922 3154 11956 3188
rect 11991 3154 12025 3188
rect 12060 3154 12094 3188
rect 12129 3154 12163 3188
rect 5505 3023 5539 3057
rect 4163 1499 4197 1533
rect 4163 1427 4197 1461
rect 4163 1355 4197 1389
rect 4163 1283 4197 1317
rect 4163 1211 4197 1245
rect 4163 1139 4197 1173
rect 4163 1067 4197 1101
rect 4163 995 4197 1029
rect 4163 923 4197 957
rect 4163 851 4197 885
rect 4163 779 4197 813
rect 4163 707 4197 741
rect 4163 635 4197 669
rect 4163 564 4197 598
rect 4163 493 4197 527
<< locali >>
rect 7920 4137 7959 4171
rect 7993 4137 8032 4171
rect 8066 4137 8106 4171
rect 6581 3335 7807 3446
rect 6474 3330 7807 3335
rect 6474 3322 8329 3330
rect 6474 3280 7114 3322
rect 7288 3280 8329 3322
rect 5505 3244 5693 3278
rect 5727 3244 5762 3278
rect 5796 3244 5831 3278
rect 5865 3244 5900 3278
rect 5934 3244 5969 3278
rect 6003 3244 6038 3278
rect 6072 3244 6106 3278
rect 6140 3244 6174 3278
rect 6208 3244 6242 3278
rect 6276 3244 6300 3278
rect 5505 3234 6300 3244
rect 5505 3188 5662 3234
rect 5505 3154 5529 3188
rect 5563 3154 5604 3188
rect 5638 3154 5662 3188
rect 5730 3166 5768 3200
rect 5505 3057 5539 3154
rect 5696 3048 5802 3166
rect 5836 3188 6300 3234
rect 5836 3154 5860 3188
rect 5894 3154 5937 3188
rect 5971 3154 6014 3188
rect 6048 3154 6090 3188
rect 6124 3154 6166 3188
rect 6200 3154 6242 3188
rect 6276 3154 6300 3188
rect 6368 3246 6406 3280
rect 6119 3039 6152 3060
rect 6334 3048 6440 3246
rect 6474 3246 6498 3280
rect 6532 3246 6568 3280
rect 6602 3246 6638 3280
rect 6672 3246 6708 3280
rect 6742 3246 6778 3280
rect 6812 3246 6848 3280
rect 6882 3246 6918 3280
rect 6952 3246 6987 3280
rect 7021 3246 7056 3280
rect 7090 3246 7114 3280
rect 6474 3188 7114 3246
rect 6474 3154 6498 3188
rect 6532 3154 6568 3188
rect 6602 3154 6638 3188
rect 6672 3154 6708 3188
rect 6742 3154 6778 3188
rect 6812 3154 6848 3188
rect 6882 3154 6918 3188
rect 6952 3154 6987 3188
rect 7021 3154 7056 3188
rect 7090 3154 7114 3188
rect 7182 3246 7220 3280
rect 7148 3048 7254 3246
rect 7288 3246 7312 3280
rect 7346 3246 7380 3280
rect 7414 3246 7448 3280
rect 7482 3246 7516 3280
rect 7550 3246 7584 3280
rect 7618 3246 7652 3280
rect 7686 3246 7720 3280
rect 7754 3246 7788 3280
rect 7822 3246 7857 3280
rect 7891 3246 7926 3280
rect 7960 3246 7995 3280
rect 8029 3246 8064 3280
rect 8098 3246 8133 3280
rect 8167 3246 8202 3280
rect 8236 3246 8271 3280
rect 8305 3246 8329 3280
rect 7288 3188 8329 3246
rect 8983 3321 9021 3355
rect 8600 3188 8638 3206
rect 8672 3188 8710 3206
rect 7288 3154 7312 3188
rect 7346 3154 7384 3188
rect 7418 3154 7455 3188
rect 7489 3154 7526 3188
rect 7560 3154 7597 3188
rect 7631 3154 7668 3188
rect 7702 3154 7739 3188
rect 7773 3154 7810 3188
rect 7844 3154 7881 3188
rect 7915 3154 7952 3188
rect 7986 3154 8023 3188
rect 8057 3154 8094 3188
rect 8128 3154 8165 3188
rect 8199 3154 8236 3188
rect 8270 3154 8307 3188
rect 8341 3154 8378 3188
rect 8412 3154 8449 3188
rect 8483 3154 8520 3188
rect 8554 3172 8566 3188
rect 8625 3172 8638 3188
rect 8696 3172 8710 3188
rect 8554 3154 8591 3172
rect 8625 3154 8662 3172
rect 8696 3154 8733 3172
rect 8767 3154 8804 3188
rect 8838 3154 8862 3188
rect 7644 3086 7682 3120
rect 7820 3086 7858 3120
rect 8458 3086 8496 3120
rect 8949 3114 9030 3321
rect 9350 3239 9351 3273
rect 9385 3239 9423 3273
rect 9137 3188 9175 3200
rect 9209 3188 9247 3200
rect 9088 3166 9103 3188
rect 9146 3166 9175 3188
rect 9219 3166 9247 3188
rect 9088 3154 9112 3166
rect 9146 3154 9185 3166
rect 9219 3154 9258 3166
rect 9292 3154 9316 3188
rect 9350 3114 9452 3239
rect 9486 3154 9510 3188
rect 9544 3154 9578 3188
rect 9612 3154 9646 3188
rect 9680 3154 9714 3188
rect 9748 3154 9783 3188
rect 9817 3154 9852 3188
rect 9886 3154 9921 3188
rect 9955 3154 9990 3188
rect 10024 3154 10059 3188
rect 10093 3154 10128 3188
rect 10162 3154 10197 3188
rect 10231 3154 10266 3188
rect 10300 3154 10335 3188
rect 10369 3154 10404 3188
rect 10438 3154 10473 3188
rect 10507 3154 10542 3188
rect 10576 3154 10611 3188
rect 10645 3154 10680 3188
rect 10714 3154 10749 3188
rect 10783 3154 10818 3188
rect 10852 3154 10887 3188
rect 10921 3154 10956 3188
rect 10990 3154 11025 3188
rect 11059 3154 11094 3188
rect 11128 3154 11163 3188
rect 11197 3154 11232 3188
rect 11266 3154 11301 3188
rect 11335 3154 11370 3188
rect 11404 3154 11439 3188
rect 11473 3154 11508 3188
rect 11542 3154 11577 3188
rect 11611 3154 11646 3188
rect 11680 3154 11715 3188
rect 11749 3154 11784 3188
rect 11818 3154 11853 3188
rect 11887 3154 11922 3188
rect 11956 3154 11991 3188
rect 12025 3154 12060 3188
rect 12094 3154 12129 3188
rect 12163 3154 12187 3188
rect 8880 3049 9030 3114
rect 9558 3086 9596 3120
rect 10834 3086 10872 3120
rect 11010 3086 11048 3120
rect 5505 2999 5539 3023
rect 6098 3005 6136 3039
rect 11393 3027 12187 3154
rect 5644 2828 5678 2866
rect 4395 2247 4429 2383
rect 4707 2247 4741 2383
rect 5820 2076 5854 2113
rect 6634 2076 6668 2113
rect 7096 2076 7130 2113
rect 7910 2076 7944 2113
rect 8548 2076 8582 2113
rect 9186 2076 9220 2122
rect 9648 2076 9682 2122
rect 10286 2076 10320 2122
rect 10748 2076 10782 2122
rect 4289 1718 4327 1752
rect 4977 1718 5015 1752
rect 4551 1586 4585 1624
rect 4163 1533 4197 1557
rect 4659 1570 4713 1605
rect 5083 1572 5187 1739
rect 4163 1461 4197 1499
rect 4693 1536 4713 1570
rect 5115 1538 5153 1572
rect 4659 1498 4713 1536
rect 4693 1464 4713 1498
rect 4163 1389 4197 1427
rect 4163 1317 4197 1355
rect 5705 1418 5759 1605
rect 5705 1384 5725 1418
rect 5705 1346 5759 1384
rect 5705 1312 5725 1346
rect 4163 1245 4197 1283
rect 4163 1173 4197 1211
rect 4163 1101 4197 1139
rect 4163 1029 4197 1067
rect 4163 957 4197 995
rect 4163 885 4197 923
rect 4163 813 4197 851
rect 4163 741 4197 779
rect 4163 669 4197 707
rect 4163 598 4197 635
rect 4163 527 4197 564
rect 4163 483 4197 493
rect 5936 1247 6082 1732
rect 10990 1706 11028 1732
rect 11325 1706 12223 1798
rect 10990 1698 11093 1706
rect 10998 1672 11093 1698
rect 11127 1672 11162 1706
rect 11196 1672 11231 1706
rect 8618 1424 8724 1664
rect 8652 1390 8690 1424
rect 8618 1389 8724 1390
rect 10998 1638 11231 1672
rect 10998 1604 11093 1638
rect 11127 1604 11162 1638
rect 11196 1604 11231 1638
rect 10998 1570 11231 1604
rect 10998 1536 11093 1570
rect 11127 1536 11162 1570
rect 11196 1536 11231 1570
rect 10998 1502 11231 1536
rect 10998 1468 11093 1502
rect 11127 1468 11162 1502
rect 11196 1468 11231 1502
rect 10998 1434 11231 1468
rect 10998 1400 11093 1434
rect 11127 1400 11162 1434
rect 11196 1400 11231 1434
rect 11877 1475 12223 1706
rect 13668 1492 13706 1526
rect 11877 1400 11901 1475
rect 10998 1345 11793 1400
rect 6361 1280 6395 1314
rect 8007 1280 8041 1314
rect 9653 1280 9687 1314
rect 11299 1280 11333 1314
rect 11483 1280 11517 1314
rect 11667 1280 11701 1314
rect 5936 1141 6057 1247
rect 5936 826 6082 1141
rect 7751 1052 7785 1086
rect 9397 984 9431 1022
rect 9907 1019 9945 1053
rect 11041 1022 11079 1056
rect 13149 1020 13183 1094
rect 13501 1020 13535 1090
rect 13149 986 13275 1020
rect 6042 720 6082 826
rect 4163 449 4281 483
rect 5936 449 6082 720
rect 7853 848 7891 882
rect 7819 574 7925 848
rect 14110 751 14144 775
rect 14110 675 14144 717
rect 14110 599 14144 641
rect 6651 540 6689 574
rect 7853 540 7891 574
rect 8261 544 8299 578
rect 11694 535 11702 569
rect 11736 535 11748 569
rect 11694 497 11748 535
rect 11694 463 11702 497
rect 11736 463 11748 497
rect 11535 281 11573 315
rect 11694 188 11748 463
rect 14110 523 14144 565
rect 14110 447 14144 489
rect 14110 372 14144 413
rect 14110 297 14144 338
rect 14110 222 14144 263
rect 14110 147 14144 188
rect 14036 113 14110 123
rect 14036 89 14144 113
<< viali >>
rect 7886 4137 7920 4171
rect 7959 4137 7993 4171
rect 8032 4137 8066 4171
rect 8106 4137 8140 4171
rect 5696 3166 5730 3200
rect 5768 3166 5802 3200
rect 6334 3246 6368 3280
rect 6406 3246 6440 3280
rect 7148 3246 7182 3280
rect 7220 3246 7254 3280
rect 8949 3321 8983 3355
rect 9021 3321 9055 3355
rect 8566 3188 8600 3206
rect 8638 3188 8672 3206
rect 8710 3188 8744 3206
rect 8566 3172 8591 3188
rect 8591 3172 8600 3188
rect 8638 3172 8662 3188
rect 8662 3172 8672 3188
rect 8710 3172 8733 3188
rect 8733 3172 8744 3188
rect 7610 3086 7644 3120
rect 7682 3086 7716 3120
rect 7786 3086 7820 3120
rect 7858 3086 7892 3120
rect 8424 3086 8458 3120
rect 8496 3086 8530 3120
rect 9351 3239 9385 3273
rect 9423 3239 9457 3273
rect 9103 3188 9137 3200
rect 9175 3188 9209 3200
rect 9247 3188 9281 3200
rect 9103 3166 9112 3188
rect 9112 3166 9137 3188
rect 9175 3166 9185 3188
rect 9185 3166 9209 3188
rect 9247 3166 9258 3188
rect 9258 3166 9281 3188
rect 9524 3086 9558 3120
rect 9596 3086 9630 3120
rect 10800 3086 10834 3120
rect 10872 3086 10906 3120
rect 10976 3086 11010 3120
rect 11048 3086 11082 3120
rect 6064 3005 6098 3039
rect 6136 3005 6170 3039
rect 5644 2866 5678 2900
rect 5644 2794 5678 2828
rect 4255 1718 4289 1752
rect 4327 1718 4361 1752
rect 4943 1718 4977 1752
rect 5015 1718 5049 1752
rect 4551 1624 4585 1658
rect 4551 1552 4585 1586
rect 4659 1536 4693 1570
rect 5081 1538 5115 1572
rect 5153 1538 5187 1572
rect 4659 1464 4693 1498
rect 5725 1384 5759 1418
rect 5725 1312 5759 1346
rect 8618 1390 8652 1424
rect 8690 1390 8724 1424
rect 13634 1492 13668 1526
rect 13706 1492 13740 1526
rect 6057 1141 6163 1247
rect 9397 1022 9431 1056
rect 9873 1019 9907 1053
rect 9945 1019 9979 1053
rect 11007 1022 11041 1056
rect 11079 1022 11113 1056
rect 9397 950 9431 984
rect 5936 720 6042 826
rect 7819 848 7853 882
rect 7891 848 7925 882
rect 6617 540 6651 574
rect 6689 540 6723 574
rect 7819 540 7853 574
rect 7891 540 7925 574
rect 8227 544 8261 578
rect 8299 544 8333 578
rect 11702 535 11736 569
rect 11702 463 11736 497
rect 11501 281 11535 315
rect 11573 281 11607 315
<< metal1 >>
tri 6809 5301 6847 5339 se
rect 6847 5333 6899 5339
rect 4633 5295 6847 5301
rect 4685 5281 6847 5295
rect 4685 5269 6899 5281
rect 4685 5249 6847 5269
rect 4685 5243 4700 5249
rect 4633 5231 4700 5243
rect 4685 5211 4700 5231
tri 4700 5211 4738 5249 nw
tri 6809 5211 6847 5249 ne
rect 6847 5211 6899 5217
tri 4685 5196 4700 5211 nw
rect 4633 5173 4685 5179
rect 1680 5153 1732 5159
rect 1680 5089 1732 5101
tri 1732 5080 1757 5105 sw
rect 5354 5090 5540 5096
rect 1732 5037 3585 5080
rect 1680 5028 3585 5037
rect 3637 5028 3649 5080
rect 3701 5028 3707 5080
rect 5354 5038 5355 5090
rect 5407 5038 5421 5090
rect 5473 5038 5487 5090
rect 5539 5038 5540 5090
rect 5354 5021 5540 5038
rect 5354 4969 5355 5021
rect 5407 4969 5421 5021
rect 5473 4969 5487 5021
rect 5539 4969 5540 5021
rect 5354 4952 5540 4969
rect 5354 4900 5355 4952
rect 5407 4900 5421 4952
rect 5473 4900 5487 4952
rect 5539 4900 5540 4952
rect 5354 4883 5540 4900
rect 5354 4831 5355 4883
rect 5407 4831 5421 4883
rect 5473 4831 5487 4883
rect 5539 4831 5540 4883
rect 5354 4814 5540 4831
rect 5354 4762 5355 4814
rect 5407 4762 5421 4814
rect 5473 4762 5487 4814
rect 5539 4762 5540 4814
rect 5354 4745 5540 4762
rect 5354 4693 5355 4745
rect 5407 4693 5421 4745
rect 5473 4693 5487 4745
rect 5539 4693 5540 4745
rect 5354 4676 5540 4693
rect 5354 4624 5355 4676
rect 5407 4624 5421 4676
rect 5473 4624 5487 4676
rect 5539 4624 5540 4676
rect 6228 4977 6542 4983
rect 6228 4669 6231 4977
rect 6539 4669 6542 4977
rect 6228 4663 6542 4669
rect 5354 4618 5540 4624
rect 6847 4392 7035 4398
rect 6899 4340 7035 4392
rect 6847 4326 7035 4340
rect 6899 4274 7035 4326
rect 6847 4268 7035 4274
tri 6979 4238 7009 4268 ne
rect 7009 4238 7035 4268
tri 11881 4238 11937 4294 se
rect 11937 4288 11989 4294
tri 7009 4212 7035 4238 ne
rect 7705 4212 8237 4238
tri 8237 4212 8263 4238 sw
tri 11855 4212 11881 4238 se
rect 11881 4236 11937 4238
rect 11881 4224 11989 4236
rect 11881 4212 11937 4224
rect 7705 4207 8263 4212
tri 8263 4207 8268 4212 sw
rect 7705 4205 8268 4207
tri 8174 4180 8199 4205 ne
rect 8199 4180 8268 4205
tri 4789 4177 4792 4180 se
rect 4792 4177 4798 4180
tri 4786 4174 4789 4177 se
rect 4789 4174 4798 4177
rect 4792 4128 4798 4174
rect 4850 4128 4862 4180
rect 4914 4177 4920 4180
tri 4920 4177 4923 4180 sw
tri 8199 4177 8202 4180 ne
rect 8202 4177 8268 4180
rect 4914 4174 4923 4177
tri 4923 4174 4926 4177 sw
rect 4914 4128 4920 4174
rect 7874 4171 8157 4177
rect 7874 4137 7886 4171
rect 7920 4137 7959 4171
rect 7993 4137 8032 4171
rect 8066 4137 8106 4171
rect 8140 4163 8157 4171
tri 8157 4163 8171 4177 sw
tri 8202 4163 8216 4177 ne
rect 8140 4146 8171 4163
tri 8171 4146 8188 4163 sw
rect 8140 4140 8188 4146
rect 7874 4131 8136 4137
tri 8058 4128 8061 4131 ne
rect 8061 4128 8136 4131
tri 8061 4091 8098 4128 ne
rect 8098 4091 8136 4128
tri 8098 4053 8136 4091 ne
rect 8136 4076 8188 4088
rect 8136 4018 8188 4024
rect 8216 4085 8268 4177
tri 11989 4212 12071 4294 sw
rect 11937 4166 11989 4172
rect 8216 4021 8268 4033
rect 8216 3963 8268 3969
rect 7000 3657 7006 3709
rect 7058 3657 7076 3709
rect 7128 3657 7146 3709
rect 7198 3657 7216 3709
rect 7268 3657 7286 3709
rect 7338 3657 7356 3709
rect 7408 3657 7426 3709
rect 7478 3657 7496 3709
rect 7548 3657 7566 3709
rect 7618 3657 7636 3709
rect 7688 3657 7705 3709
rect 7757 3657 7763 3709
rect 6862 3576 6868 3628
rect 6920 3576 6926 3628
rect 6862 3564 6926 3576
rect 6862 3512 6868 3564
rect 6920 3512 6926 3564
rect 7000 3627 7763 3657
rect 7000 3575 7006 3627
rect 7058 3575 7076 3627
rect 7128 3575 7146 3627
rect 7198 3575 7216 3627
rect 7268 3575 7286 3627
rect 7338 3575 7356 3627
rect 7408 3575 7426 3627
rect 7478 3575 7496 3627
rect 7548 3575 7566 3627
rect 7618 3575 7636 3627
rect 7688 3575 7705 3627
rect 7757 3575 7763 3627
rect 7000 3545 7763 3575
rect 7000 3493 7006 3545
rect 7058 3493 7076 3545
rect 7128 3493 7146 3545
rect 7198 3493 7216 3545
rect 7268 3493 7286 3545
rect 7338 3493 7356 3545
rect 7408 3493 7426 3545
rect 7478 3493 7496 3545
rect 7548 3493 7566 3545
rect 7618 3493 7636 3545
rect 7688 3493 7705 3545
rect 7757 3493 7763 3545
tri 9711 3493 9723 3505 se
rect 9723 3493 9729 3505
tri 9674 3456 9711 3493 se
rect 9711 3456 9729 3493
rect 9723 3453 9729 3456
rect 9781 3453 9787 3505
tri 9787 3456 9836 3505 sw
rect 9723 3441 9787 3453
tri 9702 3389 9723 3410 ne
rect 9723 3389 9729 3441
rect 9781 3389 9787 3441
tri 9787 3389 9808 3410 nw
rect 8318 3356 8648 3358
tri 8648 3356 8650 3358 sw
tri 6559 3286 6584 3311 se
rect 6584 3304 6590 3356
rect 6642 3304 6648 3356
rect 6584 3292 6648 3304
rect 6584 3286 6590 3292
rect 6322 3280 6590 3286
rect 6322 3246 6334 3280
rect 6368 3246 6406 3280
rect 6440 3246 6590 3280
rect 6322 3240 6590 3246
rect 6642 3240 6648 3292
rect 6676 3304 6682 3356
rect 6734 3304 6740 3356
rect 8318 3355 8650 3356
tri 8650 3355 8651 3356 sw
rect 8937 3355 12822 3361
rect 8318 3321 8651 3355
tri 8651 3321 8685 3355 sw
rect 8937 3321 8949 3355
rect 8983 3321 9021 3355
rect 9055 3321 12822 3355
rect 8318 3315 8685 3321
tri 8685 3315 8691 3321 sw
rect 6676 3292 6740 3304
rect 6676 3240 6682 3292
rect 6734 3286 6740 3292
tri 6740 3286 6765 3311 sw
rect 8318 3309 8691 3315
tri 8691 3309 8697 3315 sw
rect 8937 3309 12822 3321
rect 12874 3309 12886 3361
rect 12938 3309 12944 3361
rect 13606 3355 13658 3361
rect 8318 3286 8697 3309
tri 8697 3286 8720 3309 sw
tri 13588 3286 13606 3304 se
rect 13606 3291 13658 3303
rect 6734 3280 7266 3286
rect 6734 3246 7148 3280
rect 7182 3246 7220 3280
rect 7254 3246 7266 3280
rect 6734 3240 7266 3246
rect 8318 3279 8720 3286
tri 8720 3279 8727 3286 sw
tri 13581 3279 13588 3286 se
rect 13588 3279 13606 3286
rect 8318 3273 8727 3279
tri 8727 3273 8733 3279 sw
rect 9339 3273 13606 3279
rect 8318 3240 8733 3273
tri 8733 3240 8766 3273 sw
tri 8535 3239 8536 3240 ne
rect 8536 3239 8766 3240
tri 8766 3239 8767 3240 sw
rect 9339 3239 9351 3273
rect 9385 3239 9423 3273
rect 9457 3239 13606 3273
tri 8536 3218 8557 3239 ne
rect 8557 3233 8767 3239
tri 8767 3233 8773 3239 sw
rect 9339 3233 13658 3239
rect 8557 3218 8773 3233
tri 8773 3218 8788 3233 sw
tri 8557 3215 8560 3218 ne
rect 8560 3212 8788 3218
tri 8788 3212 8794 3218 sw
rect 3655 3202 3707 3208
rect 5684 3206 8188 3212
rect 5684 3200 8136 3206
rect 5684 3166 5696 3200
rect 5730 3166 5768 3200
rect 5802 3166 8136 3200
rect 5684 3160 8136 3166
tri 8081 3157 8084 3160 ne
rect 8084 3157 8136 3160
rect 3655 3138 3707 3150
rect 1022 3013 1028 3129
rect 1144 3013 1150 3129
rect 1950 3013 1956 3129
rect 2072 3013 2078 3129
tri 3707 3132 3732 3157 sw
tri 8084 3132 8109 3157 ne
rect 8109 3154 8136 3157
rect 8560 3206 8818 3212
rect 8560 3172 8566 3206
rect 8600 3172 8638 3206
rect 8672 3172 8710 3206
rect 8744 3172 8818 3206
rect 8560 3160 8818 3172
rect 8870 3160 8882 3212
rect 8934 3160 8946 3212
rect 8998 3160 9010 3212
rect 9062 3160 9074 3212
rect 9126 3200 9138 3212
rect 9190 3206 9320 3212
tri 9320 3206 9326 3212 sw
rect 9190 3205 9326 3206
tri 9326 3205 9327 3206 sw
rect 9190 3200 9713 3205
rect 9137 3166 9138 3200
rect 9209 3166 9247 3200
rect 9281 3166 9713 3200
rect 9126 3160 9138 3166
rect 9190 3160 9713 3166
rect 10303 3199 10611 3205
tri 9688 3159 9689 3160 ne
rect 8109 3142 8188 3154
rect 8109 3132 8136 3142
rect 3707 3126 3732 3132
tri 3732 3126 3738 3132 sw
rect 3707 3120 7728 3126
rect 3707 3086 7610 3120
rect 7644 3086 7682 3120
rect 7716 3086 7728 3120
rect 3655 3080 7728 3086
rect 7774 3120 7826 3132
rect 7878 3120 7890 3132
rect 7774 3086 7786 3120
rect 7820 3086 7826 3120
rect 7774 3080 7826 3086
rect 7878 3080 7890 3086
rect 7942 3080 8056 3132
tri 8109 3120 8121 3132 ne
rect 8121 3120 8136 3132
tri 8121 3105 8136 3120 ne
tri 10280 3141 10298 3159 ne
rect 10298 3147 10303 3159
rect 10355 3147 10367 3199
rect 10419 3147 10431 3199
rect 10483 3147 10495 3199
rect 10547 3147 10559 3199
rect 10298 3141 10611 3147
rect 10788 3199 10932 3205
rect 10788 3147 10880 3199
rect 10788 3135 10932 3147
rect 8136 3084 8188 3090
rect 8412 3120 8561 3132
rect 8412 3086 8424 3120
rect 8458 3086 8496 3120
rect 8530 3086 8561 3120
rect 8412 3080 8561 3086
rect 8613 3080 8625 3132
rect 8677 3080 8683 3132
rect 8711 3080 8717 3132
rect 8769 3080 8781 3132
rect 8833 3120 9642 3132
rect 8833 3086 9524 3120
rect 9558 3086 9596 3120
rect 9630 3086 9642 3120
rect 8833 3080 9642 3086
rect 10788 3120 10880 3135
rect 10788 3086 10800 3120
rect 10834 3086 10872 3120
rect 10788 3083 10880 3086
rect 10788 3077 10932 3083
rect 10960 3199 11094 3205
rect 11012 3147 11094 3199
rect 10960 3135 11094 3147
rect 11012 3120 11094 3135
rect 11012 3086 11048 3120
rect 11082 3086 11094 3120
rect 11012 3083 11094 3086
rect 10960 3077 11094 3083
tri 9809 3051 9833 3075 se
rect 9833 3051 9839 3075
rect 6058 3039 9839 3051
rect 6058 3005 6064 3039
rect 6098 3005 6136 3039
rect 6170 3023 9839 3039
rect 9891 3023 9903 3075
rect 9955 3023 9961 3075
rect 11411 3064 12189 3192
rect 6170 3005 6178 3023
rect 6058 2995 6178 3005
tri 6178 2995 6206 3023 nw
rect 6058 2993 6176 2995
tri 6176 2993 6178 2995 nw
rect 6734 2943 6740 2995
rect 6792 2943 6804 2995
rect 6856 2989 14318 2995
rect 6856 2962 14266 2989
rect 6856 2943 6862 2962
tri 6862 2943 6881 2962 nw
tri 14241 2943 14260 2962 ne
rect 14260 2943 14266 2962
tri 14260 2937 14266 2943 ne
rect 4872 2910 4924 2916
tri 4924 2906 4934 2916 sw
rect 4924 2900 5690 2906
rect 4924 2866 5644 2900
rect 5678 2866 5690 2900
rect 7820 2882 7826 2934
rect 7878 2882 7890 2934
rect 7942 2882 8226 2934
rect 8278 2882 8290 2934
rect 8342 2882 8348 2934
rect 8416 2881 8422 2933
rect 8474 2881 8486 2933
rect 8538 2927 14229 2933
rect 8538 2900 14177 2927
rect 8538 2881 8544 2900
tri 8544 2881 8563 2900 nw
tri 14152 2881 14171 2900 ne
rect 14171 2881 14177 2900
tri 14171 2875 14177 2881 ne
rect 4924 2858 5690 2866
rect 4872 2846 5690 2858
rect 4924 2828 5690 2846
rect 4924 2794 5644 2828
rect 5678 2794 5690 2828
rect 14177 2863 14229 2875
rect 14266 2925 14318 2937
rect 14266 2867 14318 2873
rect 14177 2805 14229 2811
rect 4872 2788 5690 2794
rect 5016 2706 5022 2758
rect 5074 2706 5080 2758
rect 5016 2694 5080 2706
rect 5016 2642 5022 2694
rect 5074 2688 5080 2694
tri 5080 2688 5105 2713 sw
tri 6509 2688 6534 2713 se
rect 5074 2642 6576 2688
rect 5424 2608 5540 2614
rect 2967 2415 2973 2595
rect 3089 2415 3095 2595
rect 5476 2556 5488 2608
rect 3981 2424 5143 2552
rect 5424 2538 5540 2556
rect 5476 2486 5488 2538
rect 5424 2467 5540 2486
rect 3981 2387 5025 2424
tri 5025 2387 5062 2424 nw
rect 5476 2415 5488 2467
rect 5424 2396 5540 2415
rect 3981 2088 4345 2387
rect 5476 2344 5488 2396
rect 5424 2338 5540 2344
tri 5025 2244 5050 2269 sw
rect 5025 2234 5050 2244
tri 5050 2234 5060 2244 sw
rect 6897 2238 6949 2244
tri 4345 2136 4363 2154 nw
tri 4949 2136 4967 2154 ne
rect 5025 2116 5493 2234
tri 6872 2162 6897 2187 se
rect 6897 2174 6949 2186
tri 6949 2162 6974 2187 sw
tri 9774 2162 9799 2187 se
rect 9799 2180 9805 2232
rect 9857 2180 9863 2232
rect 9799 2168 9863 2180
tri 9863 2168 9882 2187 sw
rect 6897 2116 6949 2122
rect 9799 2116 9805 2168
rect 9857 2162 9882 2168
tri 9882 2162 9888 2168 sw
tri 10450 2162 10456 2168 se
rect 9857 2116 9863 2162
rect 10456 2116 10462 2168
rect 10514 2116 10526 2168
rect 10578 2116 10584 2168
tri 10584 2162 10590 2168 sw
tri 4345 2088 4358 2101 sw
tri 4954 2088 4967 2101 se
rect 4967 2088 5498 2116
rect 14266 2107 14318 2113
rect 3981 2077 5493 2088
rect 3981 2025 4553 2077
rect 4605 2025 5493 2077
rect 3981 2013 5493 2025
rect 3981 1961 4553 2013
rect 4605 1961 5493 2013
rect 3981 1949 5493 1961
rect 3981 1897 4553 1949
rect 4605 1897 5493 1949
rect 3981 1886 5493 1897
rect 5769 2078 5885 2084
rect 10456 1972 10462 2088
rect 10578 1972 10584 2088
tri 12253 2084 12257 2088 sw
tri 13139 2084 13143 2088 se
rect 5769 1892 5885 1898
rect 12229 1886 13227 2084
rect 13428 2072 13544 2078
rect 14177 2045 14229 2051
rect 14177 1981 14229 1993
rect 14266 2043 14318 2055
tri 14318 2019 14343 2044 sw
rect 14318 1991 14389 2019
rect 14266 1985 14389 1991
tri 14229 1957 14254 1982 sw
rect 14229 1929 14305 1957
rect 14177 1923 14305 1929
rect 13428 1886 13544 1892
tri 11311 1837 11360 1886 ne
rect 11360 1826 12210 1886
tri 12210 1837 12259 1886 nw
rect 3981 1752 5405 1758
rect 3981 1700 3987 1752
rect 4039 1700 4051 1752
rect 4103 1700 4115 1752
rect 4167 1700 4179 1752
rect 4231 1700 4243 1752
rect 4295 1718 4327 1752
rect 4361 1718 4943 1752
rect 4977 1718 5015 1752
rect 5049 1718 5405 1752
rect 4295 1700 5405 1718
rect 3981 1692 5405 1700
rect 5769 1750 5885 1756
rect 5821 1698 5833 1750
rect 5769 1692 5885 1698
rect 10024 1750 10268 1756
rect 10076 1698 10088 1750
rect 10140 1698 10152 1750
rect 10204 1698 10216 1750
rect 10024 1692 10268 1698
rect 11059 1692 12253 1706
tri 11022 1664 11050 1692 ne
rect 11050 1664 12253 1692
rect 4539 1658 6662 1664
rect 4539 1624 4551 1658
rect 4585 1624 6610 1658
rect 4539 1612 6610 1624
rect 4539 1586 4597 1612
tri 4597 1587 4622 1612 nw
tri 6585 1587 6610 1612 ne
tri 11050 1655 11059 1664 ne
rect 6610 1594 6662 1606
rect 4539 1552 4551 1586
rect 4585 1552 4597 1586
rect 4539 1546 4597 1552
rect 4647 1570 4705 1576
rect 4647 1536 4659 1570
rect 4693 1536 4705 1570
rect 4647 1526 4705 1536
rect 4952 1532 4958 1584
rect 5010 1532 5022 1584
rect 5074 1572 5199 1584
rect 5074 1538 5081 1572
rect 5115 1538 5153 1572
rect 5187 1538 5199 1572
rect 5074 1532 5199 1538
tri 8455 1584 8480 1609 se
rect 8480 1596 8486 1648
rect 8538 1596 8544 1648
rect 8480 1584 8544 1596
rect 6610 1536 6662 1542
rect 7442 1532 8486 1584
rect 8538 1532 8544 1584
rect 11059 1560 12253 1664
tri 12253 1655 12290 1692 nw
tri 10325 1529 10328 1532 se
rect 10328 1529 14186 1532
tri 4705 1526 4708 1529 sw
tri 10322 1526 10325 1529 se
rect 10325 1526 14186 1529
rect 4647 1504 4708 1526
tri 4708 1504 4730 1526 sw
tri 10300 1504 10322 1526 se
rect 10322 1504 13634 1526
rect 4647 1498 13634 1504
rect 4647 1464 4659 1498
rect 4693 1492 13634 1498
rect 13668 1492 13706 1526
rect 13740 1492 14186 1526
rect 4693 1486 14186 1492
rect 4693 1464 10392 1486
rect 4647 1458 10392 1464
tri 10392 1458 10420 1486 nw
rect 5719 1424 8736 1430
rect 5719 1418 8618 1424
rect 5719 1384 5725 1418
rect 5759 1390 8618 1418
rect 8652 1390 8690 1424
rect 8724 1390 8736 1424
rect 10484 1401 10490 1453
rect 10542 1401 10554 1453
rect 10606 1401 12025 1453
rect 5759 1384 8736 1390
rect 5719 1372 5778 1384
tri 5778 1372 5790 1384 nw
rect 5719 1346 5765 1372
tri 5765 1359 5778 1372 nw
rect 5719 1312 5725 1346
rect 5759 1312 5765 1346
rect 9074 1320 9080 1372
rect 9132 1320 9144 1372
rect 9196 1320 10886 1372
rect 10938 1320 10950 1372
rect 11002 1320 11008 1372
rect 5719 1300 5765 1312
tri 6299 1286 6305 1292 se
rect 6305 1286 6312 1292
tri 6285 1272 6299 1286 se
rect 6299 1272 6312 1286
rect 4033 1247 6312 1272
rect 4033 1246 6057 1247
rect 4033 1241 5769 1246
rect 4033 1189 4553 1241
rect 4605 1189 5769 1241
rect 4033 1177 5769 1189
rect 4033 1125 4553 1177
rect 4605 1130 5769 1177
rect 5885 1141 6057 1246
rect 6163 1141 6312 1247
rect 5885 1130 6312 1141
rect 4605 1125 6312 1130
rect 4033 1090 6312 1125
rect 13428 1280 13544 1286
rect 13428 1094 13544 1100
rect 5833 860 6545 1062
rect 6690 1056 9080 1062
rect 6742 1010 9080 1056
rect 9132 1010 9138 1062
rect 6742 1004 9138 1010
rect 6690 998 9138 1004
rect 6690 992 9080 998
rect 6742 990 9080 992
rect 6742 984 6772 990
tri 6772 984 6778 990 nw
tri 9038 984 9044 990 ne
rect 9044 984 9080 990
tri 6742 954 6772 984 nw
tri 9044 954 9074 984 ne
rect 9074 946 9080 984
rect 9132 946 9138 998
rect 9166 1010 9172 1062
rect 9224 1056 9443 1062
rect 9224 1022 9397 1056
rect 9431 1022 9443 1056
rect 9224 1010 9443 1022
rect 9861 1053 10490 1062
rect 9861 1019 9873 1053
rect 9907 1019 9945 1053
rect 9979 1019 10490 1053
rect 9861 1010 10490 1019
rect 10542 1010 10554 1062
rect 10606 1010 10612 1062
rect 10995 1056 12177 1062
rect 10995 1022 11007 1056
rect 11041 1022 11079 1056
rect 11113 1022 12177 1056
rect 10995 1014 12177 1022
tri 12121 1010 12125 1014 ne
rect 12125 1010 12177 1014
rect 9166 998 9443 1010
rect 9166 946 9172 998
rect 9224 984 9443 998
tri 12125 988 12147 1010 ne
rect 12147 988 12177 1010
rect 9224 950 9397 984
rect 9431 950 9443 984
rect 9224 946 9443 950
rect 9166 944 9443 946
rect 6690 934 6742 940
rect 7807 882 7826 894
rect 7807 848 7819 882
rect 7807 842 7826 848
rect 7878 842 7890 894
rect 7942 842 7948 894
rect 13229 889 14462 895
rect 13281 855 14462 889
rect 3981 826 6054 832
rect 3981 720 5936 826
rect 6042 720 6054 826
rect 13229 825 13281 837
tri 13281 830 13306 855 nw
tri 6088 767 6135 814 se
rect 6135 767 6317 814
rect 13229 767 13281 773
rect 3981 714 6054 720
tri 6082 761 6088 767 se
rect 6088 761 6317 767
rect 6082 612 6317 761
rect 6082 584 6289 612
tri 6289 584 6317 612 nw
rect 6082 580 6285 584
tri 6285 580 6289 584 nw
rect 6082 578 6283 580
tri 6283 578 6285 580 nw
rect 4293 440 5354 492
rect 5406 440 5418 492
rect 5470 440 5482 492
rect 5534 440 5791 492
rect 6082 442 6280 578
tri 6280 575 6283 578 nw
rect 6605 574 7937 580
rect 6605 540 6617 574
rect 6651 540 6689 574
rect 6723 540 7819 574
rect 7853 540 7891 574
rect 7925 540 7937 574
rect 6605 534 7937 540
rect 8215 578 11739 584
rect 8215 544 8227 578
rect 8261 544 8299 578
rect 8333 575 11739 578
tri 11739 575 11748 584 sw
rect 8333 569 11748 575
rect 8333 544 11702 569
rect 8215 538 11702 544
tri 11665 535 11668 538 ne
rect 11668 535 11702 538
rect 11736 535 11748 569
tri 11668 534 11669 535 ne
rect 11669 534 11748 535
tri 11669 513 11690 534 ne
rect 8139 500 8447 506
tri 8121 459 8122 460 ne
rect 8122 459 8139 460
tri 6280 442 6297 459 sw
tri 8122 442 8139 459 ne
rect 8191 448 8203 500
rect 8255 448 8267 500
rect 8319 448 8331 500
rect 8383 448 8395 500
rect 9551 500 9859 506
rect 8139 442 8447 448
tri 8447 442 8465 460 nw
tri 9533 442 9551 460 ne
rect 9603 448 9615 500
rect 9667 448 9679 500
rect 9731 448 9743 500
rect 9795 448 9807 500
rect 11690 497 11748 534
rect 11690 463 11702 497
rect 11736 463 11748 497
rect 9859 457 9874 460
tri 9874 457 9877 460 nw
rect 11690 457 11748 463
rect 9551 442 9859 448
tri 9859 442 9874 457 nw
rect 6082 440 6297 442
tri 6297 440 6299 442 sw
rect 6082 437 6299 440
tri 6299 437 6302 440 sw
rect 9166 437 9230 438
rect 6082 413 6302 437
tri 6302 413 6326 437 sw
rect 6082 410 6326 413
tri 6326 410 6329 413 sw
tri 8712 410 8715 413 se
tri 4781 368 4792 379 se
rect 4792 373 4844 379
rect 3610 362 3662 368
tri 3662 349 3681 368 sw
tri 4762 349 4781 368 se
rect 4781 349 4792 368
rect 3662 330 3681 349
tri 3681 330 3700 349 sw
tri 4743 330 4762 349 se
rect 4762 330 4792 349
rect 3662 321 4792 330
rect 3662 310 4844 321
rect 3610 309 4844 310
rect 3610 298 4792 309
rect 3662 278 4792 298
rect 3662 275 3697 278
tri 3697 275 3700 278 nw
tri 4765 275 4768 278 ne
rect 4768 275 4792 278
rect 3610 240 3662 246
tri 3662 240 3697 275 nw
tri 4768 251 4792 275 ne
rect 4792 251 4844 257
rect 6082 240 8180 410
rect 8715 407 9023 413
tri 9023 410 9026 413 sw
rect 8767 355 8779 407
rect 8831 355 8843 407
rect 8895 355 8907 407
rect 8959 355 8971 407
rect 8715 349 9023 355
rect 9166 385 9172 437
rect 9224 385 9230 437
rect 9166 373 9230 385
tri 8180 324 8205 349 nw
rect 9166 321 9172 373
rect 9224 321 9230 373
rect 9258 407 9438 413
tri 9438 410 9441 413 sw
tri 11041 410 11044 413 se
rect 9310 355 9322 407
rect 9374 355 9386 407
rect 10107 358 10113 410
rect 10165 358 10177 410
rect 10229 358 10241 410
rect 10293 358 10299 410
rect 11044 407 11352 413
tri 11352 410 11355 413 sw
rect 9258 349 9438 355
rect 11096 355 11108 407
rect 11160 355 11172 407
rect 11224 355 11236 407
rect 11288 355 11300 407
rect 11044 349 11352 355
rect 9166 320 9230 321
rect 11489 315 12823 321
rect 11489 281 11501 315
rect 11535 281 11573 315
rect 11607 281 12823 315
rect 12965 291 13159 343
rect 13211 291 13223 343
rect 13275 291 13281 343
rect 11489 275 12823 281
tri 8180 240 8191 251 sw
rect 6082 226 8191 240
tri 8191 226 8205 240 sw
rect 6082 212 8180 226
tri 6082 198 6096 212 ne
rect 6096 198 8180 212
rect 3610 192 4924 198
rect 3662 140 4872 192
tri 6096 162 6132 198 ne
rect 6132 162 8180 198
rect 8715 220 9023 226
rect 8767 168 8779 220
rect 8831 168 8843 220
rect 8895 168 8907 220
rect 8959 168 8971 220
rect 8715 162 9023 168
rect 9258 220 9438 226
rect 9310 168 9322 220
rect 9374 168 9386 220
rect 11008 220 11352 226
rect 9258 162 9438 168
rect 10107 164 10113 216
rect 10165 164 10177 216
rect 10229 164 10241 216
rect 10293 164 10299 216
rect 11008 168 11044 220
rect 11096 168 11108 220
rect 11160 168 11172 220
rect 11224 168 11236 220
rect 11288 168 11300 220
rect 11008 162 11352 168
rect 3610 128 4924 140
rect 3662 76 4872 128
rect 3610 70 4924 76
rect 8140 126 8448 132
rect 8192 74 8204 126
rect 8256 74 8268 126
rect 8320 74 8332 126
rect 8384 74 8396 126
rect 8140 68 8448 74
rect 9551 126 9859 132
rect 9603 74 9615 126
rect 9667 74 9679 126
rect 9731 74 9743 126
rect 9795 74 9807 126
rect 9551 68 9859 74
rect 3610 27 3662 33
rect 3610 -37 3662 -25
rect 3610 -151 3662 -89
tri 3610 -173 3632 -151 ne
rect 3632 -173 3662 -151
tri 3662 -173 3706 -129 sw
tri 3632 -203 3662 -173 ne
rect 3662 -203 11682 -173
tri 3662 -225 3684 -203 ne
rect 3684 -225 11682 -203
rect 11734 -225 11746 -173
rect 11798 -225 11804 -173
rect 4556 -306 4562 -254
rect 4614 -306 4626 -254
rect 4678 -306 7274 -254
tri 7274 -306 7326 -254 sw
tri 7252 -352 7298 -306 ne
rect 7298 -352 7326 -306
tri 7326 -352 7372 -306 sw
tri 7298 -380 7326 -352 ne
rect 7326 -380 12242 -352
tri 7326 -404 7350 -380 ne
rect 7350 -404 12242 -380
rect 12294 -404 12306 -352
rect 12358 -404 12364 -352
<< via1 >>
rect 4633 5243 4685 5295
rect 6847 5281 6899 5333
rect 4633 5179 4685 5231
rect 6847 5217 6899 5269
rect 1680 5101 1732 5153
rect 1680 5037 1732 5089
rect 3585 5028 3637 5080
rect 3649 5028 3701 5080
rect 5355 5038 5407 5090
rect 5421 5038 5473 5090
rect 5487 5038 5539 5090
rect 5355 4969 5407 5021
rect 5421 4969 5473 5021
rect 5487 4969 5539 5021
rect 5355 4900 5407 4952
rect 5421 4900 5473 4952
rect 5487 4900 5539 4952
rect 5355 4831 5407 4883
rect 5421 4831 5473 4883
rect 5487 4831 5539 4883
rect 5355 4762 5407 4814
rect 5421 4762 5473 4814
rect 5487 4762 5539 4814
rect 5355 4693 5407 4745
rect 5421 4693 5473 4745
rect 5487 4693 5539 4745
rect 5355 4624 5407 4676
rect 5421 4624 5473 4676
rect 5487 4624 5539 4676
rect 6231 4669 6539 4977
rect 6847 4340 6899 4392
rect 6847 4274 6899 4326
rect 11937 4236 11989 4288
rect 4798 4128 4850 4180
rect 4862 4128 4914 4180
rect 8136 4137 8140 4140
rect 8140 4137 8188 4140
rect 8136 4088 8188 4137
rect 8136 4024 8188 4076
rect 11937 4172 11989 4224
rect 8216 4033 8268 4085
rect 8216 3969 8268 4021
rect 7006 3657 7058 3709
rect 7076 3657 7128 3709
rect 7146 3657 7198 3709
rect 7216 3657 7268 3709
rect 7286 3657 7338 3709
rect 7356 3657 7408 3709
rect 7426 3657 7478 3709
rect 7496 3657 7548 3709
rect 7566 3657 7618 3709
rect 7636 3657 7688 3709
rect 7705 3657 7757 3709
rect 6868 3576 6920 3628
rect 6868 3512 6920 3564
rect 7006 3575 7058 3627
rect 7076 3575 7128 3627
rect 7146 3575 7198 3627
rect 7216 3575 7268 3627
rect 7286 3575 7338 3627
rect 7356 3575 7408 3627
rect 7426 3575 7478 3627
rect 7496 3575 7548 3627
rect 7566 3575 7618 3627
rect 7636 3575 7688 3627
rect 7705 3575 7757 3627
rect 7006 3493 7058 3545
rect 7076 3493 7128 3545
rect 7146 3493 7198 3545
rect 7216 3493 7268 3545
rect 7286 3493 7338 3545
rect 7356 3493 7408 3545
rect 7426 3493 7478 3545
rect 7496 3493 7548 3545
rect 7566 3493 7618 3545
rect 7636 3493 7688 3545
rect 7705 3493 7757 3545
rect 9729 3453 9781 3505
rect 9729 3389 9781 3441
rect 6590 3304 6642 3356
rect 6590 3240 6642 3292
rect 6682 3304 6734 3356
rect 6682 3240 6734 3292
rect 12822 3309 12874 3361
rect 12886 3309 12938 3361
rect 13606 3303 13658 3355
rect 13606 3239 13658 3291
rect 3655 3150 3707 3202
rect 1028 3013 1144 3129
rect 1956 3013 2072 3129
rect 3655 3086 3707 3138
rect 8136 3154 8188 3206
rect 8818 3160 8870 3212
rect 8882 3160 8934 3212
rect 8946 3160 8998 3212
rect 9010 3160 9062 3212
rect 9074 3200 9126 3212
rect 9138 3200 9190 3212
rect 9074 3166 9103 3200
rect 9103 3166 9126 3200
rect 9138 3166 9175 3200
rect 9175 3166 9190 3200
rect 9074 3160 9126 3166
rect 9138 3160 9190 3166
rect 7826 3120 7878 3132
rect 7890 3120 7942 3132
rect 7826 3086 7858 3120
rect 7858 3086 7878 3120
rect 7890 3086 7892 3120
rect 7892 3086 7942 3120
rect 7826 3080 7878 3086
rect 7890 3080 7942 3086
rect 8136 3090 8188 3142
rect 10303 3147 10355 3199
rect 10367 3147 10419 3199
rect 10431 3147 10483 3199
rect 10495 3147 10547 3199
rect 10559 3147 10611 3199
rect 10880 3147 10932 3199
rect 8561 3080 8613 3132
rect 8625 3080 8677 3132
rect 8717 3080 8769 3132
rect 8781 3080 8833 3132
rect 10880 3120 10932 3135
rect 10880 3086 10906 3120
rect 10906 3086 10932 3120
rect 10880 3083 10932 3086
rect 10960 3147 11012 3199
rect 10960 3120 11012 3135
rect 10960 3086 10976 3120
rect 10976 3086 11010 3120
rect 11010 3086 11012 3120
rect 10960 3083 11012 3086
rect 9839 3023 9891 3075
rect 9903 3023 9955 3075
rect 6740 2943 6792 2995
rect 6804 2943 6856 2995
rect 14266 2937 14318 2989
rect 4872 2858 4924 2910
rect 7826 2882 7878 2934
rect 7890 2882 7942 2934
rect 8226 2882 8278 2934
rect 8290 2882 8342 2934
rect 8422 2881 8474 2933
rect 8486 2881 8538 2933
rect 14177 2875 14229 2927
rect 4872 2794 4924 2846
rect 14266 2873 14318 2925
rect 14177 2811 14229 2863
rect 5022 2706 5074 2758
rect 5022 2642 5074 2694
rect 2973 2415 3089 2595
rect 5424 2556 5476 2608
rect 5488 2556 5540 2608
rect 5424 2486 5476 2538
rect 5488 2486 5540 2538
rect 5424 2415 5476 2467
rect 5488 2415 5540 2467
rect 5424 2344 5476 2396
rect 5488 2344 5540 2396
rect 6897 2186 6949 2238
rect 6897 2122 6949 2174
rect 9805 2180 9857 2232
rect 9805 2116 9857 2168
rect 10462 2116 10514 2168
rect 10526 2116 10578 2168
rect 4553 2025 4605 2077
rect 4553 1961 4605 2013
rect 4553 1897 4605 1949
rect 5769 1898 5885 2078
rect 10462 1972 10578 2088
rect 13428 1892 13544 2072
rect 14266 2055 14318 2107
rect 14177 1993 14229 2045
rect 14266 1991 14318 2043
rect 14177 1929 14229 1981
rect 3987 1700 4039 1752
rect 4051 1700 4103 1752
rect 4115 1700 4167 1752
rect 4179 1700 4231 1752
rect 4243 1718 4255 1752
rect 4255 1718 4289 1752
rect 4289 1718 4295 1752
rect 4243 1700 4295 1718
rect 5769 1698 5821 1750
rect 5833 1698 5885 1750
rect 10024 1698 10076 1750
rect 10088 1698 10140 1750
rect 10152 1698 10204 1750
rect 10216 1698 10268 1750
rect 6610 1606 6662 1658
rect 4958 1532 5010 1584
rect 5022 1532 5074 1584
rect 6610 1542 6662 1594
rect 8486 1596 8538 1648
rect 8486 1532 8538 1584
rect 10490 1401 10542 1453
rect 10554 1401 10606 1453
rect 9080 1320 9132 1372
rect 9144 1320 9196 1372
rect 10886 1320 10938 1372
rect 10950 1320 11002 1372
rect 4553 1189 4605 1241
rect 4553 1125 4605 1177
rect 5769 1130 5885 1246
rect 13428 1100 13544 1280
rect 6690 1004 6742 1056
rect 9080 1010 9132 1062
rect 6690 940 6742 992
rect 9080 946 9132 998
rect 9172 1010 9224 1062
rect 10490 1010 10542 1062
rect 10554 1010 10606 1062
rect 9172 946 9224 998
rect 7826 882 7878 894
rect 7826 848 7853 882
rect 7853 848 7878 882
rect 7826 842 7878 848
rect 7890 882 7942 894
rect 7890 848 7891 882
rect 7891 848 7925 882
rect 7925 848 7942 882
rect 7890 842 7942 848
rect 13229 837 13281 889
rect 13229 773 13281 825
rect 5354 440 5406 492
rect 5418 440 5470 492
rect 5482 440 5534 492
rect 8139 448 8191 500
rect 8203 448 8255 500
rect 8267 448 8319 500
rect 8331 448 8383 500
rect 8395 448 8447 500
rect 9551 448 9603 500
rect 9615 448 9667 500
rect 9679 448 9731 500
rect 9743 448 9795 500
rect 9807 448 9859 500
rect 3610 310 3662 362
rect 4792 321 4844 373
rect 3610 246 3662 298
rect 4792 257 4844 309
rect 8715 355 8767 407
rect 8779 355 8831 407
rect 8843 355 8895 407
rect 8907 355 8959 407
rect 8971 355 9023 407
rect 9172 385 9224 437
rect 9172 321 9224 373
rect 9258 355 9310 407
rect 9322 355 9374 407
rect 9386 355 9438 407
rect 10113 358 10165 410
rect 10177 358 10229 410
rect 10241 358 10293 410
rect 11044 355 11096 407
rect 11108 355 11160 407
rect 11172 355 11224 407
rect 11236 355 11288 407
rect 11300 355 11352 407
rect 13159 291 13211 343
rect 13223 291 13275 343
rect 3610 140 3662 192
rect 4872 140 4924 192
rect 8715 168 8767 220
rect 8779 168 8831 220
rect 8843 168 8895 220
rect 8907 168 8959 220
rect 8971 168 9023 220
rect 9258 168 9310 220
rect 9322 168 9374 220
rect 9386 168 9438 220
rect 10113 164 10165 216
rect 10177 164 10229 216
rect 10241 164 10293 216
rect 11044 168 11096 220
rect 11108 168 11160 220
rect 11172 168 11224 220
rect 11236 168 11288 220
rect 11300 168 11352 220
rect 3610 76 3662 128
rect 4872 76 4924 128
rect 8140 74 8192 126
rect 8204 74 8256 126
rect 8268 74 8320 126
rect 8332 74 8384 126
rect 8396 74 8448 126
rect 9551 74 9603 126
rect 9615 74 9667 126
rect 9679 74 9731 126
rect 9743 74 9795 126
rect 9807 74 9859 126
rect 3610 -25 3662 27
rect 3610 -89 3662 -37
rect 11682 -225 11734 -173
rect 11746 -225 11798 -173
rect 4562 -306 4614 -254
rect 4626 -306 4678 -254
rect 12242 -404 12294 -352
rect 12306 -404 12358 -352
<< metal2 >>
rect 4633 5295 4685 5301
rect 4633 5231 4685 5243
rect 4633 5173 4685 5179
rect 1680 5153 1732 5159
rect 1680 5089 1732 5101
rect 1680 5031 1732 5037
rect 3579 5028 3585 5080
rect 3637 5028 3649 5080
rect 3701 5028 3707 5080
tri 3630 5021 3637 5028 ne
rect 3637 5021 3707 5028
tri 3637 5003 3655 5021 ne
rect 20 4944 136 4999
rect 651 3761 2449 3965
tri 651 3441 662 3452 ne
rect 662 3441 845 3452
tri 662 3389 714 3441 ne
rect 714 3389 845 3441
tri 714 3361 742 3389 ne
rect 742 3361 845 3389
tri 742 3356 747 3361 ne
rect 747 3356 845 3361
tri 747 3304 799 3356 ne
rect 799 3304 845 3356
tri 799 3303 800 3304 ne
rect 800 3303 845 3304
tri 800 3292 811 3303 ne
rect 811 3292 845 3303
tri 811 3258 845 3292 ne
rect 2255 3441 2438 3452
tri 2438 3441 2449 3452 nw
rect 2255 3389 2386 3441
tri 2386 3389 2438 3441 nw
rect 2255 3361 2358 3389
tri 2358 3361 2386 3389 nw
rect 2255 3356 2353 3361
tri 2353 3356 2358 3361 nw
rect 2255 3304 2301 3356
tri 2301 3304 2353 3356 nw
rect 2255 3303 2300 3304
tri 2300 3303 2301 3304 nw
rect 2255 3292 2289 3303
tri 2289 3292 2300 3303 nw
tri 2255 3258 2289 3292 nw
rect 3655 3202 3707 5021
rect 3655 3138 3707 3150
rect 1022 3013 1028 3129
rect 1144 3013 1150 3129
rect 1950 3013 1956 3129
rect 2072 3013 2078 3129
rect 3655 3080 3707 3086
rect 2967 2415 2973 2595
rect 3089 2415 3095 2595
rect 3981 1752 4301 5159
rect 3981 1700 3987 1752
rect 4039 1700 4051 1752
rect 4103 1700 4115 1752
rect 4167 1700 4179 1752
rect 4231 1700 4243 1752
rect 4295 1700 4301 1752
rect 3981 715 4301 1700
rect 4553 2077 4605 5159
rect 4553 2013 4605 2025
rect 4553 1949 4605 1961
rect 4553 1241 4605 1897
rect 4553 1177 4605 1189
rect 4553 1090 4605 1125
rect 3610 362 3662 368
rect 3610 298 3662 310
rect 3610 240 3662 246
rect 3610 192 3662 198
rect 3610 128 3662 140
rect 3610 70 3662 76
rect 3610 27 3662 33
rect 3610 -37 3662 -25
rect 3610 -95 3662 -89
tri 4585 -225 4633 -177 se
rect 4633 -225 4684 5173
rect 5348 5090 5540 5096
rect 5348 5038 5355 5090
rect 5407 5038 5421 5090
rect 5473 5038 5487 5090
rect 5539 5038 5540 5090
rect 5348 5021 5540 5038
rect 5348 4969 5355 5021
rect 5407 4969 5421 5021
rect 5473 4969 5487 5021
rect 5539 4969 5540 5021
rect 5348 4952 5540 4969
rect 5348 4900 5355 4952
rect 5407 4900 5421 4952
rect 5473 4900 5487 4952
rect 5539 4900 5540 4952
rect 5348 4883 5540 4900
rect 5348 4831 5355 4883
rect 5407 4831 5421 4883
rect 5473 4831 5487 4883
rect 5539 4831 5540 4883
rect 5348 4814 5540 4831
rect 5348 4762 5355 4814
rect 5407 4762 5421 4814
rect 5473 4762 5487 4814
rect 5539 4762 5540 4814
rect 5348 4745 5540 4762
rect 5348 4693 5355 4745
rect 5407 4693 5421 4745
rect 5473 4693 5487 4745
rect 5539 4693 5540 4745
rect 5348 4676 5540 4693
rect 5348 4624 5355 4676
rect 5407 4624 5421 4676
rect 5473 4624 5487 4676
rect 5539 4624 5540 4676
rect 4792 4128 4798 4180
rect 4850 4128 4862 4180
rect 4914 4128 4920 4180
rect 4792 4088 4880 4128
tri 4880 4088 4920 4128 nw
rect 4792 4085 4877 4088
tri 4877 4085 4880 4088 nw
rect 4792 4076 4868 4085
tri 4868 4076 4877 4085 nw
rect 4792 373 4844 4076
tri 4844 4052 4868 4076 nw
rect 4792 309 4844 321
rect 4792 251 4844 257
rect 4872 2910 4924 2916
rect 4872 2846 4924 2858
rect 4872 192 4924 2794
rect 5016 2706 5022 2758
rect 5074 2706 5080 2758
rect 5016 2694 5080 2706
rect 5016 2642 5022 2694
rect 5074 2642 5080 2694
tri 5013 1606 5016 1609 se
rect 5016 1606 5080 2642
tri 5003 1596 5013 1606 se
rect 5013 1596 5080 1606
tri 5001 1594 5003 1596 se
rect 5003 1594 5080 1596
tri 4991 1584 5001 1594 se
rect 5001 1584 5080 1594
rect 4952 1532 4958 1584
rect 5010 1532 5022 1584
rect 5074 1532 5080 1584
rect 5348 2608 5540 4624
rect 6225 4977 6545 5620
rect 6847 5333 6899 5339
rect 6847 5269 6899 5281
rect 6225 4669 6231 4977
rect 6539 4669 6545 4977
rect 5348 2556 5424 2608
rect 5476 2556 5488 2608
rect 5348 2538 5540 2556
rect 5348 2486 5424 2538
rect 5476 2486 5488 2538
rect 5348 2467 5540 2486
rect 5348 2415 5424 2467
rect 5476 2415 5488 2467
rect 5348 2396 5540 2415
rect 5348 2344 5424 2396
rect 5476 2344 5488 2396
rect 5348 492 5540 2344
rect 5769 2078 5885 4195
rect 5769 1750 5885 1898
rect 5821 1698 5833 1750
rect 5769 1246 5885 1698
rect 5769 1091 5885 1130
rect 6225 860 6545 4669
tri 6589 3361 6596 3368 se
rect 6596 3361 6648 5159
tri 6584 3356 6589 3361 se
rect 6589 3356 6648 3361
rect 6584 3304 6590 3356
rect 6642 3304 6648 3356
rect 6584 3292 6648 3304
rect 6584 3240 6590 3292
rect 6642 3240 6648 3292
rect 6676 3361 6728 5159
rect 6847 4392 6899 5217
tri 11684 5159 11826 5301 se
rect 6847 4326 6899 4340
rect 6847 4268 6899 4274
rect 6982 3709 7795 5159
rect 6982 3657 7006 3709
rect 7058 3657 7076 3709
rect 7128 3657 7146 3709
rect 7198 3657 7216 3709
rect 7268 3657 7286 3709
rect 7338 3657 7356 3709
rect 7408 3657 7426 3709
rect 7478 3657 7496 3709
rect 7548 3657 7566 3709
rect 7618 3657 7636 3709
rect 7688 3657 7705 3709
rect 7757 3657 7795 3709
rect 6862 3576 6868 3628
rect 6920 3576 6926 3628
rect 6862 3564 6926 3576
rect 6862 3512 6868 3564
rect 6920 3512 6926 3564
tri 6728 3361 6735 3368 sw
rect 6676 3356 6735 3361
tri 6735 3356 6740 3361 sw
rect 6676 3304 6682 3356
rect 6734 3304 6740 3356
rect 6676 3292 6740 3304
rect 6676 3240 6682 3292
rect 6734 3240 6740 3292
rect 6862 3082 6926 3512
rect 6982 3627 7795 3657
rect 6982 3575 7006 3627
rect 7058 3575 7076 3627
rect 7128 3575 7146 3627
rect 7198 3575 7216 3627
rect 7268 3575 7286 3627
rect 7338 3575 7356 3627
rect 7408 3575 7426 3627
rect 7478 3575 7496 3627
rect 7548 3575 7566 3627
rect 7618 3575 7636 3627
rect 7688 3575 7705 3627
rect 7757 3575 7795 3627
rect 6982 3545 7795 3575
rect 6982 3493 7006 3545
rect 7058 3493 7076 3545
rect 7128 3493 7146 3545
rect 7198 3493 7216 3545
rect 7268 3493 7286 3545
rect 7338 3493 7356 3545
rect 7408 3493 7426 3545
rect 7478 3493 7496 3545
rect 7548 3493 7566 3545
rect 7618 3493 7636 3545
rect 7688 3493 7705 3545
rect 7757 3493 7795 3545
rect 6982 3187 7795 3493
rect 6982 3157 7765 3187
tri 7765 3157 7795 3187 nw
rect 6982 3116 7764 3157
tri 7764 3156 7765 3157 nw
tri 7895 3156 7896 3157 se
rect 7896 3156 7948 5159
tri 7893 3154 7895 3156 se
rect 7895 3154 7948 3156
tri 7886 3147 7893 3154 se
rect 7893 3147 7948 3154
tri 7881 3142 7886 3147 se
rect 7886 3142 7948 3147
tri 7871 3132 7881 3142 se
rect 7881 3132 7948 3142
tri 6982 3093 7005 3116 ne
tri 6862 3080 6864 3082 ne
rect 6864 3080 6926 3082
tri 6926 3080 6938 3092 sw
tri 6864 3075 6869 3080 ne
rect 6869 3075 6938 3080
tri 6938 3075 6943 3080 sw
tri 6869 3069 6875 3075 ne
rect 6875 3069 6943 3075
tri 6943 3069 6949 3075 sw
tri 6875 3047 6897 3069 ne
rect 6734 2943 6740 2995
rect 6792 2943 6804 2995
rect 6856 2943 6862 2995
tri 6773 2937 6779 2943 ne
rect 6779 2937 6862 2943
tri 6779 2934 6782 2937 ne
rect 6782 2934 6862 2937
tri 6782 2918 6798 2934 ne
rect 6798 2308 6862 2934
rect 6897 2238 6949 3069
rect 6897 2174 6949 2186
rect 6897 2116 6949 2122
rect 7005 2827 7764 3116
rect 7820 3080 7826 3132
rect 7878 3080 7890 3132
rect 7942 3080 7948 3132
rect 8136 4140 8188 4146
rect 8136 4076 8188 4088
rect 8136 3206 8188 4024
rect 8216 4085 8268 4091
rect 8216 4021 8268 4033
rect 8216 3963 8268 3969
rect 8136 3142 8188 3154
rect 8136 3084 8188 3090
tri 8280 2943 8296 2959 se
rect 8296 2943 8348 5159
tri 8621 3147 8631 3157 se
rect 8631 3147 8683 5159
tri 8609 3135 8621 3147 se
rect 8621 3135 8683 3147
tri 8606 3132 8609 3135 se
rect 8609 3132 8683 3135
rect 8555 3080 8561 3132
rect 8613 3080 8625 3132
rect 8677 3080 8683 3132
rect 8711 3147 8775 5159
rect 8803 4006 9047 5159
rect 9167 4002 9475 4262
tri 9167 3874 9295 4002 ne
rect 9295 3781 9475 4002
rect 8812 3212 9196 3620
rect 8812 3160 8818 3212
rect 8870 3160 8882 3212
rect 8934 3160 8946 3212
rect 8998 3160 9010 3212
rect 9062 3160 9074 3212
rect 9126 3160 9138 3212
rect 9190 3160 9196 3212
rect 9723 3453 9729 3505
rect 9781 3453 9787 3505
rect 9723 3441 9787 3453
rect 9723 3389 9729 3441
rect 9781 3389 9787 3441
tri 8775 3147 8785 3157 sw
rect 8711 3135 8785 3147
tri 8785 3135 8797 3147 sw
rect 8711 3132 8797 3135
tri 8797 3132 8800 3135 sw
rect 8711 3080 8717 3132
rect 8769 3080 8781 3132
rect 8833 3080 8839 3132
tri 8274 2937 8280 2943 se
rect 8280 2937 8348 2943
tri 8271 2934 8274 2937 se
rect 8274 2934 8348 2937
rect 7820 2882 7826 2934
rect 7878 2882 7890 2934
rect 7942 2882 7948 2934
rect 8220 2882 8226 2934
rect 8278 2882 8290 2934
rect 8342 2882 8348 2934
tri 7871 2881 7872 2882 ne
rect 7872 2881 7948 2882
rect 8416 2881 8422 2933
rect 8474 2881 8486 2933
rect 8538 2881 8544 2933
tri 7872 2875 7878 2881 ne
rect 7878 2875 7948 2881
tri 8455 2875 8461 2881 ne
rect 8461 2875 8544 2881
tri 7878 2873 7880 2875 ne
rect 7880 2873 7948 2875
tri 8461 2873 8463 2875 ne
rect 8463 2873 8544 2875
tri 7880 2863 7890 2873 ne
rect 7890 2863 7948 2873
tri 8463 2863 8473 2873 ne
rect 8473 2863 8544 2873
tri 7890 2858 7895 2863 ne
rect 7895 2858 7948 2863
tri 7764 2827 7795 2858 sw
tri 7895 2857 7896 2858 ne
tri 7001 2088 7005 2092 se
rect 7005 2088 7795 2827
tri 6982 2069 7001 2088 se
rect 7001 2069 7795 2088
rect 6982 1801 7795 2069
rect 6982 1750 7744 1801
tri 7744 1750 7795 1801 nw
rect 6982 1698 7692 1750
tri 7692 1698 7744 1750 nw
rect 6610 1658 6662 1664
rect 6610 1594 6662 1606
rect 5348 440 5354 492
rect 5406 440 5418 492
rect 5470 440 5482 492
rect 5534 440 5540 492
rect 4872 128 4924 140
rect 4872 70 4924 76
rect 6610 0 6662 1542
rect 6982 1329 7684 1698
tri 7684 1690 7692 1698 nw
tri 7684 1329 7692 1337 sw
rect 6982 1090 7692 1329
rect 6690 1056 6742 1062
rect 6690 992 6742 1004
rect 6690 0 6742 940
tri 7871 894 7896 919 se
rect 7896 894 7948 2858
tri 8473 2856 8480 2863 ne
rect 8480 1648 8544 2863
rect 9723 2782 9787 3389
rect 9833 3083 9885 5159
rect 10088 4989 10124 5159
rect 10296 5106 10604 5159
rect 9952 4288 10080 4386
tri 10080 4288 10178 4386 sw
rect 9952 4262 10178 4288
tri 10178 4262 10204 4288 sw
rect 9952 3800 10268 4196
tri 9953 3389 10016 3452 ne
rect 10016 3389 10268 3452
tri 10016 3381 10024 3389 ne
tri 9885 3083 9902 3100 sw
rect 9833 3075 9902 3083
tri 9902 3075 9910 3083 sw
rect 9833 3023 9839 3075
rect 9891 3023 9903 3075
rect 9955 3023 9961 3075
tri 9723 2732 9773 2782 ne
rect 9773 2732 9787 2782
tri 9787 2732 9863 2808 sw
tri 9773 2718 9787 2732 ne
rect 9787 2718 9863 2732
tri 9787 2706 9799 2718 ne
rect 9799 2232 9863 2718
rect 9799 2180 9805 2232
rect 9857 2180 9863 2232
rect 9799 2168 9863 2180
rect 9799 2116 9805 2168
rect 9857 2116 9863 2168
rect 8480 1596 8486 1648
rect 8538 1596 8544 1648
rect 8480 1584 8544 1596
rect 8480 1532 8486 1584
rect 8538 1532 8544 1584
rect 7820 842 7826 894
rect 7878 842 7890 894
rect 7942 842 7948 894
rect 8136 500 8452 1108
rect 8136 448 8139 500
rect 8191 448 8203 500
rect 8255 448 8267 500
rect 8319 448 8331 500
rect 8383 448 8395 500
rect 8447 448 8452 500
rect 8136 126 8452 448
rect 8711 407 9027 2110
rect 10024 1750 10268 3389
rect 10303 3199 10611 3205
rect 10355 3147 10367 3199
rect 10419 3147 10431 3199
rect 10483 3147 10495 3199
rect 10547 3147 10559 3199
rect 10303 3141 10611 3147
rect 10880 3199 10932 5159
rect 10880 3135 10932 3147
rect 10880 3077 10932 3083
rect 10960 3199 11012 5142
rect 11040 5106 11356 5158
tri 11850 5076 11864 5090 sw
rect 10960 3135 11012 3147
rect 10960 3077 11012 3083
rect 11492 2544 11864 5076
rect 11937 4288 11989 4294
rect 11937 4224 11989 4236
rect 10456 2116 10462 2168
rect 10514 2116 10526 2168
rect 10578 2116 10584 2168
rect 10456 2088 10584 2116
rect 10456 1972 10462 2088
rect 10578 1972 10584 2088
tri 11915 1756 11937 1778 se
rect 11937 1756 11989 4172
tri 12847 3361 12892 3406 se
rect 12892 3361 12944 5159
rect 13429 5109 13555 5156
rect 13428 5003 13556 5079
rect 12816 3309 12822 3361
rect 12874 3309 12886 3361
rect 12938 3309 12944 3361
rect 13606 3355 13658 5159
rect 13864 5106 14149 5158
rect 13606 3291 13658 3303
rect 13879 4443 14147 4452
rect 13935 4387 13985 4443
rect 14041 4387 14091 4443
rect 13879 4362 14147 4387
rect 13935 4306 13985 4362
rect 14041 4306 14091 4362
rect 13879 4281 14147 4306
rect 13935 4225 13985 4281
rect 14041 4225 14091 4281
rect 13879 4200 14147 4225
rect 13935 4144 13985 4200
rect 14041 4144 14091 4200
rect 13879 4119 14147 4144
rect 13935 4063 13985 4119
rect 14041 4063 14091 4119
rect 13879 4038 14147 4063
rect 13935 3982 13985 4038
rect 14041 3982 14091 4038
rect 13879 3957 14147 3982
rect 13935 3901 13985 3957
rect 14041 3901 14091 3957
rect 13879 3876 14147 3901
rect 13935 3820 13985 3876
rect 14041 3820 14091 3876
rect 13879 3795 14147 3820
rect 13935 3739 13985 3795
rect 14041 3739 14091 3795
rect 13879 3714 14147 3739
rect 13935 3658 13985 3714
rect 14041 3658 14091 3714
rect 13879 3633 14147 3658
rect 13935 3577 13985 3633
rect 14041 3577 14091 3633
rect 13879 3551 14147 3577
rect 13935 3495 13985 3551
rect 14041 3495 14091 3551
rect 13879 3469 14147 3495
rect 13935 3413 13985 3469
rect 14041 3413 14091 3469
rect 13879 3387 14147 3413
rect 13935 3331 13985 3387
rect 14041 3331 14091 3387
rect 13879 3305 14147 3331
rect 13935 3249 13985 3305
rect 14041 3249 14091 3305
rect 13879 3240 14147 3249
rect 13606 3233 13658 3239
rect 14266 2989 14318 2995
rect 14177 2927 14229 2933
rect 14177 2863 14229 2875
tri 12582 2168 12584 2170 ne
rect 12584 2168 12690 2170
tri 12584 2132 12620 2168 ne
tri 12542 1972 12620 2050 se
rect 12620 2022 12690 2168
tri 12690 2150 12710 2170 nw
tri 12522 1952 12542 1972 se
rect 12542 1952 12620 1972
tri 12620 1952 12690 2022 nw
rect 13428 2072 13544 2078
tri 12462 1892 12522 1952 se
rect 12522 1892 12560 1952
tri 12560 1892 12620 1952 nw
rect 14177 2045 14229 2811
rect 14177 1981 14229 1993
rect 14266 2925 14318 2937
rect 14266 2107 14318 2873
rect 14266 2043 14318 2055
rect 14266 1985 14318 1991
rect 14177 1923 14229 1929
tri 12461 1891 12462 1892 se
rect 12462 1891 12554 1892
tri 12456 1886 12461 1891 se
rect 12461 1886 12554 1891
tri 12554 1886 12560 1892 nw
rect 13428 1886 13544 1892
tri 12424 1854 12456 1886 se
rect 12456 1854 12522 1886
tri 12522 1854 12554 1886 nw
tri 12326 1756 12424 1854 se
tri 12424 1756 12522 1854 nw
rect 10076 1698 10088 1750
rect 10140 1698 10152 1750
rect 10204 1698 10216 1750
tri 11863 1704 11915 1756 se
rect 11915 1704 11937 1756
tri 11937 1704 11989 1756 nw
tri 12274 1704 12326 1756 se
rect 12326 1704 12347 1756
rect 9074 1320 9080 1372
rect 9132 1320 9144 1372
rect 9196 1320 9202 1372
rect 9074 1062 9138 1320
tri 9138 1295 9163 1320 nw
rect 10024 1287 10268 1698
tri 11851 1692 11863 1704 se
rect 11863 1692 11925 1704
tri 11925 1692 11937 1704 nw
tri 12262 1692 12274 1704 se
rect 12274 1692 12347 1704
tri 11807 1648 11851 1692 se
rect 11851 1648 11863 1692
tri 11789 1630 11807 1648 se
rect 11807 1630 11863 1648
tri 11863 1630 11925 1692 nw
tri 12249 1679 12262 1692 se
rect 12262 1679 12347 1692
tri 12347 1679 12424 1756 nw
rect 12249 1664 12332 1679
tri 12332 1664 12347 1679 nw
tri 11752 1593 11789 1630 se
rect 11789 1593 11826 1630
tri 11826 1593 11863 1630 nw
rect 10484 1401 10490 1453
rect 10542 1401 10554 1453
rect 10606 1401 10612 1453
rect 9074 1010 9080 1062
rect 9132 1010 9138 1062
rect 9074 998 9138 1010
rect 9074 946 9080 998
rect 9132 946 9138 998
rect 9166 1010 9172 1062
rect 9224 1010 9230 1062
rect 9166 998 9230 1010
rect 9166 946 9172 998
rect 9224 946 9230 998
rect 8711 355 8715 407
rect 8767 355 8779 407
rect 8831 355 8843 407
rect 8895 355 8907 407
rect 8959 355 8971 407
rect 9023 355 9027 407
rect 8711 220 9027 355
rect 9166 437 9230 946
rect 9166 385 9172 437
rect 9224 385 9230 437
rect 9166 373 9230 385
rect 9166 321 9172 373
rect 9224 321 9230 373
rect 9258 407 9438 808
rect 9310 355 9322 407
rect 9374 355 9386 407
rect 8711 168 8715 220
rect 8767 168 8779 220
rect 8831 168 8843 220
rect 8895 168 8907 220
rect 8959 168 8971 220
rect 9023 168 9027 220
rect 8711 162 9027 168
rect 9258 220 9438 355
rect 9310 168 9322 220
rect 9374 168 9386 220
rect 9258 162 9438 168
rect 9547 500 9863 1108
rect 10484 1062 10612 1401
rect 10484 1010 10490 1062
rect 10542 1010 10554 1062
rect 10606 1010 10612 1062
rect 10880 1320 10886 1372
rect 10938 1320 10950 1372
rect 11002 1320 11008 1372
rect 10880 948 11008 1320
rect 9547 448 9551 500
rect 9603 448 9615 500
rect 9667 448 9679 500
rect 9731 448 9743 500
rect 9795 448 9807 500
rect 9859 448 9863 500
rect 8136 74 8140 126
rect 8192 74 8204 126
rect 8256 74 8268 126
rect 8320 74 8332 126
rect 8384 74 8396 126
rect 8448 74 8452 126
rect 8136 68 8452 74
rect 9547 126 9863 448
rect 10107 410 10299 808
rect 10107 358 10113 410
rect 10165 358 10177 410
rect 10229 358 10241 410
rect 10293 358 10299 410
rect 10107 216 10299 358
rect 10107 164 10113 216
rect 10165 164 10177 216
rect 10229 164 10241 216
rect 10293 164 10299 216
rect 11040 407 11356 612
rect 11040 355 11044 407
rect 11096 355 11108 407
rect 11160 355 11172 407
rect 11224 355 11236 407
rect 11288 355 11300 407
rect 11352 355 11356 407
rect 11040 220 11356 355
rect 11040 168 11044 220
rect 11096 168 11108 220
rect 11160 168 11172 220
rect 11224 168 11236 220
rect 11288 168 11300 220
rect 11352 168 11356 220
rect 11040 162 11356 168
rect 9547 74 9551 126
rect 9603 74 9615 126
rect 9667 74 9679 126
rect 9731 74 9743 126
rect 9795 74 9807 126
rect 9859 74 9863 126
rect 9547 68 9863 74
tri 11676 -173 11752 -97 se
rect 11752 -173 11804 1593
tri 11804 1571 11826 1593 nw
rect 11676 -225 11682 -173
rect 11734 -225 11746 -173
rect 11798 -225 11804 -173
tri 4556 -254 4585 -225 se
rect 4585 -254 4684 -225
rect 4556 -306 4562 -254
rect 4614 -306 4626 -254
rect 4678 -306 4684 -254
rect 12249 -339 12316 1664
tri 12316 1648 12332 1664 nw
rect 13428 1280 13544 1286
rect 13428 1094 13544 1100
rect 13229 889 13281 895
rect 13229 825 13281 837
rect 12576 467 12729 545
tri 13204 343 13229 368 se
rect 13229 343 13281 773
rect 13153 291 13159 343
rect 13211 291 13223 343
rect 13275 291 13281 343
tri 13755 54 13814 113 sw
tri 12316 -339 12351 -304 sw
tri 12236 -352 12249 -339 se
rect 12249 -352 12351 -339
tri 12351 -352 12364 -339 sw
rect 12236 -404 12242 -352
rect 12294 -404 12306 -352
rect 12358 -404 12364 -352
<< via2 >>
rect 13879 4387 13935 4443
rect 13985 4387 14041 4443
rect 14091 4387 14147 4443
rect 13879 4306 13935 4362
rect 13985 4306 14041 4362
rect 14091 4306 14147 4362
rect 13879 4225 13935 4281
rect 13985 4225 14041 4281
rect 14091 4225 14147 4281
rect 13879 4144 13935 4200
rect 13985 4144 14041 4200
rect 14091 4144 14147 4200
rect 13879 4063 13935 4119
rect 13985 4063 14041 4119
rect 14091 4063 14147 4119
rect 13879 3982 13935 4038
rect 13985 3982 14041 4038
rect 14091 3982 14147 4038
rect 13879 3901 13935 3957
rect 13985 3901 14041 3957
rect 14091 3901 14147 3957
rect 13879 3820 13935 3876
rect 13985 3820 14041 3876
rect 14091 3820 14147 3876
rect 13879 3739 13935 3795
rect 13985 3739 14041 3795
rect 14091 3739 14147 3795
rect 13879 3658 13935 3714
rect 13985 3658 14041 3714
rect 14091 3658 14147 3714
rect 13879 3577 13935 3633
rect 13985 3577 14041 3633
rect 14091 3577 14147 3633
rect 13879 3495 13935 3551
rect 13985 3495 14041 3551
rect 14091 3495 14147 3551
rect 13879 3413 13935 3469
rect 13985 3413 14041 3469
rect 14091 3413 14147 3469
rect 13879 3331 13935 3387
rect 13985 3331 14041 3387
rect 14091 3331 14147 3387
rect 13879 3249 13935 3305
rect 13985 3249 14041 3305
rect 14091 3249 14147 3305
<< metal3 >>
rect 13874 4443 14152 4448
rect 13874 4387 13879 4443
rect 13935 4387 13985 4443
rect 14041 4387 14091 4443
rect 14147 4387 14152 4443
rect 13874 4362 14152 4387
rect 13874 4306 13879 4362
rect 13935 4306 13985 4362
rect 14041 4306 14091 4362
rect 14147 4306 14152 4362
rect 13874 4281 14152 4306
rect 13874 4225 13879 4281
rect 13935 4225 13985 4281
rect 14041 4225 14091 4281
rect 14147 4225 14152 4281
rect 13874 4200 14152 4225
rect 13874 4144 13879 4200
rect 13935 4144 13985 4200
rect 14041 4144 14091 4200
rect 14147 4144 14152 4200
rect 13874 4119 14152 4144
rect 13874 4063 13879 4119
rect 13935 4063 13985 4119
rect 14041 4063 14091 4119
rect 14147 4063 14152 4119
rect 13874 4038 14152 4063
rect 13874 3982 13879 4038
rect 13935 3982 13985 4038
rect 14041 3982 14091 4038
rect 14147 3982 14152 4038
rect 13874 3957 14152 3982
rect 13874 3901 13879 3957
rect 13935 3901 13985 3957
rect 14041 3901 14091 3957
rect 14147 3901 14152 3957
rect 13874 3876 14152 3901
rect 13874 3820 13879 3876
rect 13935 3820 13985 3876
rect 14041 3820 14091 3876
rect 14147 3820 14152 3876
rect 13874 3795 14152 3820
rect 13874 3739 13879 3795
rect 13935 3739 13985 3795
rect 14041 3739 14091 3795
rect 14147 3739 14152 3795
rect 13874 3714 14152 3739
rect 13874 3658 13879 3714
rect 13935 3658 13985 3714
rect 14041 3658 14091 3714
rect 14147 3658 14152 3714
rect 13874 3633 14152 3658
rect 13874 3577 13879 3633
rect 13935 3577 13985 3633
rect 14041 3577 14091 3633
rect 14147 3577 14152 3633
rect 13874 3551 14152 3577
rect 13874 3495 13879 3551
rect 13935 3495 13985 3551
rect 14041 3495 14091 3551
rect 14147 3495 14152 3551
rect 13874 3469 14152 3495
rect 13874 3413 13879 3469
rect 13935 3413 13985 3469
rect 14041 3413 14091 3469
rect 14147 3413 14152 3469
rect 13874 3387 14152 3413
rect 13874 3331 13879 3387
rect 13935 3331 13985 3387
rect 14041 3331 14091 3387
rect 14147 3331 14152 3387
rect 13874 3305 14152 3331
rect 13874 3249 13879 3305
rect 13935 3249 13985 3305
rect 14041 3249 14091 3305
rect 14147 3249 14152 3305
rect 13874 3244 14152 3249
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_0
timestamp 1707688321
transform 0 1 6064 1 0 3005
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_1
timestamp 1707688321
transform 1 0 9397 0 -1 1056
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_2
timestamp 1707688321
transform 1 0 11702 0 -1 569
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_3
timestamp 1707688321
transform 1 0 4551 0 -1 1658
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_4
timestamp 1707688321
transform 1 0 5644 0 1 2794
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_5
timestamp 1707688321
transform 1 0 4659 0 1 1464
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_0
timestamp 1707688321
transform -1 0 8333 0 1 544
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_1
timestamp 1707688321
transform -1 0 9979 0 1 1019
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_2
timestamp 1707688321
transform -1 0 11607 0 1 281
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_3
timestamp 1707688321
transform -1 0 5049 0 1 1718
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_4
timestamp 1707688321
transform -1 0 4361 0 1 1718
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_5
timestamp 1707688321
transform -1 0 11113 0 -1 1056
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_6
timestamp 1707688321
transform 0 -1 5759 1 0 1312
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_7
timestamp 1707688321
transform 1 0 5696 0 -1 3200
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_8
timestamp 1707688321
transform 1 0 7610 0 1 3086
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_9
timestamp 1707688321
transform 1 0 9351 0 1 3239
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_10
timestamp 1707688321
transform 1 0 7148 0 1 3246
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_11
timestamp 1707688321
transform 1 0 6334 0 1 3246
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_12
timestamp 1707688321
transform 1 0 13634 0 1 1492
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_13
timestamp 1707688321
transform 1 0 5081 0 1 1538
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_14
timestamp 1707688321
transform 1 0 8618 0 1 1390
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_15
timestamp 1707688321
transform 1 0 10976 0 1 3086
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_16
timestamp 1707688321
transform 1 0 10800 0 1 3086
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_17
timestamp 1707688321
transform 1 0 9524 0 1 3086
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_18
timestamp 1707688321
transform 1 0 8949 0 1 3321
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_19
timestamp 1707688321
transform 1 0 8424 0 1 3086
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_20
timestamp 1707688321
transform 1 0 7786 0 1 3086
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_21
timestamp 1707688321
transform 1 0 6617 0 1 540
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_22
timestamp 1707688321
transform 1 0 7819 0 1 540
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_23
timestamp 1707688321
transform 1 0 7819 0 1 848
box 0 0 1 1
use L1M1_CDNS_5246887918559  L1M1_CDNS_5246887918559_0
timestamp 1707688321
transform -1 0 6042 0 -1 826
box 0 0 1 1
use L1M1_CDNS_5246887918559  L1M1_CDNS_5246887918559_1
timestamp 1707688321
transform 1 0 6057 0 1 1141
box 0 0 1 1
use L1M1_CDNS_5246887918590  L1M1_CDNS_5246887918590_0
timestamp 1707688321
transform 1 0 9103 0 1 3166
box 0 0 1 1
use L1M1_CDNS_52468879185192  L1M1_CDNS_52468879185192_0
timestamp 1707688321
transform 0 1 8566 1 0 3172
box 0 0 1 1
use L1M1_CDNS_52468879185335  L1M1_CDNS_52468879185335_0
timestamp 1707688321
transform -1 0 12241 0 1 1604
box -12 -6 1126 40
use L1M1_CDNS_52468879185381  L1M1_CDNS_52468879185381_0
timestamp 1707688321
transform -1 0 10599 0 1 3165
box -12 -6 910 40
use L1M1_CDNS_524688791851011  L1M1_CDNS_524688791851011_0
timestamp 1707688321
transform 1 0 11028 0 1 1698
box -12 -6 1198 40
use L1M1_CDNS_524688791851012  L1M1_CDNS_524688791851012_0
timestamp 1707688321
transform 1 0 4305 0 1 449
box -12 -6 1486 40
use L1M1_CDNS_524688791851040  L1M1_CDNS_524688791851040_0
timestamp 1707688321
transform -1 0 5131 0 1 2477
box -12 -6 1054 40
use L1M1_CDNS_524688791851191  L1M1_CDNS_524688791851191_0
timestamp 1707688321
transform 1 0 11423 0 -1 3186
box -12 -6 766 112
use L1M1_CDNS_524688791851192  L1M1_CDNS_524688791851192_0
timestamp 1707688321
transform 1 0 7336 0 -1 3352
box -12 -6 982 112
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_0
timestamp 1707688321
transform 0 -1 8188 -1 0 3212
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_1
timestamp 1707688321
transform 0 -1 6662 -1 0 1664
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_2
timestamp 1707688321
transform 0 -1 6742 -1 0 1062
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_3
timestamp 1707688321
transform 0 1 10960 -1 0 3205
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_4
timestamp 1707688321
transform 0 1 10880 -1 0 3205
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_5
timestamp 1707688321
transform -1 0 5080 0 1 1532
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_6
timestamp 1707688321
transform -1 0 3707 0 1 5028
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_7
timestamp 1707688321
transform -1 0 7948 0 1 3080
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_8
timestamp 1707688321
transform -1 0 8683 0 1 3080
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_9
timestamp 1707688321
transform -1 0 12944 0 -1 3361
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_10
timestamp 1707688321
transform -1 0 8544 0 -1 2933
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_11
timestamp 1707688321
transform -1 0 7948 0 -1 894
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_12
timestamp 1707688321
transform -1 0 8348 0 -1 2934
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_13
timestamp 1707688321
transform -1 0 7948 0 -1 2934
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_14
timestamp 1707688321
transform 0 1 6897 1 0 2116
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_15
timestamp 1707688321
transform 0 1 13606 1 0 3233
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_16
timestamp 1707688321
transform 0 1 3655 1 0 3080
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_17
timestamp 1707688321
transform 0 -1 1732 1 0 5031
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_18
timestamp 1707688321
transform 0 -1 13281 1 0 767
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_19
timestamp 1707688321
transform 0 -1 4605 1 0 1119
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_20
timestamp 1707688321
transform 1 0 9833 0 -1 3075
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_21
timestamp 1707688321
transform 1 0 10484 0 1 1010
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_22
timestamp 1707688321
transform 1 0 10484 0 1 1401
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_23
timestamp 1707688321
transform 1 0 8711 0 1 3080
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_24
timestamp 1707688321
transform 1 0 10880 0 1 1320
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_25
timestamp 1707688321
transform 1 0 9074 0 1 1320
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_26
timestamp 1707688321
transform 1 0 6734 0 1 2943
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_27
timestamp 1707688321
transform 1 0 13153 0 1 291
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_28
timestamp 1707688321
transform 1 0 10456 0 1 2116
box 0 0 1 1
use M1M2_CDNS_52468879185198  M1M2_CDNS_52468879185198_0
timestamp 1707688321
transform 0 1 5769 -1 0 2084
box 0 0 1 1
use M1M2_CDNS_52468879185198  M1M2_CDNS_52468879185198_1
timestamp 1707688321
transform 0 -1 13544 1 0 1094
box 0 0 1 1
use M1M2_CDNS_52468879185198  M1M2_CDNS_52468879185198_2
timestamp 1707688321
transform 0 -1 13544 1 0 1886
box 0 0 1 1
use M1M2_CDNS_52468879185199  M1M2_CDNS_52468879185199_0
timestamp 1707688321
transform 0 1 5769 -1 0 1252
box 0 0 1 1
use M1M2_CDNS_52468879185199  M1M2_CDNS_52468879185199_1
timestamp 1707688321
transform 1 0 10456 0 1 1972
box 0 0 1 1
use M1M2_CDNS_52468879185199  M1M2_CDNS_52468879185199_2
timestamp 1707688321
transform 1 0 1950 0 1 3013
box 0 0 1 1
use M1M2_CDNS_52468879185199  M1M2_CDNS_52468879185199_3
timestamp 1707688321
transform 1 0 1022 0 1 3013
box 0 0 1 1
use M1M2_CDNS_52468879185200  M1M2_CDNS_52468879185200_0
timestamp 1707688321
transform 1 0 2967 0 1 2415
box 0 0 1 1
use M1M2_CDNS_52468879185201  M1M2_CDNS_52468879185201_0
timestamp 1707688321
transform -1 0 4301 0 -1 831
box 0 0 320 116
use M1M2_CDNS_52468879185202  M1M2_CDNS_52468879185202_0
timestamp 1707688321
transform -1 0 4301 0 -1 1752
box 0 0 1 1
use M1M2_CDNS_52468879185203  M1M2_CDNS_52468879185203_0
timestamp 1707688321
transform 0 -1 4605 -1 0 2083
box 0 0 1 1
use M1M2_CDNS_52468879185203  M1M2_CDNS_52468879185203_1
timestamp 1707688321
transform 1 0 10107 0 1 358
box 0 0 1 1
use M1M2_CDNS_52468879185203  M1M2_CDNS_52468879185203_2
timestamp 1707688321
transform 1 0 10107 0 1 164
box 0 0 1 1
use M1M2_CDNS_52468879185203  M1M2_CDNS_52468879185203_3
timestamp 1707688321
transform 1 0 5348 0 1 440
box 0 0 1 1
use M1M2_CDNS_52468879185204  M1M2_CDNS_52468879185204_0
timestamp 1707688321
transform 1 0 8812 0 1 3160
box 0 0 1 1
use M1M2_CDNS_52468879185208  M1M2_CDNS_52468879185208_0
timestamp 1707688321
transform 0 -1 10268 -1 0 2084
box 0 0 192 244
use M1M2_CDNS_52468879185208  M1M2_CDNS_52468879185208_1
timestamp 1707688321
transform 0 -1 10268 -1 0 1287
box 0 0 192 244
use M1M2_CDNS_52468879185299  M1M2_CDNS_52468879185299_0
timestamp 1707688321
transform 1 0 6982 0 1 1692
box 0 0 704 52
use M1M2_CDNS_52468879185369  M1M2_CDNS_52468879185369_0
timestamp 1707688321
transform -1 0 6926 0 1 3512
box 0 0 1 1
use M1M2_CDNS_52468879185369  M1M2_CDNS_52468879185369_1
timestamp 1707688321
transform -1 0 9787 0 1 3389
box 0 0 1 1
use M1M2_CDNS_52468879185369  M1M2_CDNS_52468879185369_2
timestamp 1707688321
transform -1 0 9863 0 1 2116
box 0 0 1 1
use M1M2_CDNS_52468879185369  M1M2_CDNS_52468879185369_3
timestamp 1707688321
transform -1 0 6648 0 1 3240
box 0 0 1 1
use M1M2_CDNS_52468879185369  M1M2_CDNS_52468879185369_4
timestamp 1707688321
transform 0 -1 5885 1 0 1692
box 0 0 1 1
use M1M2_CDNS_52468879185369  M1M2_CDNS_52468879185369_5
timestamp 1707688321
transform 1 0 9074 0 -1 1062
box 0 0 1 1
use M1M2_CDNS_52468879185369  M1M2_CDNS_52468879185369_6
timestamp 1707688321
transform 1 0 9166 0 1 946
box 0 0 1 1
use M1M2_CDNS_52468879185369  M1M2_CDNS_52468879185369_7
timestamp 1707688321
transform 1 0 9166 0 1 321
box 0 0 1 1
use M1M2_CDNS_52468879185369  M1M2_CDNS_52468879185369_8
timestamp 1707688321
transform 1 0 5016 0 1 2642
box 0 0 1 1
use M1M2_CDNS_52468879185369  M1M2_CDNS_52468879185369_9
timestamp 1707688321
transform 1 0 6676 0 1 3240
box 0 0 1 1
use M1M2_CDNS_52468879185369  M1M2_CDNS_52468879185369_10
timestamp 1707688321
transform 1 0 8480 0 1 1532
box 0 0 1 1
use M1M2_CDNS_52468879185371  M1M2_CDNS_52468879185371_0
timestamp 1707688321
transform 0 1 9258 1 0 162
box 0 0 1 1
use M1M2_CDNS_52468879185371  M1M2_CDNS_52468879185371_1
timestamp 1707688321
transform 0 1 9258 1 0 349
box 0 0 1 1
use M1M2_CDNS_52468879185961  M1M2_CDNS_52468879185961_0
timestamp 1707688321
transform 0 -1 10268 1 0 1692
box 0 0 1 1
use M1M2_CDNS_52468879185972  M1M2_CDNS_52468879185972_0
timestamp 1707688321
transform 0 1 8715 -1 0 226
box 0 0 1 1
use M1M2_CDNS_52468879185972  M1M2_CDNS_52468879185972_1
timestamp 1707688321
transform 0 1 8715 -1 0 413
box 0 0 1 1
use M1M2_CDNS_52468879185972  M1M2_CDNS_52468879185972_2
timestamp 1707688321
transform 0 1 9551 1 0 68
box 0 0 1 1
use M1M2_CDNS_52468879185972  M1M2_CDNS_52468879185972_3
timestamp 1707688321
transform 0 1 9551 1 0 442
box 0 0 1 1
use M1M2_CDNS_52468879185972  M1M2_CDNS_52468879185972_4
timestamp 1707688321
transform 0 1 8140 1 0 68
box 0 0 1 1
use M1M2_CDNS_52468879185972  M1M2_CDNS_52468879185972_5
timestamp 1707688321
transform 0 1 8139 1 0 442
box 0 0 1 1
use M1M2_CDNS_52468879185972  M1M2_CDNS_52468879185972_6
timestamp 1707688321
transform 0 1 11044 1 0 349
box 0 0 1 1
use M1M2_CDNS_52468879185972  M1M2_CDNS_52468879185972_7
timestamp 1707688321
transform 0 1 11044 1 0 162
box 0 0 1 1
use M1M2_CDNS_52468879185972  M1M2_CDNS_52468879185972_8
timestamp 1707688321
transform 0 1 10303 1 0 3141
box 0 0 1 1
use M1M2_CDNS_52468879185975  M1M2_CDNS_52468879185975_0
timestamp 1707688321
transform 0 1 10113 -1 0 808
box 0 0 192 180
use M1M2_CDNS_52468879185975  M1M2_CDNS_52468879185975_1
timestamp 1707688321
transform 0 1 9258 -1 0 808
box 0 0 192 180
use M1M2_CDNS_52468879185975  M1M2_CDNS_52468879185975_2
timestamp 1707688321
transform 1 0 5348 0 -1 1052
box 0 0 192 180
use M1M2_CDNS_524688791851031  M1M2_CDNS_524688791851031_0
timestamp 1707688321
transform 0 1 11492 -1 0 3192
box 0 0 128 372
use M1M2_CDNS_524688791851032  M1M2_CDNS_524688791851032_0
timestamp 1707688321
transform 0 1 11492 -1 0 2611
box 0 0 192 372
use M1M2_CDNS_524688791851077  M1M2_CDNS_524688791851077_0
timestamp 1707688321
transform 1 0 6225 0 -1 1052
box 0 0 320 180
use M1M2_CDNS_524688791851077  M1M2_CDNS_524688791851077_1
timestamp 1707688321
transform 1 0 3981 0 1 1092
box 0 0 320 180
use M1M2_CDNS_524688791851077  M1M2_CDNS_524688791851077_2
timestamp 1707688321
transform 1 0 3981 0 1 1896
box 0 0 320 180
use M1M2_CDNS_524688791851185  M1M2_CDNS_524688791851185_0
timestamp 1707688321
transform 1 0 6225 0 -1 2592
box 0 0 320 244
use M1M2_CDNS_524688791851186  M1M2_CDNS_524688791851186_0
timestamp 1707688321
transform 0 1 8715 -1 0 808
box 0 0 192 308
use M1M2_CDNS_524688791851186  M1M2_CDNS_524688791851186_1
timestamp 1707688321
transform 1 0 920 0 1 741
box 0 0 192 308
use M1M2_CDNS_524688791851187  M1M2_CDNS_524688791851187_0
timestamp 1707688321
transform 1 0 7008 0 -1 2079
box 0 0 768 180
use M1M2_CDNS_524688791851193  M1M2_CDNS_524688791851193_0
timestamp 1707688321
transform 1 0 6982 0 -1 1283
box 0 0 704 180
use M1M2_CDNS_524688791851194  M1M2_CDNS_524688791851194_0
timestamp 1707688321
transform -1 0 4301 0 1 2116
box 0 0 320 436
use M2M3_CDNS_524688791851182  M2M3_CDNS_524688791851182_0
timestamp 1707688321
transform 1 0 3992 0 1 3462
box -5 0 301 794
use M2M3_CDNS_524688791851183  M2M3_CDNS_524688791851183_0
timestamp 1707688321
transform 1 0 5799 0 1 3378
box -5 0 61 794
use M2M3_CDNS_524688791851183  M2M3_CDNS_524688791851183_1
timestamp 1707688321
transform 1 0 3004 0 1 3378
box -5 0 61 794
use M2M3_CDNS_524688791851183  M2M3_CDNS_524688791851183_2
timestamp 1707688321
transform 1 0 13466 0 1 3458
box -5 0 61 794
use M2M3_CDNS_524688791851184  M2M3_CDNS_524688791851184_0
timestamp 1707688321
transform 1 0 14383 0 1 3458
box -5 0 141 794
use sky130_fd_io__sio_buf_localesd  sky130_fd_io__sio_buf_localesd_0
timestamp 1707688321
transform 1 0 19 0 1 349
box 0 -729 4014 4714
use sky130_fd_io__sio_com_inbuf_hv_dis  sky130_fd_io__sio_com_inbuf_hv_dis_0
timestamp 1707688321
transform -1 0 5827 0 -1 2418
box -74 -25 1622 2035
use sky130_fd_io__sio_com_inbuf_lv_dis  sky130_fd_io__sio_com_inbuf_lv_dis_0
timestamp 1707688321
transform 1 0 8097 0 1 123
box 0 -77 3817 1251
use sky130_fd_io__sio_com_m2m3_strap  sky130_fd_io__sio_com_m2m3_strap_0
timestamp 1707688321
transform -1 0 11832 0 -1 5644
box 0 0 364 858
use sky130_fd_io__sio_com_m2m3_strap  sky130_fd_io__sio_com_m2m3_strap_1
timestamp 1707688321
transform 0 -1 1485 1 0 3428
box 0 0 364 858
use sky130_fd_io__sio_com_m2m3_strap  sky130_fd_io__sio_com_m2m3_strap_2
timestamp 1707688321
transform 0 -1 2473 1 0 3428
box 0 0 364 858
use sky130_fd_io__sio_com_m2m3_strap  sky130_fd_io__sio_com_m2m3_strap_3
timestamp 1707688321
transform 1 0 11016 0 1 2070
box 0 0 364 858
use sky130_fd_io__sio_com_m2m3_strap  sky130_fd_io__sio_com_m2m3_strap_4
timestamp 1707688321
transform 1 0 12477 0 1 712
box 0 0 364 858
use sky130_fd_io__sio_com_m2m3_strap  sky130_fd_io__sio_com_m2m3_strap_5
timestamp 1707688321
transform 1 0 9523 0 1 712
box 0 0 364 858
use sky130_fd_io__sio_com_m2m3_strap  sky130_fd_io__sio_com_m2m3_strap_6
timestamp 1707688321
transform 1 0 8112 0 1 712
box 0 0 364 858
use sky130_fd_io__sio_com_m2m3_strap  sky130_fd_io__sio_com_m2m3_strap_7
timestamp 1707688321
transform 1 0 8687 0 1 2070
box 0 0 364 858
use sky130_fd_io__sio_com_m2m3_strap  sky130_fd_io__sio_com_m2m3_strap_8
timestamp 1707688321
transform 1 0 6961 0 1 3428
box 0 0 364 858
use sky130_fd_io__sio_com_m2m3_strap  sky130_fd_io__sio_com_m2m3_strap_9
timestamp 1707688321
transform 1 0 10272 0 1 4786
box 0 0 364 858
use sky130_fd_io__sio_com_m2m3_strap  sky130_fd_io__sio_com_m2m3_strap_10
timestamp 1707688321
transform 1 0 6203 0 1 4786
box 0 0 364 858
use sky130_fd_io__sio_com_m2m3_strap  sky130_fd_io__sio_com_m2m3_strap_11
timestamp 1707688321
transform 1 0 9271 0 1 3428
box 0 0 364 858
use sky130_fd_io__sio_com_m2m3_strap  sky130_fd_io__sio_com_m2m3_strap_12
timestamp 1707688321
transform 1 0 9928 0 1 3428
box 0 0 364 858
use sky130_fd_io__sio_com_m2m3_strap  sky130_fd_io__sio_com_m2m3_strap_13
timestamp 1707688321
transform 1 0 7455 0 1 3428
box 0 0 364 858
use sky130_fd_io__sio_ibuf_se  sky130_fd_io__sio_ibuf_se_0
timestamp 1707688321
transform 1 0 3800 0 1 3414
box -251 -3429 10369 3645
use sky130_fd_io__sio_ictl  sky130_fd_io__sio_ictl_0
timestamp 1707688321
transform -1 0 11206 0 1 430
box -210 -9 5801 2684
<< labels >>
flabel comment s 13688 1511 13688 1511 0 FreeSans 200 0 0 0 ibufmux_out_h_n
flabel comment s 10919 1513 10919 1513 0 FreeSans 200 0 0 0 ibufmux_out_h_n
flabel comment s 10284 1488 10284 1488 0 FreeSans 200 0 0 0 ibufmux_out_h_n
flabel comment s 6092 1480 6092 1480 0 FreeSans 200 0 0 0 ibufmux_out_h_n
flabel comment s 4120 2847 4120 2847 0 FreeSans 200 0 0 0 tripsel_i_h
flabel metal1 s 14425 855 14462 895 7 FreeSans 400 0 0 0 ibufmux_out_n
port 4 nsew
flabel metal1 s 14147 1486 14186 1532 7 FreeSans 400 0 0 0 ibufmux_out_h_n
port 5 nsew
flabel metal1 s 14262 1923 14305 1957 3 FreeSans 400 0 0 0 ie_diff_sel_h_n
port 2 nsew
flabel metal1 s 14346 1985 14389 2019 3 FreeSans 400 0 0 0 ie_diff_sel_h
port 3 nsew
flabel locali s 7751 1052 7785 1086 0 FreeSans 200 180 0 0 ie_diff_sel
port 6 nsew
flabel metal2 s 10296 5106 10604 5159 0 FreeSans 200 0 0 0 vcc_io
port 7 nsew
flabel metal2 s 7896 5112 7948 5159 7 FreeSans 200 90 0 0 dm_h_n<1>
port 8 nsew
flabel metal2 s 10088 5112 10124 5159 7 FreeSans 200 90 0 0 vtrip_sel_h_n
port 9 nsew
flabel metal2 s 8631 5112 8683 5159 7 FreeSans 200 90 0 0 dm_h_n<2>
port 10 nsew
flabel metal2 s 12892 5108 12944 5159 7 FreeSans 200 90 0 0 inp_dis_h_n
port 11 nsew
flabel metal2 s 8711 5112 8775 5159 7 FreeSans 200 90 0 0 dm_h<0>
port 12 nsew
flabel metal2 s 10880 5112 10932 5159 7 FreeSans 200 90 0 0 dm_h<2>
port 13 nsew
flabel metal2 s 10965 5090 11002 5142 3 FreeSans 200 270 0 0 dm_h<1>
port 14 nsew
flabel metal2 s 6610 0 6662 45 3 FreeSans 200 90 0 0 out_h
port 15 nsew
flabel metal2 s 9833 5112 9885 5159 7 FreeSans 200 90 0 0 vtrip_sel_h
port 16 nsew
flabel metal2 s 20 4944 136 4999 0 FreeSans 200 0 0 0 pad
port 17 nsew
flabel metal2 s 12576 467 12729 545 0 FreeSans 200 0 0 0 vpb_ka
port 18 nsew
flabel metal2 s 13429 5109 13555 5156 0 FreeSans 200 0 0 0 vgnd
port 19 nsew
flabel metal2 s 13864 5106 14149 5158 0 FreeSans 200 0 0 0 vgnd
port 19 nsew
flabel metal2 s 11040 5106 11356 5158 0 FreeSans 200 0 0 0 vpwr_ka
port 20 nsew
flabel metal2 s 6690 0 6742 45 3 FreeSans 200 90 0 0 out
port 21 nsew
flabel metal2 s 6596 5110 6648 5159 7 FreeSans 200 90 0 0 ibuf_sel_h
port 22 nsew
flabel metal2 s 6676 5110 6728 5159 7 FreeSans 200 90 0 0 ibuf_sel_h_n
port 23 nsew
flabel metal2 s 13606 5108 13658 5159 7 FreeSans 200 90 0 0 inp_dis_h
port 24 nsew
flabel metal2 s 1680 5118 1732 5159 7 FreeSans 200 90 0 0 dm_h_n<0>
port 25 nsew
flabel metal2 s 8296 5115 8348 5159 7 FreeSans 200 90 0 0 ie_diff_sel_n
port 26 nsew
<< properties >>
string GDS_END 85944678
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 85884042
string path 350.325 81.100 350.325 111.200 
<< end >>
