magic
tech sky130B
magscale 1 2
timestamp 1707688321
<< metal1 >>
rect 0 1 2 403
rect 2268 1 2270 403
use s8_esd_res250_sub_small  s8_esd_res250_sub_small_0
timestamp 1707688321
transform 1 0 0 0 1 0
box 0 0 2270 404
<< labels >>
flabel comment s 1156 206 1156 206 0 FreeSans 400 0 0 0 250 ohm
flabel metal1 s 2268 1 2270 403 0 FreeSans 400 0 0 0 rout
port 1 nsew
flabel metal1 s 0 1 2 403 0 FreeSans 200 0 0 0 pad
port 2 nsew
<< properties >>
string GDS_END 6066596
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 6065580
<< end >>
