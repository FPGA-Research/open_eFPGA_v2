magic
tech sky130A
magscale 1 2
timestamp 1707688321
<< nwell >>
rect -36 -36 89 1036
<< pdiff >>
rect 0 930 53 1000
rect 0 896 11 930
rect 45 896 53 930
rect 0 862 53 896
rect 0 828 11 862
rect 45 828 53 862
rect 0 794 53 828
rect 0 760 11 794
rect 45 760 53 794
rect 0 726 53 760
rect 0 692 11 726
rect 45 692 53 726
rect 0 658 53 692
rect 0 624 11 658
rect 45 624 53 658
rect 0 590 53 624
rect 0 556 11 590
rect 45 556 53 590
rect 0 522 53 556
rect 0 488 11 522
rect 45 488 53 522
rect 0 454 53 488
rect 0 420 11 454
rect 45 420 53 454
rect 0 386 53 420
rect 0 352 11 386
rect 45 352 53 386
rect 0 318 53 352
rect 0 284 11 318
rect 45 284 53 318
rect 0 250 53 284
rect 0 216 11 250
rect 45 216 53 250
rect 0 182 53 216
rect 0 148 11 182
rect 45 148 53 182
rect 0 114 53 148
rect 0 80 11 114
rect 45 80 53 114
rect 0 46 53 80
rect 0 12 11 46
rect 45 12 53 46
rect 0 0 53 12
<< pdiffc >>
rect 11 896 45 930
rect 11 828 45 862
rect 11 760 45 794
rect 11 692 45 726
rect 11 624 45 658
rect 11 556 45 590
rect 11 488 45 522
rect 11 420 45 454
rect 11 352 45 386
rect 11 284 45 318
rect 11 216 45 250
rect 11 148 45 182
rect 11 80 45 114
rect 11 12 45 46
<< locali >>
rect 11 930 45 932
rect 11 894 45 896
rect 11 822 45 828
rect 11 750 45 760
rect 11 678 45 692
rect 11 606 45 624
rect 11 534 45 556
rect 11 462 45 488
rect 11 390 45 420
rect 11 318 45 352
rect 11 250 45 284
rect 11 182 45 212
rect 11 114 45 140
rect 11 46 45 68
<< viali >>
rect 11 932 45 966
rect 11 862 45 894
rect 11 860 45 862
rect 11 794 45 822
rect 11 788 45 794
rect 11 726 45 750
rect 11 716 45 726
rect 11 658 45 678
rect 11 644 45 658
rect 11 590 45 606
rect 11 572 45 590
rect 11 522 45 534
rect 11 500 45 522
rect 11 454 45 462
rect 11 428 45 454
rect 11 386 45 390
rect 11 356 45 386
rect 11 284 45 318
rect 11 216 45 246
rect 11 212 45 216
rect 11 148 45 174
rect 11 140 45 148
rect 11 80 45 102
rect 11 68 45 80
rect 11 12 45 30
rect 11 -4 45 12
<< metal1 >>
rect 5 966 51 978
rect 5 932 11 966
rect 45 932 51 966
rect 5 894 51 932
rect 5 860 11 894
rect 45 860 51 894
rect 5 822 51 860
rect 5 788 11 822
rect 45 788 51 822
rect 5 750 51 788
rect 5 716 11 750
rect 45 716 51 750
rect 5 678 51 716
rect 5 644 11 678
rect 45 644 51 678
rect 5 606 51 644
rect 5 572 11 606
rect 45 572 51 606
rect 5 534 51 572
rect 5 500 11 534
rect 45 500 51 534
rect 5 462 51 500
rect 5 428 11 462
rect 45 428 51 462
rect 5 390 51 428
rect 5 356 11 390
rect 45 356 51 390
rect 5 318 51 356
rect 5 284 11 318
rect 45 284 51 318
rect 5 246 51 284
rect 5 212 11 246
rect 45 212 51 246
rect 5 174 51 212
rect 5 140 11 174
rect 45 140 51 174
rect 5 102 51 140
rect 5 68 11 102
rect 45 68 51 102
rect 5 30 51 68
rect 5 -4 11 30
rect 45 -4 51 30
rect 5 -16 51 -4
<< properties >>
string GDS_END 86590332
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 86588216
<< end >>
