magic
tech sky130B
timestamp 1707688321
<< locali >>
rect 17 0 36 17
rect 53 0 72 17
rect 89 0 108 17
rect 125 0 144 17
rect 161 0 180 17
rect 197 0 216 17
rect 233 0 252 17
rect 269 0 288 17
rect 305 0 324 17
rect 341 0 360 17
rect 377 0 396 17
rect 413 0 432 17
rect 449 0 468 17
rect 485 0 504 17
rect 521 0 540 17
rect 557 0 576 17
rect 593 0 612 17
rect 629 0 648 17
rect 665 0 684 17
rect 701 0 720 17
rect 737 0 756 17
rect 773 0 792 17
rect 809 0 828 17
rect 845 0 864 17
rect 881 0 900 17
rect 917 0 936 17
rect 953 0 972 17
rect 989 0 1008 17
rect 1025 0 1044 17
rect 1061 0 1080 17
rect 1097 0 1116 17
rect 1133 0 1152 17
rect 1169 0 1188 17
rect 1205 0 1224 17
rect 1241 0 1260 17
rect 1277 0 1296 17
rect 1313 0 1332 17
rect 1349 0 1368 17
rect 1385 0 1404 17
rect 1421 0 1440 17
rect 1457 0 1476 17
rect 1493 0 1512 17
rect 1529 0 1548 17
rect 1565 0 1584 17
rect 1601 0 1620 17
rect 1637 0 1656 17
rect 1673 0 1692 17
rect 1709 0 1728 17
rect 1745 0 1764 17
rect 1781 0 1800 17
rect 1817 0 1836 17
rect 1853 0 1872 17
rect 1889 0 1908 17
rect 1925 0 1944 17
rect 1961 0 1980 17
rect 1997 0 2016 17
rect 2033 0 2052 17
rect 2069 0 2088 17
rect 2105 0 2124 17
rect 2141 0 2160 17
rect 2177 0 2196 17
rect 2213 0 2232 17
rect 2249 0 2268 17
rect 2285 0 2304 17
rect 2321 0 2340 17
rect 2357 0 2376 17
rect 2393 0 2412 17
rect 2429 0 2448 17
rect 2465 0 2484 17
rect 2501 0 2520 17
rect 2537 0 2556 17
rect 2573 0 2592 17
rect 2609 0 2628 17
rect 2645 0 2664 17
rect 2681 0 2700 17
rect 2717 0 2736 17
rect 2753 0 2772 17
rect 2789 0 2808 17
rect 2825 0 2844 17
rect 2861 0 2880 17
rect 2897 0 2916 17
rect 2933 0 2952 17
rect 2969 0 2988 17
rect 3005 0 3024 17
rect 3041 0 3060 17
rect 3077 0 3096 17
rect 3113 0 3132 17
rect 3149 0 3168 17
rect 3185 0 3204 17
rect 3221 0 3240 17
rect 3257 0 3276 17
rect 3293 0 3312 17
rect 3329 0 3348 17
rect 3365 0 3384 17
rect 3401 0 3420 17
rect 3437 0 3456 17
rect 3473 0 3492 17
rect 3509 0 3528 17
rect 3545 0 3564 17
rect 3581 0 3600 17
rect 3617 0 3636 17
rect 3653 0 3672 17
rect 3689 0 3708 17
rect 3725 0 3744 17
rect 3761 0 3780 17
rect 3797 0 3816 17
rect 3833 0 3852 17
rect 3869 0 3888 17
rect 3905 0 3924 17
rect 3941 0 3960 17
rect 3977 0 3996 17
rect 4013 0 4032 17
rect 4049 0 4068 17
rect 4085 0 4104 17
rect 4121 0 4140 17
rect 4157 0 4176 17
rect 4193 0 4212 17
rect 4229 0 4248 17
rect 4265 0 4284 17
rect 4301 0 4320 17
rect 4337 0 4356 17
rect 4373 0 4392 17
rect 4409 0 4428 17
rect 4445 0 4464 17
rect 4481 0 4500 17
rect 4517 0 4536 17
rect 4553 0 4572 17
rect 4589 0 4608 17
rect 4625 0 4644 17
rect 4661 0 4680 17
rect 4697 0 4716 17
rect 4733 0 4752 17
rect 4769 0 4788 17
rect 4805 0 4824 17
rect 4841 0 4860 17
rect 4877 0 4896 17
rect 4913 0 4932 17
rect 4949 0 4968 17
rect 4985 0 5004 17
rect 5021 0 5040 17
rect 5057 0 5076 17
rect 5093 0 5112 17
rect 5129 0 5148 17
rect 5165 0 5184 17
rect 5201 0 5220 17
rect 5237 0 5256 17
rect 5273 0 5292 17
rect 5309 0 5328 17
rect 5345 0 5364 17
rect 5381 0 5400 17
rect 5417 0 5436 17
rect 5453 0 5472 17
rect 5489 0 5508 17
rect 5525 0 5544 17
rect 5561 0 5580 17
rect 5597 0 5616 17
rect 5633 0 5652 17
rect 5669 0 5688 17
rect 5705 0 5724 17
rect 5741 0 5760 17
rect 5777 0 5796 17
<< viali >>
rect 0 0 17 17
rect 36 0 53 17
rect 72 0 89 17
rect 108 0 125 17
rect 144 0 161 17
rect 180 0 197 17
rect 216 0 233 17
rect 252 0 269 17
rect 288 0 305 17
rect 324 0 341 17
rect 360 0 377 17
rect 396 0 413 17
rect 432 0 449 17
rect 468 0 485 17
rect 504 0 521 17
rect 540 0 557 17
rect 576 0 593 17
rect 612 0 629 17
rect 648 0 665 17
rect 684 0 701 17
rect 720 0 737 17
rect 756 0 773 17
rect 792 0 809 17
rect 828 0 845 17
rect 864 0 881 17
rect 900 0 917 17
rect 936 0 953 17
rect 972 0 989 17
rect 1008 0 1025 17
rect 1044 0 1061 17
rect 1080 0 1097 17
rect 1116 0 1133 17
rect 1152 0 1169 17
rect 1188 0 1205 17
rect 1224 0 1241 17
rect 1260 0 1277 17
rect 1296 0 1313 17
rect 1332 0 1349 17
rect 1368 0 1385 17
rect 1404 0 1421 17
rect 1440 0 1457 17
rect 1476 0 1493 17
rect 1512 0 1529 17
rect 1548 0 1565 17
rect 1584 0 1601 17
rect 1620 0 1637 17
rect 1656 0 1673 17
rect 1692 0 1709 17
rect 1728 0 1745 17
rect 1764 0 1781 17
rect 1800 0 1817 17
rect 1836 0 1853 17
rect 1872 0 1889 17
rect 1908 0 1925 17
rect 1944 0 1961 17
rect 1980 0 1997 17
rect 2016 0 2033 17
rect 2052 0 2069 17
rect 2088 0 2105 17
rect 2124 0 2141 17
rect 2160 0 2177 17
rect 2196 0 2213 17
rect 2232 0 2249 17
rect 2268 0 2285 17
rect 2304 0 2321 17
rect 2340 0 2357 17
rect 2376 0 2393 17
rect 2412 0 2429 17
rect 2448 0 2465 17
rect 2484 0 2501 17
rect 2520 0 2537 17
rect 2556 0 2573 17
rect 2592 0 2609 17
rect 2628 0 2645 17
rect 2664 0 2681 17
rect 2700 0 2717 17
rect 2736 0 2753 17
rect 2772 0 2789 17
rect 2808 0 2825 17
rect 2844 0 2861 17
rect 2880 0 2897 17
rect 2916 0 2933 17
rect 2952 0 2969 17
rect 2988 0 3005 17
rect 3024 0 3041 17
rect 3060 0 3077 17
rect 3096 0 3113 17
rect 3132 0 3149 17
rect 3168 0 3185 17
rect 3204 0 3221 17
rect 3240 0 3257 17
rect 3276 0 3293 17
rect 3312 0 3329 17
rect 3348 0 3365 17
rect 3384 0 3401 17
rect 3420 0 3437 17
rect 3456 0 3473 17
rect 3492 0 3509 17
rect 3528 0 3545 17
rect 3564 0 3581 17
rect 3600 0 3617 17
rect 3636 0 3653 17
rect 3672 0 3689 17
rect 3708 0 3725 17
rect 3744 0 3761 17
rect 3780 0 3797 17
rect 3816 0 3833 17
rect 3852 0 3869 17
rect 3888 0 3905 17
rect 3924 0 3941 17
rect 3960 0 3977 17
rect 3996 0 4013 17
rect 4032 0 4049 17
rect 4068 0 4085 17
rect 4104 0 4121 17
rect 4140 0 4157 17
rect 4176 0 4193 17
rect 4212 0 4229 17
rect 4248 0 4265 17
rect 4284 0 4301 17
rect 4320 0 4337 17
rect 4356 0 4373 17
rect 4392 0 4409 17
rect 4428 0 4445 17
rect 4464 0 4481 17
rect 4500 0 4517 17
rect 4536 0 4553 17
rect 4572 0 4589 17
rect 4608 0 4625 17
rect 4644 0 4661 17
rect 4680 0 4697 17
rect 4716 0 4733 17
rect 4752 0 4769 17
rect 4788 0 4805 17
rect 4824 0 4841 17
rect 4860 0 4877 17
rect 4896 0 4913 17
rect 4932 0 4949 17
rect 4968 0 4985 17
rect 5004 0 5021 17
rect 5040 0 5057 17
rect 5076 0 5093 17
rect 5112 0 5129 17
rect 5148 0 5165 17
rect 5184 0 5201 17
rect 5220 0 5237 17
rect 5256 0 5273 17
rect 5292 0 5309 17
rect 5328 0 5345 17
rect 5364 0 5381 17
rect 5400 0 5417 17
rect 5436 0 5453 17
rect 5472 0 5489 17
rect 5508 0 5525 17
rect 5544 0 5561 17
rect 5580 0 5597 17
rect 5616 0 5633 17
rect 5652 0 5669 17
rect 5688 0 5705 17
rect 5724 0 5741 17
rect 5760 0 5777 17
rect 5796 0 5813 17
<< metal1 >>
rect -6 17 5819 20
rect -6 0 0 17
rect 17 0 36 17
rect 53 0 72 17
rect 89 0 108 17
rect 125 0 144 17
rect 161 0 180 17
rect 197 0 216 17
rect 233 0 252 17
rect 269 0 288 17
rect 305 0 324 17
rect 341 0 360 17
rect 377 0 396 17
rect 413 0 432 17
rect 449 0 468 17
rect 485 0 504 17
rect 521 0 540 17
rect 557 0 576 17
rect 593 0 612 17
rect 629 0 648 17
rect 665 0 684 17
rect 701 0 720 17
rect 737 0 756 17
rect 773 0 792 17
rect 809 0 828 17
rect 845 0 864 17
rect 881 0 900 17
rect 917 0 936 17
rect 953 0 972 17
rect 989 0 1008 17
rect 1025 0 1044 17
rect 1061 0 1080 17
rect 1097 0 1116 17
rect 1133 0 1152 17
rect 1169 0 1188 17
rect 1205 0 1224 17
rect 1241 0 1260 17
rect 1277 0 1296 17
rect 1313 0 1332 17
rect 1349 0 1368 17
rect 1385 0 1404 17
rect 1421 0 1440 17
rect 1457 0 1476 17
rect 1493 0 1512 17
rect 1529 0 1548 17
rect 1565 0 1584 17
rect 1601 0 1620 17
rect 1637 0 1656 17
rect 1673 0 1692 17
rect 1709 0 1728 17
rect 1745 0 1764 17
rect 1781 0 1800 17
rect 1817 0 1836 17
rect 1853 0 1872 17
rect 1889 0 1908 17
rect 1925 0 1944 17
rect 1961 0 1980 17
rect 1997 0 2016 17
rect 2033 0 2052 17
rect 2069 0 2088 17
rect 2105 0 2124 17
rect 2141 0 2160 17
rect 2177 0 2196 17
rect 2213 0 2232 17
rect 2249 0 2268 17
rect 2285 0 2304 17
rect 2321 0 2340 17
rect 2357 0 2376 17
rect 2393 0 2412 17
rect 2429 0 2448 17
rect 2465 0 2484 17
rect 2501 0 2520 17
rect 2537 0 2556 17
rect 2573 0 2592 17
rect 2609 0 2628 17
rect 2645 0 2664 17
rect 2681 0 2700 17
rect 2717 0 2736 17
rect 2753 0 2772 17
rect 2789 0 2808 17
rect 2825 0 2844 17
rect 2861 0 2880 17
rect 2897 0 2916 17
rect 2933 0 2952 17
rect 2969 0 2988 17
rect 3005 0 3024 17
rect 3041 0 3060 17
rect 3077 0 3096 17
rect 3113 0 3132 17
rect 3149 0 3168 17
rect 3185 0 3204 17
rect 3221 0 3240 17
rect 3257 0 3276 17
rect 3293 0 3312 17
rect 3329 0 3348 17
rect 3365 0 3384 17
rect 3401 0 3420 17
rect 3437 0 3456 17
rect 3473 0 3492 17
rect 3509 0 3528 17
rect 3545 0 3564 17
rect 3581 0 3600 17
rect 3617 0 3636 17
rect 3653 0 3672 17
rect 3689 0 3708 17
rect 3725 0 3744 17
rect 3761 0 3780 17
rect 3797 0 3816 17
rect 3833 0 3852 17
rect 3869 0 3888 17
rect 3905 0 3924 17
rect 3941 0 3960 17
rect 3977 0 3996 17
rect 4013 0 4032 17
rect 4049 0 4068 17
rect 4085 0 4104 17
rect 4121 0 4140 17
rect 4157 0 4176 17
rect 4193 0 4212 17
rect 4229 0 4248 17
rect 4265 0 4284 17
rect 4301 0 4320 17
rect 4337 0 4356 17
rect 4373 0 4392 17
rect 4409 0 4428 17
rect 4445 0 4464 17
rect 4481 0 4500 17
rect 4517 0 4536 17
rect 4553 0 4572 17
rect 4589 0 4608 17
rect 4625 0 4644 17
rect 4661 0 4680 17
rect 4697 0 4716 17
rect 4733 0 4752 17
rect 4769 0 4788 17
rect 4805 0 4824 17
rect 4841 0 4860 17
rect 4877 0 4896 17
rect 4913 0 4932 17
rect 4949 0 4968 17
rect 4985 0 5004 17
rect 5021 0 5040 17
rect 5057 0 5076 17
rect 5093 0 5112 17
rect 5129 0 5148 17
rect 5165 0 5184 17
rect 5201 0 5220 17
rect 5237 0 5256 17
rect 5273 0 5292 17
rect 5309 0 5328 17
rect 5345 0 5364 17
rect 5381 0 5400 17
rect 5417 0 5436 17
rect 5453 0 5472 17
rect 5489 0 5508 17
rect 5525 0 5544 17
rect 5561 0 5580 17
rect 5597 0 5616 17
rect 5633 0 5652 17
rect 5669 0 5688 17
rect 5705 0 5724 17
rect 5741 0 5760 17
rect 5777 0 5796 17
rect 5813 0 5819 17
rect -6 -3 5819 0
<< properties >>
string GDS_END 78539446
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 78528946
<< end >>
