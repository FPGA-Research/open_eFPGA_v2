magic
tech sky130A
magscale 1 2
timestamp 1707688321
use padPLhp_CDNS_5246887918516  padPLhp_CDNS_5246887918516_0
timestamp 1707688321
transform 1 0 1500 0 1 24759
box -540 -540 12540 14540
<< properties >>
string GDS_END 85509694
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 85509640
<< end >>
