magic
tech sky130B
timestamp 1707688321
<< metal1 >>
rect 0 0 3 90
rect 253 0 256 90
<< via1 >>
rect 3 0 253 90
<< metal2 >>
rect 0 0 3 90
rect 253 0 256 90
<< properties >>
string GDS_END 79746460
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 79744792
<< end >>
