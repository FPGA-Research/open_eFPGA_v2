magic
tech sky130A
magscale 1 2
timestamp 1707688321
<< nwell >>
rect -38 261 866 582
<< pwell >>
rect 98 157 820 203
rect 1 21 820 157
rect 30 -17 64 21
<< locali >>
rect 212 401 278 493
rect 380 401 446 493
rect 212 391 446 401
rect 652 401 702 493
rect 652 391 810 401
rect 212 357 810 391
rect 86 215 156 255
rect 212 215 348 255
rect 390 215 628 255
rect 770 181 810 357
rect 652 127 810 181
<< obsli1 >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 828 561
rect 18 413 82 493
rect 18 323 52 413
rect 116 367 178 527
rect 312 435 346 527
rect 480 435 530 527
rect 568 435 618 527
rect 752 435 810 527
rect 18 289 730 323
rect 18 131 52 289
rect 664 215 730 289
rect 18 51 82 131
rect 116 17 178 181
rect 212 143 550 181
rect 212 51 278 143
rect 400 127 550 143
rect 312 17 362 109
rect 584 93 618 181
rect 400 51 810 93
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 828 17
<< obsli1c >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
<< metal1 >>
rect 0 561 828 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 828 561
rect 0 496 828 527
rect 0 17 828 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 828 17
rect 0 -48 828 -17
<< labels >>
rlabel locali s 86 215 156 255 6 A_N
port 1 nsew signal input
rlabel locali s 390 215 628 255 6 B
port 2 nsew signal input
rlabel locali s 212 215 348 255 6 C
port 3 nsew signal input
rlabel metal1 s 0 -48 828 48 8 VGND
port 4 nsew ground bidirectional abutment
rlabel pwell s 30 -17 64 21 6 VNB
port 5 nsew ground bidirectional
rlabel pwell s 1 21 820 157 6 VNB
port 5 nsew ground bidirectional
rlabel pwell s 98 157 820 203 6 VNB
port 5 nsew ground bidirectional
rlabel nwell s -38 261 866 582 6 VPB
port 6 nsew power bidirectional
rlabel metal1 s 0 496 828 592 6 VPWR
port 7 nsew power bidirectional abutment
rlabel locali s 652 127 810 181 6 Y
port 8 nsew signal output
rlabel locali s 770 181 810 357 6 Y
port 8 nsew signal output
rlabel locali s 212 357 810 391 6 Y
port 8 nsew signal output
rlabel locali s 652 391 810 401 6 Y
port 8 nsew signal output
rlabel locali s 652 401 702 493 6 Y
port 8 nsew signal output
rlabel locali s 212 391 446 401 6 Y
port 8 nsew signal output
rlabel locali s 380 401 446 493 6 Y
port 8 nsew signal output
rlabel locali s 212 401 278 493 6 Y
port 8 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 828 544
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_END 1850952
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_START 1844004
<< end >>
